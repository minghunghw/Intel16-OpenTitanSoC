module mem_tlul (clk_i,
    rst_ni,
    en_ifetch_i,
    tl_i,
    tl_o);
 input clk_i;
 input rst_ni;
 input [3:0] en_ifetch_i;
 input [108:0] tl_i;
 output [65:0] tl_o;

 wire N1;
 wire n126;
 wire n131;
 wire n170;
 wire n175;
 wire n188;
 wire n189;
 wire n192;
 wire n197;
 wire n211;
 wire n322;
 wire n323;
 wire n324;
 wire n325;
 wire n326;
 wire n327;
 wire n328;
 wire n329;
 wire n330;
 wire n331;
 wire n332;
 wire n333;
 wire n334;
 wire n335;
 wire n336;
 wire n337;
 wire n338;
 wire n339;
 wire n340;
 wire n341;
 wire n342;
 wire n343;
 wire n344;
 wire n345;
 wire n346;
 wire n347;
 wire n348;
 wire n349;
 wire n350;
 wire n351;
 wire n352;
 wire n353;
 wire n354;
 wire n355;
 wire n356;
 wire n357;
 wire n358;
 wire n359;
 wire n360;
 wire n361;
 wire n362;
 wire n363;
 wire n364;
 wire n365;
 wire n366;
 wire n367;
 wire n368;
 wire n369;
 wire n370;
 wire n371;
 wire n372;
 wire n373;
 wire n374;
 wire n375;
 wire n376;
 wire n377;
 wire n378;
 wire n379;
 wire n380;
 wire n381;
 wire n382;
 wire n383;
 wire n384;
 wire n385;
 wire n386;
 wire n387;
 wire n388;
 wire n389;
 wire n390;
 wire n391;
 wire n392;
 wire n393;
 wire n394;
 wire n395;
 wire n396;
 wire n397;
 wire n401;
 wire n402;
 wire n403;
 wire n404;
 wire n405;
 wire n409;
 wire n410;
 wire n411;
 wire n412;
 wire n413;
 wire n414;
 wire n415;
 wire n416;
 wire n417;
 wire n418;
 wire n419;
 wire n420;
 wire n421;
 wire n424;
 wire n426;
 wire n427;
 wire n428;
 wire n429;
 wire n430;
 wire n431;
 wire n432;
 wire n433;
 wire n434;
 wire n438;
 wire n439;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire n_0_net_;
 wire clknet_0_clk_i;
 wire rvalid;
 wire u_tlul_adapter_sram_N210;
 wire u_tlul_adapter_sram_reqfifo_wdata_op__0_;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_rptr_1_;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_wptr_1_;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_rptr_value_0_;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N11;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N23;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N25;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_wptr_value_0_;
 wire u_tlul_adapter_sram_u_reqfifo_net644;
 wire u_tlul_adapter_sram_u_reqfifo_net650;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_rptr_1_;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_wptr_1_;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_rptr_value_0_;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N11;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N23;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N25;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_wptr_value_0_;
 wire u_tlul_adapter_sram_u_rspfifo_net616;
 wire u_tlul_adapter_sram_u_rspfifo_net622;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_rptr_1_;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_wptr_1_;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_rptr_value_0_;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N11;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N23;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N25;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_wptr_value_0_;
 wire wen;
 wire net313;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_1_1__leaf_clk_i;
 wire clknet_0_u_tlul_adapter_sram_u_rspfifo_net616;
 wire clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net616;
 wire clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net616;
 wire clknet_0_u_tlul_adapter_sram_u_rspfifo_net622;
 wire clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622;
 wire clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622;
 wire clknet_0_u_tlul_adapter_sram_u_reqfifo_net644;
 wire clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net644;
 wire clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net644;
 wire clknet_0_u_tlul_adapter_sram_u_reqfifo_net650;
 wire clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net650;
 wire clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net650;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire [10:0] addr;
 wire [31:0] rdata;
 wire [31:0] u_tlul_adapter_sram_rdata_tlword;
 wire [16:0] u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata;
 wire [39:0] u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata;
 wire [4:0] u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata;
 wire [31:0] wdata;

 b15inv000as1n80x5 U430 (.a(net12),
    .o1(n328));
 b15nonb02aq1n16x5 U431 (.a(net57),
    .b(net186),
    .out0(addr[2]));
 b15nonb02ah1n16x5 U432 (.a(net56),
    .b(net187),
    .out0(addr[1]));
 b15nonb02ah1n16x5 U433 (.a(net55),
    .b(net187),
    .out0(addr[0]));
 b15nonb02ah1n16x5 U434 (.a(net191),
    .b(net187),
    .out0(addr[6]));
 b15nonb02ah1n16x5 U435 (.a(net59),
    .b(net187),
    .out0(addr[4]));
 b15nonb02as1n16x5 U436 (.a(net58),
    .b(net187),
    .out0(addr[3]));
 b15nonb02aq1n16x5 U437 (.a(net63),
    .b(net186),
    .out0(addr[8]));
 b15nonb02aq1n16x5 U438 (.a(net60),
    .b(net186),
    .out0(addr[5]));
 b15nonb02al1n04x5 U439 (.a(net190),
    .b(net187),
    .out0(addr[10]));
 b15nonb02al1n08x5 U440 (.a(net64),
    .b(net186),
    .out0(addr[9]));
 b15nonb02as1n16x5 U441 (.a(net62),
    .b(net186),
    .out0(addr[7]));
 b15norp03as1n24x5 U442 (.a(net11),
    .b(net10),
    .c(n328),
    .o1(wen));
 b15nandp2as1n32x5 U443 (.a(net199),
    .b(net174),
    .o1(n322));
 b15nonb02al1n16x5 U444 (.a(net24),
    .b(n322),
    .out0(wdata[7]));
 b15nonb02aq1n12x5 U445 (.a(net23),
    .b(n322),
    .out0(wdata[6]));
 b15nonb02aq1n12x5 U446 (.a(net22),
    .b(n322),
    .out0(wdata[5]));
 b15nonb02an1n12x5 U447 (.a(net21),
    .b(n322),
    .out0(wdata[4]));
 b15nonb02as1n08x5 U448 (.a(net20),
    .b(n322),
    .out0(wdata[3]));
 b15nonb02ah1n08x5 U449 (.a(net19),
    .b(n322),
    .out0(wdata[2]));
 b15nonb02al1n12x5 U450 (.a(net18),
    .b(n322),
    .out0(wdata[1]));
 b15nonb02aq1n08x5 U451 (.a(net17),
    .b(n322),
    .out0(wdata[0]));
 b15nand02ah1n48x5 U452 (.a(net196),
    .b(net174),
    .o1(n323));
 b15nonb02ah1n08x5 U453 (.a(net26),
    .b(n323),
    .out0(wdata[9]));
 b15nonb02al1n12x5 U454 (.a(net25),
    .b(n323),
    .out0(wdata[8]));
 b15nonb02ar1n16x5 U455 (.a(net28),
    .b(n323),
    .out0(wdata[11]));
 b15nonb02as1n08x5 U456 (.a(net27),
    .b(n323),
    .out0(wdata[10]));
 b15nonb02al1n16x5 U457 (.a(net32),
    .b(n323),
    .out0(wdata[15]));
 b15nonb02al1n16x5 U458 (.a(net31),
    .b(n323),
    .out0(wdata[14]));
 b15nonb02ah1n12x5 U459 (.a(net30),
    .b(n323),
    .out0(wdata[13]));
 b15nonb02al1n16x5 U460 (.a(net29),
    .b(n323),
    .out0(wdata[12]));
 b15inv000ah1n40x5 U461 (.a(wen),
    .o1(n_0_net_));
 b15inv020ar1n40x5 U462 (.a(net193),
    .o1(n347));
 b15norp02as1n48x5 U463 (.a(n347),
    .b(n_0_net_),
    .o1(n324));
 b15and002an1n16x5 U464 (.a(n324),
    .b(net48),
    .o(wdata[31]));
 b15and002an1n16x5 U465 (.a(n324),
    .b(net47),
    .o(wdata[30]));
 b15and002ah1n16x5 U466 (.a(n324),
    .b(net46),
    .o(wdata[29]));
 b15and002ar1n24x5 U467 (.a(n324),
    .b(net45),
    .o(wdata[28]));
 b15and002al1n24x5 U468 (.a(n324),
    .b(net44),
    .o(wdata[27]));
 b15and002as1n12x5 U469 (.a(n324),
    .b(net43),
    .o(wdata[26]));
 b15and002aq1n12x5 U470 (.a(n324),
    .b(net42),
    .o(wdata[25]));
 b15and002aq1n12x5 U471 (.a(n324),
    .b(net41),
    .o(wdata[24]));
 b15inv000ah1n12x5 U472 (.a(net194),
    .o1(n345));
 b15norp02ar1n32x5 U473 (.a(n345),
    .b(n_0_net_),
    .o1(n325));
 b15and002al1n16x5 U474 (.a(net156),
    .b(net40),
    .o(wdata[23]));
 b15and002aq1n16x5 U475 (.a(net156),
    .b(net39),
    .o(wdata[22]));
 b15and002ar1n24x5 U476 (.a(net156),
    .b(net38),
    .o(wdata[21]));
 b15and002al1n16x5 U477 (.a(net156),
    .b(net37),
    .o(wdata[20]));
 b15and002aq1n12x5 U478 (.a(net156),
    .b(net36),
    .o(wdata[19]));
 b15and002al1n16x5 U479 (.a(net156),
    .b(net35),
    .o(wdata[18]));
 b15and002al1n16x5 U480 (.a(net156),
    .b(net34),
    .o(wdata[17]));
 b15and002ah1n12x5 U481 (.a(n325),
    .b(net200),
    .o(wdata[16]));
 b15xor002an1n16x5 U482 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_wptr_1_),
    .b(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_rptr_1_),
    .out0(n360));
 b15inv020ah1n10x5 U483 (.a(net380),
    .o1(n327));
 b15inv040aq1n08x5 U484 (.a(net179),
    .o1(n365));
 b15aoi022ah1n24x5 U485 (.a(net179),
    .b(n327),
    .c(net380),
    .d(n365),
    .o1(n359));
 b15nanb02ah1n16x5 U486 (.a(n360),
    .b(net381),
    .out0(n418));
 b15inv000ah1n16x5 U487 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst),
    .o1(n356));
 b15xor002as1n12x5 U488 (.a(net406),
    .b(net183),
    .out0(n358));
 b15inv040al1n04x5 U489 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_rptr_1_),
    .o1(n326));
 b15aboi22aq1n24x5 U490 (.a(net584),
    .b(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_rptr_1_),
    .c(net584),
    .d(n326),
    .out0(n357));
 b15nanb02ah1n24x5 U491 (.a(net407),
    .b(n357),
    .out0(n384));
 b15nand02ah1n16x5 U492 (.a(n356),
    .b(net408),
    .o1(n374));
 b15inv040an1n08x5 U493 (.a(net409),
    .o1(n373));
 b15nandp2al1n24x5 U494 (.a(n373),
    .b(net481),
    .o1(n369));
 b15nonb03as1n12x5 U495 (.a(n418),
    .b(net178),
    .c(n369),
    .out0(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N23));
 b15nor002ah1n16x5 U496 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .b(n327),
    .o1(n175));
 b15aoi112as1n08x5 U497 (.a(net10),
    .b(n328),
    .c(net13),
    .d(net15),
    .o1(n355));
 b15norp02al1n12x5 U498 (.a(net193),
    .b(net195),
    .o1(n330));
 b15norp02an1n12x5 U499 (.a(net194),
    .b(net198),
    .o1(n329));
 b15inv040ah1n12x5 U500 (.a(net192),
    .o1(n343));
 b15aoi022al1n32x5 U501 (.a(net192),
    .b(n330),
    .c(n329),
    .d(n343),
    .o1(n331));
 b15aboi22ah1n24x5 U502 (.a(net189),
    .b(n331),
    .c(net198),
    .d(net195),
    .out0(n334));
 b15inv000ar1n03x5 U503 (.a(net8),
    .o1(n332));
 b15aoai13as1n08x5 U504 (.a(net194),
    .b(n332),
    .c(net198),
    .d(net195),
    .o1(n333));
 b15oai022ar1n24x5 U505 (.a(net8),
    .b(n334),
    .c(n333),
    .d(n347),
    .o1(n340));
 b15inv040as1n04x5 U506 (.a(net11),
    .o1(n439));
 b15inv040aq1n03x5 U507 (.a(net14),
    .o1(n336));
 b15nor004an1n03x5 U508 (.a(net4),
    .b(net1),
    .c(n439),
    .d(n336),
    .o1(n335));
 b15aoi013ar1n04x5 U509 (.a(net16),
    .b(net2),
    .c(net3),
    .d(n335),
    .o1(n338));
 b15obai22ar1n08x5 U510 (.a(net16),
    .b(net13),
    .c(net15),
    .d(n336),
    .out0(n337));
 b15aoi112aq1n06x5 U511 (.a(n338),
    .b(n337),
    .c(net189),
    .d(net192),
    .o1(n339));
 b15oai013ah1n08x5 U512 (.a(n339),
    .b(n340),
    .c(net9),
    .d(net11),
    .o1(n341));
 b15aoi012as1n06x5 U513 (.a(n341),
    .b(net9),
    .c(net11),
    .o1(n354));
 b15aoi022ah1n08x5 U514 (.a(net192),
    .b(net198),
    .c(net195),
    .d(n343),
    .o1(n344));
 b15nor002al1n12x5 U515 (.a(net54),
    .b(net194),
    .o1(n348));
 b15inv020as1n06x5 U516 (.a(net54),
    .o1(n342));
 b15norp03as1n16x5 U517 (.a(net198),
    .b(net195),
    .c(n342),
    .o1(n346));
 b15aoi022ah1n12x5 U518 (.a(n344),
    .b(n348),
    .c(n346),
    .d(n343),
    .o1(n351));
 b15aoi013as1n03x5 U519 (.a(net8),
    .b(net192),
    .c(n346),
    .d(n345),
    .o1(n350));
 b15aoai13as1n04x5 U520 (.a(net189),
    .b(n346),
    .c(n348),
    .d(n347),
    .o1(n349));
 b15oai112aq1n16x5 U521 (.a(n350),
    .b(n349),
    .c(net193),
    .d(n351),
    .o1(n353));
 b15oai013as1n12x5 U522 (.a(net8),
    .b(net54),
    .c(net192),
    .d(net189),
    .o1(n352));
 b15nand04as1n16x5 U523 (.a(n355),
    .b(n354),
    .c(n353),
    .d(n352),
    .o1(u_tlul_adapter_sram_N210));
 b15oai012aq1n32x5 U524 (.a(n356),
    .b(net407),
    .c(net585),
    .o1(n361));
 b15norp03as1n24x5 U525 (.a(wen),
    .b(n361),
    .c(u_tlul_adapter_sram_N210),
    .o1(N1));
 b15aoi012ar1n16x5 U526 (.a(net178),
    .b(n360),
    .c(net381),
    .o1(n362));
 b15nand02an1n24x5 U527 (.a(n362),
    .b(N1),
    .o1(n364));
 b15nor002an1n08x5 U528 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_wptr_1_),
    .b(n364),
    .o1(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N11));
 b15nonb02al1n08x5 U529 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .b(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_rptr_1_),
    .out0(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N25));
 b15nonb02aq1n16x5 U530 (.a(net382),
    .b(n361),
    .out0(net74));
 b15nand02ar1n24x5 U531 (.a(net12),
    .b(net74),
    .o1(n363));
 b15nor002ah1n06x5 U532 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_wptr_1_),
    .b(n363),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N11));
 b15inv020ah1n28x5 U533 (.a(n363),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9));
 b15nonb02ah1n16x5 U534 (.a(net183),
    .b(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .out0(n170));
 b15inv000ah1n20x5 U535 (.a(n364),
    .o1(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9));
 b15nor002ah1n16x5 U536 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .b(n365),
    .o1(n192));
 b15nonb02ah1n12x5 U537 (.a(n188),
    .b(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .out0(n189));
 b15inv040aq1n05x5 U538 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_rptr_1_),
    .o1(n372));
 b15obai22as1n16x5 U539 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_wptr_1_),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_rptr_1_),
    .c(n372),
    .d(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_wptr_1_),
    .out0(n367));
 b15inv020as1n10x5 U540 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_wptr_value_0_),
    .o1(n366));
 b15inv000as1n10x5 U541 (.a(net392),
    .o1(n370));
 b15aoi022aq1n32x5 U542 (.a(net392),
    .b(n366),
    .c(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_wptr_value_0_),
    .d(n370),
    .o1(n368));
 b15aoi112as1n08x5 U543 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst),
    .b(n369),
    .c(n367),
    .d(n368),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9));
 b15nor002ar1n16x5 U544 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .b(n366),
    .o1(n126));
 b15nonb02as1n16x5 U545 (.a(net393),
    .b(n367),
    .out0(n380));
 b15inv020as1n24x5 U546 (.a(net394),
    .o1(n386));
 b15ao0012al1n08x5 U547 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst),
    .b(net482),
    .c(net394),
    .o(n375));
 b15nanb02ah1n24x5 U548 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[16]),
    .b(net449),
    .out0(n379));
 b15nor004as1n12x5 U549 (.a(n375),
    .b(n379),
    .c(net409),
    .d(net399),
    .o1(n385));
 b15aob012as1n24x5 U550 (.a(net400),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[6]),
    .c(net395),
    .out0(net125));
 b15aob012as1n24x5 U551 (.a(net411),
    .b(net414),
    .c(net395),
    .out0(net101));
 b15aob012as1n24x5 U552 (.a(net411),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[4]),
    .c(net395),
    .out0(net121));
 b15nonb02as1n06x5 U553 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_wptr_1_),
    .out0(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N11));
 b15inv000al1n24x5 U554 (.a(net400),
    .o1(n382));
 b15nonb02aq1n16x5 U555 (.a(net6),
    .b(n382),
    .out0(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N23));
 b15norp02an1n08x5 U556 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .b(n370),
    .o1(n131));
 b15nor002as1n16x5 U557 (.a(net394),
    .b(net401),
    .o1(n371));
 b15and002an1n24x5 U558 (.a(net402),
    .b(net429),
    .o(net90));
 b15and002ah1n16x5 U559 (.a(net402),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[5]),
    .o(net124));
 b15and002ah1n16x5 U560 (.a(net402),
    .b(net420),
    .o(net126));
 b15and002ah1n16x5 U561 (.a(net402),
    .b(net417),
    .o(net111));
 b15and002ar1n08x5 U562 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .b(n372),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N25));
 b15nand02ah1n24x5 U563 (.a(n373),
    .b(net450),
    .o1(net122));
 b15inv020aq1n05x5 U564 (.a(net399),
    .o1(n377));
 b15aoai13as1n08x5 U565 (.a(net451),
    .b(net409),
    .c(n377),
    .d(net483),
    .o1(net123));
 b15inv000as1n48x5 U566 (.a(net484),
    .o1(n376));
 b15nonb02al1n12x5 U567 (.a(net529),
    .b(net139),
    .out0(net119));
 b15nonb02aq1n12x5 U568 (.a(net388),
    .b(net139),
    .out0(net113));
 b15nonb02as1n08x5 U569 (.a(net376),
    .b(net139),
    .out0(net117));
 b15nonb02as1n08x5 U570 (.a(net541),
    .b(net139),
    .out0(net110));
 b15nonb02as1n08x5 U571 (.a(net538),
    .b(net139),
    .out0(net115));
 b15nonb02ar1n12x5 U572 (.a(net559),
    .b(net139),
    .out0(net116));
 b15nonb02ar1n16x5 U573 (.a(net446),
    .b(net139),
    .out0(net114));
 b15nonb02ar1n16x5 U574 (.a(net523),
    .b(n376),
    .out0(net120));
 b15nonb02as1n08x5 U575 (.a(net385),
    .b(net139),
    .out0(net118));
 b15nonb02aq1n08x5 U576 (.a(net526),
    .b(net139),
    .out0(net112));
 b15nonb02ah1n16x5 U577 (.a(net6),
    .b(n376),
    .out0(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N23));
 b15nonb02ah1n16x5 U578 (.a(net184),
    .b(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .out0(n197));
 b15nonb02ar1n06x5 U579 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .b(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_rptr_1_),
    .out0(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N25));
 b15nandp2ah1n05x5 U580 (.a(net425),
    .b(net395),
    .o1(n378));
 b15oaoi13as1n08x5 U581 (.a(n376),
    .b(n377),
    .c(net450),
    .d(net426),
    .o1(net79));
 b15nandp2aq1n48x5 U582 (.a(net494),
    .b(net155),
    .o1(n397));
 b15nonb02as1n16x5 U583 (.a(rdata[26]),
    .b(net153),
    .out0(u_tlul_adapter_sram_rdata_tlword[26]));
 b15norp03as1n24x5 U584 (.a(net394),
    .b(net171),
    .c(net401),
    .o1(n381));
 b15inv000ar1n03x5 U585 (.a(net313),
    .o1(tl_o[9]));
 b15norp02ah1n24x5 U587 (.a(net395),
    .b(net401),
    .o1(n383));
 b15inv000ar1n03x5 U588 (.a(net314),
    .o1(tl_o[10]));
 b15aoi022an1n48x5 U590 (.a(net135),
    .b(net547),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[26]),
    .o1(n390));
 b15nand03an1n12x5 U591 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[12]),
    .b(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[11]),
    .c(net408),
    .o1(n388));
 b15aob012al1n16x5 U592 (.a(net400),
    .b(net171),
    .c(net395),
    .out0(n387));
 b15oai013as1n12x5 U593 (.a(n387),
    .b(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[13]),
    .c(net485),
    .d(n388),
    .o1(n389));
 b15inv000ar1n03x5 U594 (.a(net315),
    .o1(tl_o[11]));
 b15nand02ah1n06x5 U596 (.a(net548),
    .b(net130),
    .o1(net104));
 b15nonb02as1n16x5 U597 (.a(rdata[27]),
    .b(net153),
    .out0(u_tlul_adapter_sram_rdata_tlword[27]));
 b15aoi022al1n48x5 U598 (.a(net135),
    .b(net514),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[27]),
    .o1(n391));
 b15nand02al1n08x5 U599 (.a(net515),
    .b(net130),
    .o1(net105));
 b15nonb02ah1n16x5 U600 (.a(rdata[24]),
    .b(net153),
    .out0(u_tlul_adapter_sram_rdata_tlword[24]));
 b15aoi022ar1n32x5 U601 (.a(net135),
    .b(net532),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[24]),
    .o1(n392));
 b15inv000ar1n03x5 U602 (.a(net316),
    .o1(tl_o[12]));
 b15nandp2ar1n12x5 U603 (.a(net533),
    .b(net130),
    .o1(net102));
 b15nonb02ar1n04x5 U604 (.a(rdata[25]),
    .b(net153),
    .out0(u_tlul_adapter_sram_rdata_tlword[25]));
 b15aoi022ah1n32x5 U605 (.a(net135),
    .b(net556),
    .c(net131),
    .d(net150),
    .o1(n393));
 b15nandp2ah1n05x5 U606 (.a(net557),
    .b(net130),
    .o1(net103));
 b15nonb02as1n16x5 U607 (.a(rdata[30]),
    .b(net153),
    .out0(u_tlul_adapter_sram_rdata_tlword[30]));
 b15aoi022as1n32x5 U608 (.a(net135),
    .b(net553),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[30]),
    .o1(n394));
 b15qgbna2an1n05x5 U609 (.o1(net108),
    .a(net554),
    .b(net128));
 b15nonb02as1n16x5 U610 (.a(net201),
    .b(net495),
    .out0(u_tlul_adapter_sram_rdata_tlword[31]));
 b15aoi022ah1n48x5 U611 (.a(net135),
    .b(net499),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[31]),
    .o1(n395));
 b15nandp2al1n08x5 U612 (.a(net500),
    .b(net130),
    .o1(net109));
 b15nonb02as1n16x5 U613 (.a(rdata[28]),
    .b(net153),
    .out0(u_tlul_adapter_sram_rdata_tlword[28]));
 b15aoi022al1n06x5 U614 (.a(net138),
    .b(net470),
    .c(net134),
    .d(u_tlul_adapter_sram_rdata_tlword[28]),
    .o1(n396));
 b15nandp2ah1n03x5 U615 (.a(net471),
    .b(net128),
    .o1(net106));
 b15nonb02as1n16x5 U616 (.a(net202),
    .b(net495),
    .out0(u_tlul_adapter_sram_rdata_tlword[29]));
 b15aoi022ah1n48x5 U617 (.a(net135),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[37]),
    .c(net131),
    .d(net496),
    .o1(n401));
 b15qgbna2an1n05x5 U618 (.o1(net107),
    .a(net497),
    .b(net128));
 b15nandp2ar1n24x5 U619 (.a(net181),
    .b(net155),
    .o1(n434));
 b15nonb02as1n16x5 U620 (.a(rdata[20]),
    .b(net152),
    .out0(u_tlul_adapter_sram_rdata_tlword[20]));
 b15inv000ar1n03x5 U622 (.a(net317),
    .o1(tl_o[13]));
 b15aoi022aq1n48x5 U623 (.a(net135),
    .b(net571),
    .c(net131),
    .d(net149),
    .o1(n402));
 b15nandp2as1n03x5 U624 (.a(net572),
    .b(net128),
    .o1(net97));
 b15nonb02as1n16x5 U625 (.a(net204),
    .b(net152),
    .out0(u_tlul_adapter_sram_rdata_tlword[21]));
 b15aoi022an1n16x5 U626 (.a(net135),
    .b(net520),
    .c(net131),
    .d(net148),
    .o1(n403));
 b15nand02ah1n24x5 U627 (.a(net521),
    .b(net130),
    .o1(net98));
 b15nonb02as1n16x5 U628 (.a(net203),
    .b(net152),
    .out0(u_tlul_adapter_sram_rdata_tlword[22]));
 b15aoi022aq1n48x5 U629 (.a(net135),
    .b(net580),
    .c(net131),
    .d(net147),
    .o1(n404));
 b15nand02ar1n12x5 U630 (.a(net581),
    .b(net130),
    .o1(net99));
 b15nonb02as1n16x5 U631 (.a(rdata[23]),
    .b(net151),
    .out0(u_tlul_adapter_sram_rdata_tlword[23]));
 b15aoi022an1n48x5 U632 (.a(net135),
    .b(net550),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[23]),
    .o1(n405));
 b15nand02al1n08x5 U633 (.a(net551),
    .b(net130),
    .o1(net100));
 b15nandp2as1n48x5 U634 (.a(net458),
    .b(net155),
    .o1(n416));
 b15nonb02as1n16x5 U635 (.a(rdata[0]),
    .b(net459),
    .out0(u_tlul_adapter_sram_rdata_tlword[0]));
 b15inv000ar1n03x5 U637 (.a(net318),
    .o1(tl_o[14]));
 b15aoi022ar1n32x5 U638 (.a(net136),
    .b(net510),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[0]),
    .o1(n409));
 b15nandp2an1n12x5 U640 (.a(net511),
    .b(net127),
    .o1(net75));
 b15nonb02as1n16x5 U641 (.a(rdata[1]),
    .b(n416),
    .out0(u_tlul_adapter_sram_rdata_tlword[1]));
 b15aoi022as1n16x5 U642 (.a(net136),
    .b(net432),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[1]),
    .o1(n410));
 b15nandp2ah1n08x5 U643 (.a(net433),
    .b(net127),
    .o1(net76));
 b15nonb02as1n16x5 U644 (.a(rdata[2]),
    .b(net459),
    .out0(u_tlul_adapter_sram_rdata_tlword[2]));
 b15aoi022al1n32x5 U645 (.a(net136),
    .b(net503),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[2]),
    .o1(n411));
 b15nandp2al1n12x5 U646 (.a(net504),
    .b(net127),
    .o1(net77));
 b15nonb02as1n16x5 U647 (.a(rdata[3]),
    .b(n416),
    .out0(u_tlul_adapter_sram_rdata_tlword[3]));
 b15aoi022as1n16x5 U648 (.a(net136),
    .b(net442),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[3]),
    .o1(n412));
 b15nandp2ah1n08x5 U649 (.a(net443),
    .b(net486),
    .o1(net78));
 b15nonb02as1n16x5 U650 (.a(rdata[4]),
    .b(n416),
    .out0(u_tlul_adapter_sram_rdata_tlword[4]));
 b15aoi022ar1n32x5 U651 (.a(net137),
    .b(net454),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[4]),
    .o1(n413));
 b15nand02al1n32x5 U652 (.a(net455),
    .b(net129),
    .o1(net80));
 b15nonb02as1n16x5 U653 (.a(rdata[5]),
    .b(net459),
    .out0(u_tlul_adapter_sram_rdata_tlword[5]));
 b15aoi022aq1n24x5 U654 (.a(net136),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[13]),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[5]),
    .o1(n414));
 b15nand02al1n32x5 U655 (.a(n414),
    .b(net487),
    .o1(net81));
 b15nonb02as1n16x5 U656 (.a(rdata[6]),
    .b(net459),
    .out0(u_tlul_adapter_sram_rdata_tlword[6]));
 b15aoi022aq1n32x5 U657 (.a(net136),
    .b(net491),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[6]),
    .o1(n415));
 b15nand02ar1n16x5 U658 (.a(net492),
    .b(net127),
    .o1(net82));
 b15nonb02as1n16x5 U659 (.a(rdata[7]),
    .b(net459),
    .out0(u_tlul_adapter_sram_rdata_tlword[7]));
 b15aoi022aq1n32x5 U660 (.a(net136),
    .b(net166),
    .c(net132),
    .d(net460),
    .o1(n417));
 b15nand02aq1n12x5 U661 (.a(net461),
    .b(net127),
    .o1(net83));
 b15nandp2as1n48x5 U662 (.a(net474),
    .b(net155),
    .o1(n429));
 b15nonb02as1n16x5 U663 (.a(rdata[8]),
    .b(net475),
    .out0(u_tlul_adapter_sram_rdata_tlword[8]));
 b15aoi022ah1n32x5 U664 (.a(net136),
    .b(net165),
    .c(net132),
    .d(net476),
    .o1(n419));
 b15nand02aq1n24x5 U665 (.a(net477),
    .b(net127),
    .o1(net84));
 b15nonb02as1n16x5 U666 (.a(rdata[9]),
    .b(n429),
    .out0(u_tlul_adapter_sram_rdata_tlword[9]));
 b15aoi022aq1n32x5 U667 (.a(n381),
    .b(net437),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[9]),
    .o1(n420));
 b15nandp2ah1n16x5 U668 (.a(net438),
    .b(net127),
    .o1(net85));
 b15nonb02ar1n04x5 U669 (.a(rdata[10]),
    .b(net475),
    .out0(u_tlul_adapter_sram_rdata_tlword[10]));
 b15aoi022ah1n24x5 U670 (.a(net138),
    .b(net562),
    .c(net134),
    .d(net146),
    .o1(n421));
 b15nand02aq1n16x5 U671 (.a(net563),
    .b(net130),
    .o1(net86));
 b15nonb02as1n16x5 U672 (.a(rdata[11]),
    .b(n429),
    .out0(u_tlul_adapter_sram_rdata_tlword[11]));
 b15aoi022as1n16x5 U673 (.a(net136),
    .b(net465),
    .c(n383),
    .d(u_tlul_adapter_sram_rdata_tlword[11]),
    .o1(n424));
 b15nandp2aq1n24x5 U674 (.a(net466),
    .b(net127),
    .o1(net87));
 b15nonb02as1n16x5 U675 (.a(rdata[12]),
    .b(net475),
    .out0(u_tlul_adapter_sram_rdata_tlword[12]));
 b15aoi022aq1n32x5 U676 (.a(net138),
    .b(net574),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[12]),
    .o1(n426));
 b15nand02al1n24x5 U677 (.a(net575),
    .b(net130),
    .o1(net88));
 b15nonb02ar1n04x5 U678 (.a(rdata[13]),
    .b(net475),
    .out0(u_tlul_adapter_sram_rdata_tlword[13]));
 b15aoi022al1n32x5 U679 (.a(net138),
    .b(net577),
    .c(net134),
    .d(net145),
    .o1(n427));
 b15nand02ar1n24x5 U680 (.a(net578),
    .b(net130),
    .o1(net89));
 b15nonb02as1n16x5 U681 (.a(rdata[14]),
    .b(net475),
    .out0(u_tlul_adapter_sram_rdata_tlword[14]));
 b15aoi022al1n16x5 U682 (.a(net138),
    .b(net506),
    .c(net134),
    .d(u_tlul_adapter_sram_rdata_tlword[14]),
    .o1(n428));
 b15nandp2an1n05x5 U683 (.a(net507),
    .b(net128),
    .o1(net91));
 b15nonb02as1n16x5 U684 (.a(rdata[15]),
    .b(net475),
    .out0(u_tlul_adapter_sram_rdata_tlword[15]));
 b15aoi022ah1n32x5 U685 (.a(net135),
    .b(net565),
    .c(net134),
    .d(u_tlul_adapter_sram_rdata_tlword[15]),
    .o1(n430));
 b15nandp2ar1n24x5 U686 (.a(net566),
    .b(net130),
    .o1(net92));
 b15nonb02an1n16x5 U687 (.a(net207),
    .b(net152),
    .out0(u_tlul_adapter_sram_rdata_tlword[16]));
 b15aoi022aq1n32x5 U688 (.a(net135),
    .b(net544),
    .c(net131),
    .d(net144),
    .o1(n431));
 b15nandp2an1n04x5 U689 (.a(net545),
    .b(net128),
    .o1(net93));
 b15nonb02as1n16x5 U690 (.a(net206),
    .b(net152),
    .out0(u_tlul_adapter_sram_rdata_tlword[17]));
 b15aoi022ah1n48x5 U691 (.a(net135),
    .b(net568),
    .c(net131),
    .d(net143),
    .o1(n432));
 b15nandp2ah1n03x5 U692 (.a(net569),
    .b(net128),
    .o1(net94));
 b15nonb02as1n16x5 U693 (.a(net205),
    .b(net152),
    .out0(u_tlul_adapter_sram_rdata_tlword[18]));
 b15aoi022aq1n48x5 U694 (.a(net135),
    .b(net535),
    .c(net131),
    .d(net142),
    .o1(n433));
 b15nand02al1n08x5 U695 (.a(net536),
    .b(net130),
    .o1(net95));
 b15nonb02as1n16x5 U696 (.a(rdata[19]),
    .b(net152),
    .out0(u_tlul_adapter_sram_rdata_tlword[19]));
 b15aoi022as1n48x5 U697 (.a(net135),
    .b(net517),
    .c(net131),
    .d(net141),
    .o1(n438));
 b15nandp2aq1n05x5 U698 (.a(net518),
    .b(net128),
    .o1(net96));
 b15norp03as1n24x5 U700 (.a(net9),
    .b(net10),
    .c(n439),
    .o1(u_tlul_adapter_sram_reqfifo_wdata_op__0_));
 b15inv000ar1n03x5 U702 (.a(net319),
    .o1(tl_o[15]));
 b15inv000ar1n03x5 U704 (.a(net320),
    .o1(tl_o[48]));
 b15inv000ar1n03x5 U706 (.a(net321),
    .o1(tl_o[59]));
 b15inv000ar1n03x5 U708 (.a(net322),
    .o1(tl_o[60]));
 b15inv000ar1n03x5 U710 (.a(net323),
    .o1(tl_o[61]));
 b15inv000ar1n03x5 U712 (.a(net324),
    .o1(tl_o[63]));
 b15inv000ar1n03x5 U714 (.a(net325),
    .o1(tl_o[64]));
 b15ztpn00an1n08x5 PHY_5 ();
 b15ztpn00an1n08x5 PHY_4 ();
 b15ztpn00an1n08x5 PHY_3 ();
 b15ztpn00an1n08x5 PHY_2 ();
 b15ztpn00an1n08x5 PHY_1 ();
 b15ztpn00an1n08x5 PHY_0 ();
 b15fqy203ar1n02x5 rvalid_reg_u_tlul_adapter_sram_intg_error_q_reg (.rb(net197),
    .clk(clknet_1_1__leaf_clk_i),
    .d1(N1),
    .d2(net583),
    .o1(rvalid),
    .o2(n211),
    .si1(net208),
    .si2(net209),
    .ssb(net326));
 ip224uhdlp1p11rf_2048x32m8b2c1s0_t0r0p0d0a1m1h u_sram (.clkbyp(net210),
    .fwen(net211),
    .mcen(net215),
    .ren(net157),
    .wen(net174),
    .wpulseen(net327),
    .clk(clknet_1_1__leaf_clk_i),
    .adr({net176,
    net175,
    addr[8],
    addr[7],
    addr[6],
    addr[5],
    addr[4],
    addr[3],
    net177,
    addr[1],
    addr[0]}),
    .din({wdata[31],
    wdata[30],
    wdata[29],
    wdata[28],
    wdata[27],
    wdata[26],
    wdata[25],
    wdata[24],
    wdata[23],
    wdata[22],
    wdata[21],
    wdata[20],
    wdata[19],
    wdata[18],
    wdata[17],
    net154,
    wdata[15],
    wdata[14],
    wdata[13],
    wdata[12],
    wdata[11],
    wdata[10],
    wdata[9],
    wdata[8],
    wdata[7],
    wdata[6],
    wdata[5],
    wdata[4],
    wdata[3],
    wdata[2],
    wdata[1],
    wdata[0]}),
    .mc({net214,
    net213,
    net212}),
    .q({rdata[31],
    rdata[30],
    rdata[29],
    rdata[28],
    rdata[27],
    rdata[26],
    rdata[25],
    rdata[24],
    rdata[23],
    rdata[22],
    rdata[21],
    rdata[20],
    rdata[19],
    rdata[18],
    rdata[17],
    rdata[16],
    rdata[15],
    rdata[14],
    rdata[13],
    rdata[12],
    rdata[11],
    rdata[10],
    rdata[9],
    rdata[8],
    rdata[7],
    rdata[6],
    rdata[5],
    rdata[4],
    rdata[3],
    rdata[2],
    rdata[1],
    rdata[0]}),
    .wa({net217,
    net216}),
    .wpulse({net219,
    net218}));
 b15cilb05ah1n02x3 u_tlul_adapter_sram_u_reqfifo_clk_gate_gen_normal_fifo_storage_reg_0__0_latch (.clk(clknet_1_0__leaf_clk_i),
    .clkout(u_tlul_adapter_sram_u_reqfifo_net650),
    .en(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .te(net220));
 b15cilb05ah1n02x3 u_tlul_adapter_sram_u_reqfifo_clk_gate_gen_normal_fifo_storage_reg_0__latch (.clk(clknet_1_0__leaf_clk_i),
    .clkout(u_tlul_adapter_sram_u_reqfifo_net644),
    .en(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .te(net221));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__1_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net644),
    .d1(net66),
    .d2(net67),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[0]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[1]),
    .si1(net222),
    .si2(net223),
    .ssb(net328));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__11__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__12_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net650),
    .d1(net14),
    .d2(net15),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[11]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[12]),
    .si1(net224),
    .si2(net225),
    .ssb(net329));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__13__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__14_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net650),
    .d1(net16),
    .d2(u_tlul_adapter_sram_N210),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[13]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[14]),
    .si1(net226),
    .si2(net227),
    .ssb(net330));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__15__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__16_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net650),
    .d1(u_tlul_adapter_sram_reqfifo_wdata_op__0_),
    .d2(net228),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[15]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[16]),
    .si1(net229),
    .si2(net230),
    .ssb(net331));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__3_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net644),
    .d1(net68),
    .d2(net69),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[2]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[3]),
    .si1(net231),
    .si2(net232),
    .ssb(net332));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__5_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net644),
    .d1(net70),
    .d2(net71),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[4]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[5]),
    .si1(net233),
    .si2(net234),
    .ssb(net333));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__7_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net644),
    .d1(net72),
    .d2(net73),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[6]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[7]),
    .si1(net235),
    .si2(net236),
    .ssb(net334));
 b15fpy000ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__8_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net644),
    .d(net189),
    .o(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[8]),
    .si(net237),
    .ssb(net335));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__9__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__10_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net650),
    .d1(net8),
    .d2(net13),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[9]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[10]),
    .si1(net238),
    .si2(net239),
    .ssb(net336));
 b15fqy203ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0_ (.rb(net197),
    .clk(clknet_1_1__leaf_clk_i),
    .d1(n197),
    .d2(n170),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_rptr_value_0_),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_wptr_value_0_),
    .si1(net240),
    .si2(net241),
    .ssb(net337));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N25),
    .den(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .o(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_rptr_1_),
    .rb(net197),
    .si(net242),
    .ssb(net338));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N11),
    .den(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .o(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_wptr_1_),
    .rb(net197),
    .si(net243),
    .ssb(net339));
 b15fqy00car1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst_reg (.clk(clknet_1_1__leaf_clk_i),
    .d(net244),
    .o(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst),
    .psb(net197),
    .si(net245),
    .ssb(net340));
 b15cilb05ah1n02x3 u_tlul_adapter_sram_u_rspfifo_clk_gate_gen_normal_fifo_storage_reg_0__0_latch (.clk(clknet_1_0__leaf_clk_i),
    .clkout(u_tlul_adapter_sram_u_rspfifo_net622),
    .en(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .te(net246));
 b15cilb05ah1n02x3 u_tlul_adapter_sram_u_rspfifo_clk_gate_gen_normal_fifo_storage_reg_0__latch (.clk(clknet_1_1__leaf_clk_i),
    .clkout(u_tlul_adapter_sram_u_rspfifo_net616),
    .en(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .te(net247));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(net248),
    .d2(net249),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[0]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[1]),
    .si1(net250),
    .si2(net251),
    .ssb(net341));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__10__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__11_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(u_tlul_adapter_sram_rdata_tlword[2]),
    .d2(u_tlul_adapter_sram_rdata_tlword[3]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[10]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[11]),
    .si1(net252),
    .si2(net253),
    .ssb(net342));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__12__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__13_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(u_tlul_adapter_sram_rdata_tlword[4]),
    .d2(u_tlul_adapter_sram_rdata_tlword[5]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[12]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[13]),
    .si1(net254),
    .si2(net255),
    .ssb(net343));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__14__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__15_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[6]),
    .d2(u_tlul_adapter_sram_rdata_tlword[7]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[14]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[15]),
    .si1(net256),
    .si2(net257),
    .ssb(net344));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__16__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__17_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[8]),
    .d2(u_tlul_adapter_sram_rdata_tlword[9]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[16]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[17]),
    .si1(net258),
    .si2(net259),
    .ssb(net345));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__18__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__19_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(net146),
    .d2(u_tlul_adapter_sram_rdata_tlword[11]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[18]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[19]),
    .si1(net260),
    .si2(net261),
    .ssb(net346));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__20__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__21_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[12]),
    .d2(net145),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[20]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[21]),
    .si1(net262),
    .si2(net263),
    .ssb(net347));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__22__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__23_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[14]),
    .d2(u_tlul_adapter_sram_rdata_tlword[15]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[22]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[23]),
    .si1(net264),
    .si2(net265),
    .ssb(net348));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__24__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__25_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(net144),
    .d2(net143),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[24]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[25]),
    .si1(net266),
    .si2(net267),
    .ssb(net349));
 b15fpy000ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__26_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d(net142),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[26]),
    .si(net268),
    .ssb(net350));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__27__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__28_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(net141),
    .d2(net149),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[27]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[28]),
    .si1(net269),
    .si2(net270),
    .ssb(net351));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__29__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__30_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(net148),
    .d2(net147),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[29]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[30]),
    .si1(net271),
    .si2(net272),
    .ssb(net352));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(net273),
    .d2(net274),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[2]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[3]),
    .si1(net275),
    .si2(net276),
    .ssb(net353));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__31__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__32_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[23]),
    .d2(u_tlul_adapter_sram_rdata_tlword[24]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[31]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[32]),
    .si1(net277),
    .si2(net278),
    .ssb(net354));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__33__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__34_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(net150),
    .d2(u_tlul_adapter_sram_rdata_tlword[26]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[33]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[34]),
    .si1(net279),
    .si2(net280),
    .ssb(net355));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__35__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__36_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[27]),
    .d2(u_tlul_adapter_sram_rdata_tlword[28]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[35]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[36]),
    .si1(net281),
    .si2(net282),
    .ssb(net356));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__37__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__38_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[29]),
    .d2(u_tlul_adapter_sram_rdata_tlword[30]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[37]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[38]),
    .si1(net283),
    .si2(net284),
    .ssb(net357));
 b15fpy000ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__39_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d(u_tlul_adapter_sram_rdata_tlword[31]),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[39]),
    .si(net285),
    .ssb(net358));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(net286),
    .d2(net287),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[4]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[5]),
    .si1(net288),
    .si2(net289),
    .ssb(net359));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(net290),
    .d2(net291),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[6]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[7]),
    .si1(net292),
    .si2(net293),
    .ssb(net360));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__8__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__9_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(u_tlul_adapter_sram_rdata_tlword[0]),
    .d2(u_tlul_adapter_sram_rdata_tlword[1]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[8]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[9]),
    .si1(net294),
    .si2(net295),
    .ssb(net361));
 b15fqy203ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0_ (.rb(net197),
    .clk(clknet_1_0__leaf_clk_i),
    .d1(n131),
    .d2(n126),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_rptr_value_0_),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_wptr_value_0_),
    .si1(net296),
    .si2(net297),
    .ssb(net362));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N25),
    .den(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_rptr_1_),
    .rb(net197),
    .si(net298),
    .ssb(net363));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N11),
    .den(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_wptr_1_),
    .rb(net197),
    .si(net299),
    .ssb(net364));
 b15fqy00car1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst_reg (.clk(clknet_1_1__leaf_clk_i),
    .d(net300),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst),
    .psb(net197),
    .si(net301),
    .ssb(net365));
 b15fpy000ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__0_ (.clk(clknet_1_0__leaf_clk_i),
    .d(n189),
    .o(n188),
    .si(net302),
    .ssb(net366));
 b15fpy040ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__1_ (.clk(clknet_1_1__leaf_clk_i),
    .d(net199),
    .den(net140),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[1]),
    .si(net303),
    .ssb(net367));
 b15fpy040ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__2_ (.clk(clknet_1_1__leaf_clk_i),
    .d(net196),
    .den(net140),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[2]),
    .si(net304),
    .ssb(net368));
 b15fpy040ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__3_ (.clk(clknet_1_0__leaf_clk_i),
    .d(net51),
    .den(net140),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[3]),
    .si(net305),
    .ssb(net369));
 b15fpy040ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__4_ (.clk(clknet_1_0__leaf_clk_i),
    .d(net52),
    .den(net140),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[4]),
    .si(net306),
    .ssb(net370));
 b15fqy203ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0_ (.rb(net197),
    .clk(clknet_1_0__leaf_clk_i),
    .d1(n175),
    .d2(n192),
    .o1(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_rptr_value_0_),
    .o2(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_wptr_value_0_),
    .si1(net307),
    .si2(net308),
    .ssb(net371));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N25),
    .den(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_rptr_1_),
    .rb(net197),
    .si(net309),
    .ssb(net372));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N11),
    .den(net140),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_wptr_1_),
    .rb(net197),
    .si(net310),
    .ssb(net373));
 b15fqy00car1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst_reg (.clk(clknet_1_1__leaf_clk_i),
    .d(net311),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst),
    .psb(net197),
    .si(net312),
    .ssb(net374));
 b15tihi00an1n03x5 U585_313 (.o(net313));
 b15cbf000an1n16x5 clkbuf_0_clk_i (.clk(net375),
    .clkout(clknet_0_clk_i));
 b15ztpn00an1n08x5 PHY_6 ();
 b15ztpn00an1n08x5 PHY_7 ();
 b15ztpn00an1n08x5 PHY_8 ();
 b15ztpn00an1n08x5 PHY_9 ();
 b15ztpn00an1n08x5 PHY_10 ();
 b15ztpn00an1n08x5 PHY_11 ();
 b15ztpn00an1n08x5 PHY_12 ();
 b15ztpn00an1n08x5 PHY_13 ();
 b15ztpn00an1n08x5 PHY_14 ();
 b15ztpn00an1n08x5 PHY_15 ();
 b15ztpn00an1n08x5 PHY_16 ();
 b15ztpn00an1n08x5 PHY_17 ();
 b15ztpn00an1n08x5 PHY_18 ();
 b15ztpn00an1n08x5 PHY_19 ();
 b15ztpn00an1n08x5 PHY_20 ();
 b15ztpn00an1n08x5 PHY_21 ();
 b15ztpn00an1n08x5 PHY_22 ();
 b15ztpn00an1n08x5 PHY_23 ();
 b15ztpn00an1n08x5 PHY_24 ();
 b15ztpn00an1n08x5 PHY_25 ();
 b15ztpn00an1n08x5 PHY_26 ();
 b15ztpn00an1n08x5 PHY_27 ();
 b15ztpn00an1n08x5 PHY_28 ();
 b15ztpn00an1n08x5 PHY_29 ();
 b15ztpn00an1n08x5 PHY_30 ();
 b15ztpn00an1n08x5 PHY_31 ();
 b15ztpn00an1n08x5 PHY_32 ();
 b15ztpn00an1n08x5 PHY_33 ();
 b15ztpn00an1n08x5 PHY_34 ();
 b15ztpn00an1n08x5 PHY_35 ();
 b15ztpn00an1n08x5 PHY_36 ();
 b15ztpn00an1n08x5 PHY_37 ();
 b15ztpn00an1n08x5 PHY_38 ();
 b15ztpn00an1n08x5 PHY_39 ();
 b15ztpn00an1n08x5 PHY_40 ();
 b15ztpn00an1n08x5 PHY_41 ();
 b15ztpn00an1n08x5 PHY_42 ();
 b15ztpn00an1n08x5 PHY_43 ();
 b15ztpn00an1n08x5 PHY_44 ();
 b15ztpn00an1n08x5 PHY_45 ();
 b15ztpn00an1n08x5 PHY_46 ();
 b15ztpn00an1n08x5 PHY_47 ();
 b15ztpn00an1n08x5 PHY_48 ();
 b15ztpn00an1n08x5 PHY_49 ();
 b15ztpn00an1n08x5 PHY_50 ();
 b15ztpn00an1n08x5 PHY_51 ();
 b15ztpn00an1n08x5 PHY_52 ();
 b15ztpn00an1n08x5 PHY_53 ();
 b15ztpn00an1n08x5 PHY_54 ();
 b15ztpn00an1n08x5 PHY_55 ();
 b15ztpn00an1n08x5 PHY_56 ();
 b15ztpn00an1n08x5 PHY_57 ();
 b15ztpn00an1n08x5 PHY_58 ();
 b15ztpn00an1n08x5 PHY_59 ();
 b15ztpn00an1n08x5 PHY_60 ();
 b15ztpn00an1n08x5 PHY_61 ();
 b15ztpn00an1n08x5 PHY_62 ();
 b15ztpn00an1n08x5 PHY_63 ();
 b15ztpn00an1n08x5 PHY_64 ();
 b15ztpn00an1n08x5 PHY_65 ();
 b15ztpn00an1n08x5 PHY_66 ();
 b15ztpn00an1n08x5 PHY_67 ();
 b15ztpn00an1n08x5 PHY_68 ();
 b15ztpn00an1n08x5 PHY_69 ();
 b15ztpn00an1n08x5 PHY_70 ();
 b15ztpn00an1n08x5 PHY_71 ();
 b15ztpn00an1n08x5 PHY_72 ();
 b15ztpn00an1n08x5 PHY_73 ();
 b15ztpn00an1n08x5 PHY_74 ();
 b15ztpn00an1n08x5 PHY_75 ();
 b15ztpn00an1n08x5 PHY_76 ();
 b15ztpn00an1n08x5 PHY_77 ();
 b15ztpn00an1n08x5 PHY_78 ();
 b15ztpn00an1n08x5 PHY_79 ();
 b15ztpn00an1n08x5 PHY_80 ();
 b15ztpn00an1n08x5 PHY_81 ();
 b15ztpn00an1n08x5 PHY_82 ();
 b15ztpn00an1n08x5 PHY_83 ();
 b15ztpn00an1n08x5 PHY_84 ();
 b15ztpn00an1n08x5 PHY_85 ();
 b15ztpn00an1n08x5 PHY_86 ();
 b15ztpn00an1n08x5 PHY_87 ();
 b15ztpn00an1n08x5 PHY_88 ();
 b15ztpn00an1n08x5 PHY_89 ();
 b15ztpn00an1n08x5 PHY_90 ();
 b15ztpn00an1n08x5 PHY_91 ();
 b15ztpn00an1n08x5 PHY_92 ();
 b15ztpn00an1n08x5 PHY_93 ();
 b15ztpn00an1n08x5 PHY_94 ();
 b15ztpn00an1n08x5 PHY_95 ();
 b15ztpn00an1n08x5 PHY_96 ();
 b15ztpn00an1n08x5 PHY_97 ();
 b15ztpn00an1n08x5 PHY_98 ();
 b15ztpn00an1n08x5 PHY_99 ();
 b15ztpn00an1n08x5 PHY_100 ();
 b15ztpn00an1n08x5 PHY_101 ();
 b15ztpn00an1n08x5 PHY_102 ();
 b15ztpn00an1n08x5 PHY_103 ();
 b15ztpn00an1n08x5 PHY_104 ();
 b15ztpn00an1n08x5 PHY_105 ();
 b15ztpn00an1n08x5 PHY_106 ();
 b15ztpn00an1n08x5 PHY_107 ();
 b15ztpn00an1n08x5 PHY_108 ();
 b15ztpn00an1n08x5 PHY_109 ();
 b15ztpn00an1n08x5 PHY_110 ();
 b15ztpn00an1n08x5 PHY_111 ();
 b15ztpn00an1n08x5 PHY_112 ();
 b15ztpn00an1n08x5 PHY_113 ();
 b15ztpn00an1n08x5 PHY_114 ();
 b15ztpn00an1n08x5 PHY_115 ();
 b15ztpn00an1n08x5 PHY_116 ();
 b15ztpn00an1n08x5 PHY_117 ();
 b15ztpn00an1n08x5 PHY_118 ();
 b15ztpn00an1n08x5 PHY_119 ();
 b15ztpn00an1n08x5 PHY_120 ();
 b15ztpn00an1n08x5 PHY_121 ();
 b15ztpn00an1n08x5 PHY_122 ();
 b15ztpn00an1n08x5 PHY_123 ();
 b15ztpn00an1n08x5 PHY_124 ();
 b15ztpn00an1n08x5 PHY_125 ();
 b15ztpn00an1n08x5 PHY_126 ();
 b15ztpn00an1n08x5 PHY_127 ();
 b15ztpn00an1n08x5 PHY_128 ();
 b15ztpn00an1n08x5 PHY_129 ();
 b15ztpn00an1n08x5 PHY_130 ();
 b15ztpn00an1n08x5 PHY_131 ();
 b15ztpn00an1n08x5 PHY_132 ();
 b15ztpn00an1n08x5 PHY_133 ();
 b15ztpn00an1n08x5 PHY_134 ();
 b15ztpn00an1n08x5 PHY_135 ();
 b15ztpn00an1n08x5 PHY_136 ();
 b15ztpn00an1n08x5 PHY_137 ();
 b15ztpn00an1n08x5 PHY_138 ();
 b15ztpn00an1n08x5 PHY_139 ();
 b15ztpn00an1n08x5 PHY_140 ();
 b15ztpn00an1n08x5 PHY_141 ();
 b15ztpn00an1n08x5 PHY_142 ();
 b15ztpn00an1n08x5 PHY_143 ();
 b15ztpn00an1n08x5 PHY_144 ();
 b15ztpn00an1n08x5 PHY_145 ();
 b15ztpn00an1n08x5 PHY_146 ();
 b15ztpn00an1n08x5 PHY_147 ();
 b15ztpn00an1n08x5 PHY_148 ();
 b15ztpn00an1n08x5 PHY_149 ();
 b15ztpn00an1n08x5 PHY_150 ();
 b15ztpn00an1n08x5 PHY_151 ();
 b15ztpn00an1n08x5 PHY_152 ();
 b15ztpn00an1n08x5 PHY_153 ();
 b15ztpn00an1n08x5 PHY_154 ();
 b15ztpn00an1n08x5 PHY_155 ();
 b15ztpn00an1n08x5 PHY_156 ();
 b15ztpn00an1n08x5 PHY_157 ();
 b15ztpn00an1n08x5 PHY_158 ();
 b15ztpn00an1n08x5 PHY_159 ();
 b15ztpn00an1n08x5 PHY_160 ();
 b15ztpn00an1n08x5 PHY_161 ();
 b15ztpn00an1n08x5 PHY_162 ();
 b15ztpn00an1n08x5 PHY_163 ();
 b15ztpn00an1n08x5 PHY_164 ();
 b15ztpn00an1n08x5 PHY_165 ();
 b15ztpn00an1n08x5 PHY_166 ();
 b15ztpn00an1n08x5 PHY_167 ();
 b15ztpn00an1n08x5 PHY_168 ();
 b15ztpn00an1n08x5 PHY_169 ();
 b15ztpn00an1n08x5 PHY_170 ();
 b15ztpn00an1n08x5 PHY_171 ();
 b15ztpn00an1n08x5 PHY_172 ();
 b15ztpn00an1n08x5 PHY_173 ();
 b15ztpn00an1n08x5 PHY_174 ();
 b15ztpn00an1n08x5 PHY_175 ();
 b15ztpn00an1n08x5 PHY_176 ();
 b15ztpn00an1n08x5 PHY_177 ();
 b15ztpn00an1n08x5 PHY_178 ();
 b15ztpn00an1n08x5 PHY_179 ();
 b15ztpn00an1n08x5 PHY_180 ();
 b15ztpn00an1n08x5 PHY_181 ();
 b15ztpn00an1n08x5 PHY_182 ();
 b15ztpn00an1n08x5 PHY_183 ();
 b15ztpn00an1n08x5 PHY_184 ();
 b15ztpn00an1n08x5 PHY_185 ();
 b15ztpn00an1n08x5 PHY_186 ();
 b15ztpn00an1n08x5 PHY_187 ();
 b15ztpn00an1n08x5 PHY_188 ();
 b15ztpn00an1n08x5 PHY_189 ();
 b15ztpn00an1n08x5 PHY_190 ();
 b15ztpn00an1n08x5 PHY_191 ();
 b15ztpn00an1n08x5 PHY_192 ();
 b15ztpn00an1n08x5 PHY_193 ();
 b15ztpn00an1n08x5 PHY_194 ();
 b15ztpn00an1n08x5 PHY_195 ();
 b15ztpn00an1n08x5 PHY_196 ();
 b15ztpn00an1n08x5 PHY_197 ();
 b15ztpn00an1n08x5 PHY_198 ();
 b15ztpn00an1n08x5 PHY_199 ();
 b15ztpn00an1n08x5 PHY_200 ();
 b15ztpn00an1n08x5 PHY_201 ();
 b15ztpn00an1n08x5 PHY_202 ();
 b15ztpn00an1n08x5 PHY_203 ();
 b15ztpn00an1n08x5 PHY_204 ();
 b15ztpn00an1n08x5 PHY_205 ();
 b15ztpn00an1n08x5 PHY_206 ();
 b15ztpn00an1n08x5 PHY_207 ();
 b15ztpn00an1n08x5 PHY_208 ();
 b15ztpn00an1n08x5 PHY_209 ();
 b15ztpn00an1n08x5 PHY_210 ();
 b15ztpn00an1n08x5 PHY_211 ();
 b15ztpn00an1n08x5 PHY_212 ();
 b15ztpn00an1n08x5 PHY_213 ();
 b15ztpn00an1n08x5 PHY_214 ();
 b15ztpn00an1n08x5 PHY_215 ();
 b15ztpn00an1n08x5 PHY_216 ();
 b15ztpn00an1n08x5 PHY_217 ();
 b15ztpn00an1n08x5 PHY_218 ();
 b15ztpn00an1n08x5 PHY_219 ();
 b15ztpn00an1n08x5 PHY_220 ();
 b15ztpn00an1n08x5 PHY_221 ();
 b15ztpn00an1n08x5 PHY_222 ();
 b15ztpn00an1n08x5 PHY_223 ();
 b15ztpn00an1n08x5 PHY_224 ();
 b15ztpn00an1n08x5 PHY_225 ();
 b15ztpn00an1n08x5 PHY_226 ();
 b15ztpn00an1n08x5 PHY_227 ();
 b15ztpn00an1n08x5 PHY_228 ();
 b15ztpn00an1n08x5 PHY_229 ();
 b15ztpn00an1n08x5 PHY_230 ();
 b15ztpn00an1n08x5 PHY_231 ();
 b15ztpn00an1n08x5 PHY_232 ();
 b15ztpn00an1n08x5 PHY_233 ();
 b15ztpn00an1n08x5 PHY_234 ();
 b15ztpn00an1n08x5 PHY_235 ();
 b15ztpn00an1n08x5 PHY_236 ();
 b15ztpn00an1n08x5 PHY_237 ();
 b15ztpn00an1n08x5 PHY_238 ();
 b15ztpn00an1n08x5 PHY_239 ();
 b15ztpn00an1n08x5 PHY_240 ();
 b15ztpn00an1n08x5 PHY_241 ();
 b15ztpn00an1n08x5 PHY_242 ();
 b15ztpn00an1n08x5 PHY_243 ();
 b15ztpn00an1n08x5 PHY_244 ();
 b15ztpn00an1n08x5 PHY_245 ();
 b15ztpn00an1n08x5 PHY_246 ();
 b15ztpn00an1n08x5 PHY_247 ();
 b15ztpn00an1n08x5 PHY_248 ();
 b15ztpn00an1n08x5 PHY_249 ();
 b15ztpn00an1n08x5 PHY_250 ();
 b15ztpn00an1n08x5 PHY_251 ();
 b15ztpn00an1n08x5 PHY_252 ();
 b15ztpn00an1n08x5 PHY_253 ();
 b15ztpn00an1n08x5 PHY_254 ();
 b15ztpn00an1n08x5 PHY_255 ();
 b15ztpn00an1n08x5 PHY_256 ();
 b15ztpn00an1n08x5 PHY_257 ();
 b15ztpn00an1n08x5 PHY_258 ();
 b15ztpn00an1n08x5 PHY_259 ();
 b15ztpn00an1n08x5 PHY_260 ();
 b15ztpn00an1n08x5 PHY_261 ();
 b15ztpn00an1n08x5 PHY_262 ();
 b15ztpn00an1n08x5 PHY_263 ();
 b15ztpn00an1n08x5 PHY_264 ();
 b15ztpn00an1n08x5 PHY_265 ();
 b15ztpn00an1n08x5 PHY_266 ();
 b15ztpn00an1n08x5 PHY_267 ();
 b15ztpn00an1n08x5 PHY_268 ();
 b15ztpn00an1n08x5 PHY_269 ();
 b15ztpn00an1n08x5 PHY_270 ();
 b15ztpn00an1n08x5 PHY_271 ();
 b15ztpn00an1n08x5 PHY_272 ();
 b15ztpn00an1n08x5 PHY_273 ();
 b15ztpn00an1n08x5 PHY_274 ();
 b15ztpn00an1n08x5 PHY_275 ();
 b15ztpn00an1n08x5 PHY_276 ();
 b15ztpn00an1n08x5 PHY_277 ();
 b15ztpn00an1n08x5 PHY_278 ();
 b15ztpn00an1n08x5 PHY_279 ();
 b15ztpn00an1n08x5 PHY_280 ();
 b15ztpn00an1n08x5 PHY_281 ();
 b15ztpn00an1n08x5 PHY_282 ();
 b15ztpn00an1n08x5 PHY_283 ();
 b15ztpn00an1n08x5 PHY_284 ();
 b15ztpn00an1n08x5 PHY_285 ();
 b15ztpn00an1n08x5 PHY_286 ();
 b15ztpn00an1n08x5 PHY_287 ();
 b15ztpn00an1n08x5 PHY_288 ();
 b15ztpn00an1n08x5 PHY_289 ();
 b15ztpn00an1n08x5 PHY_290 ();
 b15ztpn00an1n08x5 PHY_291 ();
 b15ztpn00an1n08x5 PHY_292 ();
 b15ztpn00an1n08x5 PHY_293 ();
 b15ztpn00an1n08x5 PHY_294 ();
 b15ztpn00an1n08x5 PHY_295 ();
 b15ztpn00an1n08x5 PHY_296 ();
 b15ztpn00an1n08x5 PHY_297 ();
 b15ztpn00an1n08x5 PHY_298 ();
 b15ztpn00an1n08x5 PHY_299 ();
 b15ztpn00an1n08x5 PHY_300 ();
 b15ztpn00an1n08x5 PHY_301 ();
 b15ztpn00an1n08x5 PHY_302 ();
 b15ztpn00an1n08x5 PHY_303 ();
 b15ztpn00an1n08x5 PHY_304 ();
 b15ztpn00an1n08x5 PHY_305 ();
 b15ztpn00an1n08x5 PHY_306 ();
 b15ztpn00an1n08x5 PHY_307 ();
 b15ztpn00an1n08x5 PHY_308 ();
 b15ztpn00an1n08x5 PHY_309 ();
 b15ztpn00an1n08x5 PHY_310 ();
 b15ztpn00an1n08x5 PHY_311 ();
 b15ztpn00an1n08x5 PHY_312 ();
 b15ztpn00an1n08x5 PHY_313 ();
 b15ztpn00an1n08x5 PHY_314 ();
 b15ztpn00an1n08x5 PHY_315 ();
 b15ztpn00an1n08x5 PHY_316 ();
 b15ztpn00an1n08x5 PHY_317 ();
 b15ztpn00an1n08x5 PHY_318 ();
 b15ztpn00an1n08x5 PHY_319 ();
 b15ztpn00an1n08x5 PHY_320 ();
 b15ztpn00an1n08x5 PHY_321 ();
 b15ztpn00an1n08x5 PHY_322 ();
 b15ztpn00an1n08x5 PHY_323 ();
 b15ztpn00an1n08x5 PHY_324 ();
 b15ztpn00an1n08x5 PHY_325 ();
 b15ztpn00an1n08x5 PHY_326 ();
 b15ztpn00an1n08x5 PHY_327 ();
 b15ztpn00an1n08x5 PHY_328 ();
 b15ztpn00an1n08x5 PHY_329 ();
 b15ztpn00an1n08x5 PHY_330 ();
 b15ztpn00an1n08x5 PHY_331 ();
 b15ztpn00an1n08x5 PHY_332 ();
 b15ztpn00an1n08x5 PHY_333 ();
 b15ztpn00an1n08x5 PHY_334 ();
 b15ztpn00an1n08x5 PHY_335 ();
 b15ztpn00an1n08x5 PHY_336 ();
 b15ztpn00an1n08x5 PHY_337 ();
 b15ztpn00an1n08x5 PHY_338 ();
 b15ztpn00an1n08x5 PHY_339 ();
 b15ztpn00an1n08x5 PHY_340 ();
 b15ztpn00an1n08x5 PHY_341 ();
 b15ztpn00an1n08x5 PHY_342 ();
 b15ztpn00an1n08x5 PHY_343 ();
 b15ztpn00an1n08x5 PHY_344 ();
 b15ztpn00an1n08x5 PHY_345 ();
 b15ztpn00an1n08x5 PHY_346 ();
 b15ztpn00an1n08x5 PHY_347 ();
 b15ztpn00an1n08x5 PHY_348 ();
 b15ztpn00an1n08x5 PHY_349 ();
 b15ztpn00an1n08x5 PHY_350 ();
 b15ztpn00an1n08x5 PHY_351 ();
 b15ztpn00an1n08x5 PHY_352 ();
 b15ztpn00an1n08x5 PHY_353 ();
 b15ztpn00an1n08x5 PHY_354 ();
 b15ztpn00an1n08x5 PHY_355 ();
 b15ztpn00an1n08x5 PHY_356 ();
 b15ztpn00an1n08x5 PHY_357 ();
 b15ztpn00an1n08x5 PHY_358 ();
 b15ztpn00an1n08x5 PHY_359 ();
 b15ztpn00an1n08x5 PHY_360 ();
 b15ztpn00an1n08x5 PHY_361 ();
 b15ztpn00an1n08x5 PHY_362 ();
 b15ztpn00an1n08x5 PHY_363 ();
 b15ztpn00an1n08x5 PHY_364 ();
 b15ztpn00an1n08x5 PHY_365 ();
 b15ztpn00an1n08x5 PHY_366 ();
 b15ztpn00an1n08x5 PHY_367 ();
 b15ztpn00an1n08x5 PHY_368 ();
 b15ztpn00an1n08x5 PHY_369 ();
 b15ztpn00an1n08x5 PHY_370 ();
 b15ztpn00an1n08x5 PHY_371 ();
 b15ztpn00an1n08x5 PHY_372 ();
 b15ztpn00an1n08x5 PHY_373 ();
 b15ztpn00an1n08x5 PHY_374 ();
 b15ztpn00an1n08x5 PHY_375 ();
 b15ztpn00an1n08x5 PHY_376 ();
 b15ztpn00an1n08x5 PHY_377 ();
 b15ztpn00an1n08x5 PHY_378 ();
 b15ztpn00an1n08x5 PHY_379 ();
 b15ztpn00an1n08x5 PHY_380 ();
 b15ztpn00an1n08x5 PHY_381 ();
 b15ztpn00an1n08x5 PHY_382 ();
 b15ztpn00an1n08x5 PHY_383 ();
 b15ztpn00an1n08x5 PHY_384 ();
 b15ztpn00an1n08x5 PHY_385 ();
 b15ztpn00an1n08x5 PHY_386 ();
 b15ztpn00an1n08x5 PHY_387 ();
 b15ztpn00an1n08x5 PHY_388 ();
 b15ztpn00an1n08x5 PHY_389 ();
 b15ztpn00an1n08x5 PHY_390 ();
 b15ztpn00an1n08x5 PHY_391 ();
 b15ztpn00an1n08x5 PHY_392 ();
 b15ztpn00an1n08x5 PHY_393 ();
 b15ztpn00an1n08x5 PHY_394 ();
 b15ztpn00an1n08x5 PHY_395 ();
 b15ztpn00an1n08x5 PHY_396 ();
 b15ztpn00an1n08x5 PHY_397 ();
 b15ztpn00an1n08x5 PHY_398 ();
 b15ztpn00an1n08x5 PHY_399 ();
 b15ztpn00an1n08x5 PHY_400 ();
 b15ztpn00an1n08x5 PHY_401 ();
 b15ztpn00an1n08x5 PHY_402 ();
 b15ztpn00an1n08x5 PHY_403 ();
 b15ztpn00an1n08x5 PHY_404 ();
 b15ztpn00an1n08x5 PHY_405 ();
 b15ztpn00an1n08x5 PHY_406 ();
 b15ztpn00an1n08x5 PHY_407 ();
 b15ztpn00an1n08x5 PHY_408 ();
 b15ztpn00an1n08x5 PHY_409 ();
 b15ztpn00an1n08x5 PHY_410 ();
 b15ztpn00an1n08x5 PHY_411 ();
 b15ztpn00an1n08x5 PHY_412 ();
 b15ztpn00an1n08x5 PHY_413 ();
 b15ztpn00an1n08x5 PHY_414 ();
 b15ztpn00an1n08x5 PHY_415 ();
 b15ztpn00an1n08x5 PHY_416 ();
 b15ztpn00an1n08x5 PHY_417 ();
 b15ztpn00an1n08x5 PHY_418 ();
 b15ztpn00an1n08x5 PHY_419 ();
 b15ztpn00an1n08x5 PHY_420 ();
 b15ztpn00an1n08x5 PHY_421 ();
 b15ztpn00an1n08x5 PHY_422 ();
 b15ztpn00an1n08x5 PHY_423 ();
 b15ztpn00an1n08x5 PHY_424 ();
 b15ztpn00an1n08x5 PHY_425 ();
 b15ztpn00an1n08x5 PHY_426 ();
 b15ztpn00an1n08x5 PHY_427 ();
 b15ztpn00an1n08x5 PHY_428 ();
 b15ztpn00an1n08x5 PHY_429 ();
 b15ztpn00an1n08x5 PHY_430 ();
 b15ztpn00an1n08x5 PHY_431 ();
 b15ztpn00an1n08x5 PHY_432 ();
 b15ztpn00an1n08x5 PHY_433 ();
 b15ztpn00an1n08x5 PHY_434 ();
 b15ztpn00an1n08x5 PHY_435 ();
 b15ztpn00an1n08x5 PHY_436 ();
 b15ztpn00an1n08x5 PHY_437 ();
 b15ztpn00an1n08x5 PHY_438 ();
 b15ztpn00an1n08x5 PHY_439 ();
 b15ztpn00an1n08x5 PHY_440 ();
 b15ztpn00an1n08x5 PHY_441 ();
 b15ztpn00an1n08x5 PHY_442 ();
 b15ztpn00an1n08x5 PHY_443 ();
 b15ztpn00an1n08x5 PHY_444 ();
 b15ztpn00an1n08x5 PHY_445 ();
 b15ztpn00an1n08x5 PHY_446 ();
 b15ztpn00an1n08x5 PHY_447 ();
 b15ztpn00an1n08x5 PHY_448 ();
 b15ztpn00an1n08x5 PHY_449 ();
 b15ztpn00an1n08x5 PHY_450 ();
 b15ztpn00an1n08x5 PHY_451 ();
 b15ztpn00an1n08x5 PHY_452 ();
 b15ztpn00an1n08x5 PHY_453 ();
 b15ztpn00an1n08x5 PHY_454 ();
 b15ztpn00an1n08x5 PHY_455 ();
 b15ztpn00an1n08x5 PHY_456 ();
 b15ztpn00an1n08x5 PHY_457 ();
 b15ztpn00an1n08x5 PHY_458 ();
 b15ztpn00an1n08x5 PHY_459 ();
 b15ztpn00an1n08x5 PHY_460 ();
 b15ztpn00an1n08x5 PHY_461 ();
 b15ztpn00an1n08x5 PHY_462 ();
 b15ztpn00an1n08x5 PHY_463 ();
 b15ztpn00an1n08x5 PHY_464 ();
 b15ztpn00an1n08x5 PHY_465 ();
 b15ztpn00an1n08x5 PHY_466 ();
 b15ztpn00an1n08x5 PHY_467 ();
 b15ztpn00an1n08x5 PHY_468 ();
 b15ztpn00an1n08x5 PHY_469 ();
 b15ztpn00an1n08x5 PHY_470 ();
 b15ztpn00an1n08x5 PHY_471 ();
 b15ztpn00an1n08x5 PHY_472 ();
 b15ztpn00an1n08x5 PHY_473 ();
 b15ztpn00an1n08x5 PHY_474 ();
 b15ztpn00an1n08x5 PHY_475 ();
 b15ztpn00an1n08x5 PHY_476 ();
 b15ztpn00an1n08x5 PHY_477 ();
 b15ztpn00an1n08x5 PHY_478 ();
 b15ztpn00an1n08x5 PHY_479 ();
 b15ztpn00an1n08x5 PHY_480 ();
 b15ztpn00an1n08x5 PHY_481 ();
 b15ztpn00an1n08x5 PHY_482 ();
 b15ztpn00an1n08x5 PHY_483 ();
 b15ztpn00an1n08x5 PHY_484 ();
 b15ztpn00an1n08x5 PHY_485 ();
 b15ztpn00an1n08x5 PHY_486 ();
 b15ztpn00an1n08x5 PHY_487 ();
 b15ztpn00an1n08x5 PHY_488 ();
 b15ztpn00an1n08x5 PHY_489 ();
 b15ztpn00an1n08x5 PHY_490 ();
 b15ztpn00an1n08x5 PHY_491 ();
 b15ztpn00an1n08x5 PHY_492 ();
 b15ztpn00an1n08x5 PHY_493 ();
 b15ztpn00an1n08x5 PHY_494 ();
 b15ztpn00an1n08x5 PHY_495 ();
 b15ztpn00an1n08x5 PHY_496 ();
 b15ztpn00an1n08x5 PHY_497 ();
 b15ztpn00an1n08x5 PHY_498 ();
 b15ztpn00an1n08x5 PHY_499 ();
 b15ztpn00an1n08x5 PHY_500 ();
 b15ztpn00an1n08x5 PHY_501 ();
 b15ztpn00an1n08x5 PHY_502 ();
 b15ztpn00an1n08x5 PHY_503 ();
 b15ztpn00an1n08x5 PHY_504 ();
 b15ztpn00an1n08x5 PHY_505 ();
 b15ztpn00an1n08x5 PHY_506 ();
 b15ztpn00an1n08x5 PHY_507 ();
 b15ztpn00an1n08x5 PHY_508 ();
 b15ztpn00an1n08x5 PHY_509 ();
 b15ztpn00an1n08x5 PHY_510 ();
 b15ztpn00an1n08x5 PHY_511 ();
 b15ztpn00an1n08x5 PHY_512 ();
 b15ztpn00an1n08x5 PHY_513 ();
 b15ztpn00an1n08x5 PHY_514 ();
 b15ztpn00an1n08x5 PHY_515 ();
 b15ztpn00an1n08x5 PHY_516 ();
 b15ztpn00an1n08x5 PHY_517 ();
 b15ztpn00an1n08x5 PHY_518 ();
 b15ztpn00an1n08x5 PHY_519 ();
 b15ztpn00an1n08x5 PHY_520 ();
 b15ztpn00an1n08x5 PHY_521 ();
 b15ztpn00an1n08x5 PHY_522 ();
 b15ztpn00an1n08x5 PHY_523 ();
 b15ztpn00an1n08x5 PHY_524 ();
 b15ztpn00an1n08x5 PHY_525 ();
 b15ztpn00an1n08x5 PHY_526 ();
 b15ztpn00an1n08x5 PHY_527 ();
 b15ztpn00an1n08x5 PHY_528 ();
 b15ztpn00an1n08x5 PHY_529 ();
 b15ztpn00an1n08x5 PHY_530 ();
 b15ztpn00an1n08x5 PHY_531 ();
 b15ztpn00an1n08x5 PHY_532 ();
 b15ztpn00an1n08x5 PHY_533 ();
 b15ztpn00an1n08x5 PHY_534 ();
 b15ztpn00an1n08x5 PHY_535 ();
 b15ztpn00an1n08x5 PHY_536 ();
 b15ztpn00an1n08x5 PHY_537 ();
 b15ztpn00an1n08x5 PHY_538 ();
 b15ztpn00an1n08x5 PHY_539 ();
 b15ztpn00an1n08x5 PHY_540 ();
 b15ztpn00an1n08x5 PHY_541 ();
 b15ztpn00an1n08x5 PHY_542 ();
 b15ztpn00an1n08x5 PHY_543 ();
 b15ztpn00an1n08x5 PHY_544 ();
 b15ztpn00an1n08x5 PHY_545 ();
 b15ztpn00an1n08x5 PHY_546 ();
 b15ztpn00an1n08x5 PHY_547 ();
 b15ztpn00an1n08x5 PHY_548 ();
 b15ztpn00an1n08x5 PHY_549 ();
 b15ztpn00an1n08x5 PHY_550 ();
 b15ztpn00an1n08x5 PHY_551 ();
 b15ztpn00an1n08x5 PHY_552 ();
 b15ztpn00an1n08x5 PHY_553 ();
 b15ztpn00an1n08x5 PHY_554 ();
 b15ztpn00an1n08x5 PHY_555 ();
 b15ztpn00an1n08x5 PHY_556 ();
 b15ztpn00an1n08x5 PHY_557 ();
 b15ztpn00an1n08x5 PHY_558 ();
 b15ztpn00an1n08x5 PHY_559 ();
 b15ztpn00an1n08x5 PHY_560 ();
 b15ztpn00an1n08x5 PHY_561 ();
 b15ztpn00an1n08x5 PHY_562 ();
 b15ztpn00an1n08x5 PHY_563 ();
 b15ztpn00an1n08x5 PHY_564 ();
 b15ztpn00an1n08x5 PHY_565 ();
 b15ztpn00an1n08x5 PHY_566 ();
 b15ztpn00an1n08x5 PHY_567 ();
 b15ztpn00an1n08x5 PHY_568 ();
 b15ztpn00an1n08x5 PHY_569 ();
 b15ztpn00an1n08x5 PHY_570 ();
 b15ztpn00an1n08x5 PHY_571 ();
 b15ztpn00an1n08x5 PHY_572 ();
 b15ztpn00an1n08x5 PHY_573 ();
 b15ztpn00an1n08x5 PHY_574 ();
 b15ztpn00an1n08x5 PHY_575 ();
 b15ztpn00an1n08x5 PHY_576 ();
 b15ztpn00an1n08x5 PHY_577 ();
 b15ztpn00an1n08x5 PHY_578 ();
 b15ztpn00an1n08x5 PHY_579 ();
 b15ztpn00an1n08x5 PHY_580 ();
 b15ztpn00an1n08x5 PHY_581 ();
 b15ztpn00an1n08x5 PHY_582 ();
 b15ztpn00an1n08x5 PHY_583 ();
 b15ztpn00an1n08x5 TAP_584 ();
 b15ztpn00an1n08x5 TAP_585 ();
 b15ztpn00an1n08x5 TAP_586 ();
 b15ztpn00an1n08x5 TAP_587 ();
 b15ztpn00an1n08x5 TAP_588 ();
 b15ztpn00an1n08x5 TAP_589 ();
 b15ztpn00an1n08x5 TAP_590 ();
 b15ztpn00an1n08x5 TAP_591 ();
 b15ztpn00an1n08x5 TAP_592 ();
 b15ztpn00an1n08x5 TAP_593 ();
 b15ztpn00an1n08x5 TAP_594 ();
 b15ztpn00an1n08x5 TAP_595 ();
 b15ztpn00an1n08x5 TAP_596 ();
 b15ztpn00an1n08x5 TAP_597 ();
 b15ztpn00an1n08x5 TAP_598 ();
 b15ztpn00an1n08x5 TAP_599 ();
 b15ztpn00an1n08x5 TAP_600 ();
 b15ztpn00an1n08x5 TAP_601 ();
 b15ztpn00an1n08x5 TAP_602 ();
 b15ztpn00an1n08x5 TAP_603 ();
 b15ztpn00an1n08x5 TAP_604 ();
 b15ztpn00an1n08x5 TAP_605 ();
 b15ztpn00an1n08x5 TAP_606 ();
 b15ztpn00an1n08x5 TAP_607 ();
 b15ztpn00an1n08x5 TAP_608 ();
 b15ztpn00an1n08x5 TAP_609 ();
 b15ztpn00an1n08x5 TAP_610 ();
 b15ztpn00an1n08x5 TAP_611 ();
 b15ztpn00an1n08x5 TAP_612 ();
 b15ztpn00an1n08x5 TAP_613 ();
 b15ztpn00an1n08x5 TAP_614 ();
 b15ztpn00an1n08x5 TAP_615 ();
 b15ztpn00an1n08x5 TAP_616 ();
 b15ztpn00an1n08x5 TAP_617 ();
 b15ztpn00an1n08x5 TAP_618 ();
 b15ztpn00an1n08x5 TAP_619 ();
 b15ztpn00an1n08x5 TAP_620 ();
 b15ztpn00an1n08x5 TAP_621 ();
 b15ztpn00an1n08x5 TAP_622 ();
 b15ztpn00an1n08x5 TAP_623 ();
 b15ztpn00an1n08x5 TAP_624 ();
 b15ztpn00an1n08x5 TAP_625 ();
 b15ztpn00an1n08x5 TAP_626 ();
 b15ztpn00an1n08x5 TAP_627 ();
 b15ztpn00an1n08x5 TAP_628 ();
 b15ztpn00an1n08x5 TAP_629 ();
 b15ztpn00an1n08x5 TAP_630 ();
 b15ztpn00an1n08x5 TAP_631 ();
 b15ztpn00an1n08x5 TAP_632 ();
 b15ztpn00an1n08x5 TAP_633 ();
 b15ztpn00an1n08x5 TAP_634 ();
 b15ztpn00an1n08x5 TAP_635 ();
 b15ztpn00an1n08x5 TAP_636 ();
 b15ztpn00an1n08x5 TAP_637 ();
 b15ztpn00an1n08x5 TAP_638 ();
 b15ztpn00an1n08x5 TAP_639 ();
 b15ztpn00an1n08x5 TAP_640 ();
 b15ztpn00an1n08x5 TAP_641 ();
 b15ztpn00an1n08x5 TAP_642 ();
 b15ztpn00an1n08x5 TAP_643 ();
 b15ztpn00an1n08x5 TAP_644 ();
 b15ztpn00an1n08x5 TAP_645 ();
 b15ztpn00an1n08x5 TAP_646 ();
 b15ztpn00an1n08x5 TAP_647 ();
 b15ztpn00an1n08x5 TAP_648 ();
 b15ztpn00an1n08x5 TAP_649 ();
 b15ztpn00an1n08x5 TAP_650 ();
 b15ztpn00an1n08x5 TAP_651 ();
 b15ztpn00an1n08x5 TAP_652 ();
 b15ztpn00an1n08x5 TAP_653 ();
 b15ztpn00an1n08x5 TAP_654 ();
 b15ztpn00an1n08x5 TAP_655 ();
 b15ztpn00an1n08x5 TAP_656 ();
 b15ztpn00an1n08x5 TAP_657 ();
 b15ztpn00an1n08x5 TAP_658 ();
 b15ztpn00an1n08x5 TAP_659 ();
 b15ztpn00an1n08x5 TAP_660 ();
 b15ztpn00an1n08x5 TAP_661 ();
 b15ztpn00an1n08x5 TAP_662 ();
 b15ztpn00an1n08x5 TAP_663 ();
 b15ztpn00an1n08x5 TAP_664 ();
 b15ztpn00an1n08x5 TAP_665 ();
 b15ztpn00an1n08x5 TAP_666 ();
 b15ztpn00an1n08x5 TAP_667 ();
 b15ztpn00an1n08x5 TAP_668 ();
 b15ztpn00an1n08x5 TAP_669 ();
 b15ztpn00an1n08x5 TAP_670 ();
 b15ztpn00an1n08x5 TAP_671 ();
 b15ztpn00an1n08x5 TAP_672 ();
 b15ztpn00an1n08x5 TAP_673 ();
 b15ztpn00an1n08x5 TAP_674 ();
 b15ztpn00an1n08x5 TAP_675 ();
 b15ztpn00an1n08x5 TAP_676 ();
 b15ztpn00an1n08x5 TAP_677 ();
 b15ztpn00an1n08x5 TAP_678 ();
 b15ztpn00an1n08x5 TAP_679 ();
 b15ztpn00an1n08x5 TAP_680 ();
 b15ztpn00an1n08x5 TAP_681 ();
 b15ztpn00an1n08x5 TAP_682 ();
 b15ztpn00an1n08x5 TAP_683 ();
 b15ztpn00an1n08x5 TAP_684 ();
 b15ztpn00an1n08x5 TAP_685 ();
 b15ztpn00an1n08x5 TAP_686 ();
 b15ztpn00an1n08x5 TAP_687 ();
 b15ztpn00an1n08x5 TAP_688 ();
 b15ztpn00an1n08x5 TAP_689 ();
 b15ztpn00an1n08x5 TAP_690 ();
 b15ztpn00an1n08x5 TAP_691 ();
 b15ztpn00an1n08x5 TAP_692 ();
 b15ztpn00an1n08x5 TAP_693 ();
 b15ztpn00an1n08x5 TAP_694 ();
 b15ztpn00an1n08x5 TAP_695 ();
 b15ztpn00an1n08x5 TAP_696 ();
 b15ztpn00an1n08x5 TAP_697 ();
 b15ztpn00an1n08x5 TAP_698 ();
 b15ztpn00an1n08x5 TAP_699 ();
 b15ztpn00an1n08x5 TAP_700 ();
 b15ztpn00an1n08x5 TAP_701 ();
 b15ztpn00an1n08x5 TAP_702 ();
 b15ztpn00an1n08x5 TAP_703 ();
 b15ztpn00an1n08x5 TAP_704 ();
 b15ztpn00an1n08x5 TAP_705 ();
 b15ztpn00an1n08x5 TAP_706 ();
 b15ztpn00an1n08x5 TAP_707 ();
 b15ztpn00an1n08x5 TAP_708 ();
 b15ztpn00an1n08x5 TAP_709 ();
 b15ztpn00an1n08x5 TAP_710 ();
 b15ztpn00an1n08x5 TAP_711 ();
 b15ztpn00an1n08x5 TAP_712 ();
 b15ztpn00an1n08x5 TAP_713 ();
 b15ztpn00an1n08x5 TAP_714 ();
 b15ztpn00an1n08x5 TAP_715 ();
 b15ztpn00an1n08x5 TAP_716 ();
 b15ztpn00an1n08x5 TAP_717 ();
 b15ztpn00an1n08x5 TAP_718 ();
 b15ztpn00an1n08x5 TAP_719 ();
 b15ztpn00an1n08x5 TAP_720 ();
 b15ztpn00an1n08x5 TAP_721 ();
 b15ztpn00an1n08x5 TAP_722 ();
 b15ztpn00an1n08x5 TAP_723 ();
 b15ztpn00an1n08x5 TAP_724 ();
 b15ztpn00an1n08x5 TAP_725 ();
 b15ztpn00an1n08x5 TAP_726 ();
 b15ztpn00an1n08x5 TAP_727 ();
 b15ztpn00an1n08x5 TAP_728 ();
 b15ztpn00an1n08x5 TAP_729 ();
 b15ztpn00an1n08x5 TAP_730 ();
 b15ztpn00an1n08x5 TAP_731 ();
 b15ztpn00an1n08x5 TAP_732 ();
 b15ztpn00an1n08x5 TAP_733 ();
 b15ztpn00an1n08x5 TAP_734 ();
 b15ztpn00an1n08x5 TAP_735 ();
 b15ztpn00an1n08x5 TAP_736 ();
 b15ztpn00an1n08x5 TAP_737 ();
 b15ztpn00an1n08x5 TAP_738 ();
 b15ztpn00an1n08x5 TAP_739 ();
 b15ztpn00an1n08x5 TAP_740 ();
 b15ztpn00an1n08x5 TAP_741 ();
 b15ztpn00an1n08x5 TAP_742 ();
 b15ztpn00an1n08x5 TAP_743 ();
 b15ztpn00an1n08x5 TAP_744 ();
 b15ztpn00an1n08x5 TAP_745 ();
 b15ztpn00an1n08x5 TAP_746 ();
 b15ztpn00an1n08x5 TAP_747 ();
 b15ztpn00an1n08x5 TAP_748 ();
 b15ztpn00an1n08x5 TAP_749 ();
 b15ztpn00an1n08x5 TAP_750 ();
 b15ztpn00an1n08x5 TAP_751 ();
 b15ztpn00an1n08x5 TAP_752 ();
 b15ztpn00an1n08x5 TAP_753 ();
 b15ztpn00an1n08x5 TAP_754 ();
 b15ztpn00an1n08x5 TAP_755 ();
 b15ztpn00an1n08x5 TAP_756 ();
 b15ztpn00an1n08x5 TAP_757 ();
 b15ztpn00an1n08x5 TAP_758 ();
 b15ztpn00an1n08x5 TAP_759 ();
 b15ztpn00an1n08x5 TAP_760 ();
 b15ztpn00an1n08x5 TAP_761 ();
 b15ztpn00an1n08x5 TAP_762 ();
 b15ztpn00an1n08x5 TAP_763 ();
 b15ztpn00an1n08x5 TAP_764 ();
 b15ztpn00an1n08x5 TAP_765 ();
 b15ztpn00an1n08x5 TAP_766 ();
 b15ztpn00an1n08x5 TAP_767 ();
 b15ztpn00an1n08x5 TAP_768 ();
 b15ztpn00an1n08x5 TAP_769 ();
 b15ztpn00an1n08x5 TAP_770 ();
 b15ztpn00an1n08x5 TAP_771 ();
 b15ztpn00an1n08x5 TAP_772 ();
 b15ztpn00an1n08x5 TAP_773 ();
 b15ztpn00an1n08x5 TAP_774 ();
 b15ztpn00an1n08x5 TAP_775 ();
 b15ztpn00an1n08x5 TAP_776 ();
 b15ztpn00an1n08x5 TAP_777 ();
 b15ztpn00an1n08x5 TAP_778 ();
 b15ztpn00an1n08x5 TAP_779 ();
 b15ztpn00an1n08x5 TAP_780 ();
 b15ztpn00an1n08x5 TAP_781 ();
 b15ztpn00an1n08x5 TAP_782 ();
 b15ztpn00an1n08x5 TAP_783 ();
 b15ztpn00an1n08x5 TAP_784 ();
 b15ztpn00an1n08x5 TAP_785 ();
 b15ztpn00an1n08x5 TAP_786 ();
 b15ztpn00an1n08x5 TAP_787 ();
 b15ztpn00an1n08x5 TAP_788 ();
 b15ztpn00an1n08x5 TAP_789 ();
 b15ztpn00an1n08x5 TAP_790 ();
 b15ztpn00an1n08x5 TAP_791 ();
 b15ztpn00an1n08x5 TAP_792 ();
 b15ztpn00an1n08x5 TAP_793 ();
 b15ztpn00an1n08x5 TAP_794 ();
 b15ztpn00an1n08x5 TAP_795 ();
 b15ztpn00an1n08x5 TAP_796 ();
 b15ztpn00an1n08x5 TAP_797 ();
 b15ztpn00an1n08x5 TAP_798 ();
 b15ztpn00an1n08x5 TAP_799 ();
 b15ztpn00an1n08x5 TAP_800 ();
 b15ztpn00an1n08x5 TAP_801 ();
 b15ztpn00an1n08x5 TAP_802 ();
 b15ztpn00an1n08x5 TAP_803 ();
 b15ztpn00an1n08x5 TAP_804 ();
 b15ztpn00an1n08x5 TAP_805 ();
 b15ztpn00an1n08x5 TAP_806 ();
 b15ztpn00an1n08x5 TAP_807 ();
 b15ztpn00an1n08x5 TAP_808 ();
 b15ztpn00an1n08x5 TAP_809 ();
 b15ztpn00an1n08x5 TAP_810 ();
 b15ztpn00an1n08x5 TAP_811 ();
 b15ztpn00an1n08x5 TAP_812 ();
 b15ztpn00an1n08x5 TAP_813 ();
 b15ztpn00an1n08x5 TAP_814 ();
 b15ztpn00an1n08x5 TAP_815 ();
 b15ztpn00an1n08x5 TAP_816 ();
 b15ztpn00an1n08x5 TAP_817 ();
 b15ztpn00an1n08x5 TAP_818 ();
 b15ztpn00an1n08x5 TAP_819 ();
 b15ztpn00an1n08x5 TAP_820 ();
 b15ztpn00an1n08x5 TAP_821 ();
 b15ztpn00an1n08x5 TAP_822 ();
 b15ztpn00an1n08x5 TAP_823 ();
 b15ztpn00an1n08x5 TAP_824 ();
 b15ztpn00an1n08x5 TAP_825 ();
 b15ztpn00an1n08x5 TAP_826 ();
 b15ztpn00an1n08x5 TAP_827 ();
 b15ztpn00an1n08x5 TAP_828 ();
 b15ztpn00an1n08x5 TAP_829 ();
 b15ztpn00an1n08x5 TAP_830 ();
 b15ztpn00an1n08x5 TAP_831 ();
 b15ztpn00an1n08x5 TAP_832 ();
 b15ztpn00an1n08x5 TAP_833 ();
 b15ztpn00an1n08x5 TAP_834 ();
 b15ztpn00an1n08x5 TAP_835 ();
 b15ztpn00an1n08x5 TAP_836 ();
 b15ztpn00an1n08x5 TAP_837 ();
 b15ztpn00an1n08x5 TAP_838 ();
 b15ztpn00an1n08x5 TAP_839 ();
 b15ztpn00an1n08x5 TAP_840 ();
 b15ztpn00an1n08x5 TAP_841 ();
 b15ztpn00an1n08x5 TAP_842 ();
 b15ztpn00an1n08x5 TAP_843 ();
 b15ztpn00an1n08x5 TAP_844 ();
 b15ztpn00an1n08x5 TAP_845 ();
 b15ztpn00an1n08x5 TAP_846 ();
 b15ztpn00an1n08x5 TAP_847 ();
 b15ztpn00an1n08x5 TAP_848 ();
 b15ztpn00an1n08x5 TAP_849 ();
 b15ztpn00an1n08x5 TAP_850 ();
 b15ztpn00an1n08x5 TAP_851 ();
 b15ztpn00an1n08x5 TAP_852 ();
 b15ztpn00an1n08x5 TAP_853 ();
 b15ztpn00an1n08x5 TAP_854 ();
 b15ztpn00an1n08x5 TAP_855 ();
 b15ztpn00an1n08x5 TAP_856 ();
 b15ztpn00an1n08x5 TAP_857 ();
 b15ztpn00an1n08x5 TAP_858 ();
 b15ztpn00an1n08x5 TAP_859 ();
 b15ztpn00an1n08x5 TAP_860 ();
 b15ztpn00an1n08x5 TAP_861 ();
 b15ztpn00an1n08x5 TAP_862 ();
 b15ztpn00an1n08x5 TAP_863 ();
 b15ztpn00an1n08x5 TAP_864 ();
 b15ztpn00an1n08x5 TAP_865 ();
 b15ztpn00an1n08x5 TAP_866 ();
 b15ztpn00an1n08x5 TAP_867 ();
 b15ztpn00an1n08x5 TAP_868 ();
 b15ztpn00an1n08x5 TAP_869 ();
 b15ztpn00an1n08x5 TAP_870 ();
 b15ztpn00an1n08x5 TAP_871 ();
 b15ztpn00an1n08x5 TAP_872 ();
 b15ztpn00an1n08x5 TAP_873 ();
 b15ztpn00an1n08x5 TAP_874 ();
 b15ztpn00an1n08x5 TAP_875 ();
 b15ztpn00an1n08x5 TAP_876 ();
 b15ztpn00an1n08x5 TAP_877 ();
 b15ztpn00an1n08x5 TAP_878 ();
 b15bfn000as1n02x5 input1 (.a(en_ifetch_i[0]),
    .o(net1));
 b15bfn000as1n02x5 input2 (.a(en_ifetch_i[1]),
    .o(net2));
 b15bfn000as1n02x5 input3 (.a(en_ifetch_i[2]),
    .o(net3));
 b15bfn000as1n02x5 input4 (.a(en_ifetch_i[3]),
    .o(net4));
 b15bfn001as1n16x5 input5 (.a(rst_ni),
    .o(net5));
 b15bfn001as1n12x5 input6 (.a(tl_i[0]),
    .o(net6));
 b15bfn001as1n16x5 input7 (.a(tl_i[100]),
    .o(net7));
 b15bfn000as1n32x5 input8 (.a(tl_i[101]),
    .o(net8));
 b15bfn001as1n12x5 input9 (.a(tl_i[105]),
    .o(net9));
 b15bfn001ah1n16x5 input10 (.a(tl_i[106]),
    .o(net10));
 b15bfn001as1n12x5 input11 (.a(tl_i[107]),
    .o(net11));
 b15bfn001ah1n24x5 input12 (.a(tl_i[108]),
    .o(net12));
 b15bfn001as1n16x5 input13 (.a(tl_i[15]),
    .o(net13));
 b15bfn001as1n16x5 input14 (.a(tl_i[16]),
    .o(net14));
 b15bfn001as1n16x5 input15 (.a(tl_i[17]),
    .o(net15));
 b15bfn001as1n16x5 input16 (.a(tl_i[18]),
    .o(net16));
 b15bfn000as1n04x5 input17 (.a(tl_i[24]),
    .o(net17));
 b15bfn000as1n04x5 input18 (.a(tl_i[25]),
    .o(net18));
 b15bfn000as1n04x5 input19 (.a(tl_i[26]),
    .o(net19));
 b15bfn000as1n04x5 input20 (.a(tl_i[27]),
    .o(net20));
 b15bfm201as1n04x5 input21 (.a(tl_i[28]),
    .o(net21));
 b15qgbbf1an1n05x5 input22 (.a(tl_i[29]),
    .o(net22));
 b15bfn000ah1n04x5 input23 (.a(tl_i[30]),
    .o(net23));
 b15bfm201as1n04x5 input24 (.a(tl_i[31]),
    .o(net24));
 b15bfn001ah1n12x5 input25 (.a(tl_i[32]),
    .o(net25));
 b15bfn001ah1n12x5 input26 (.a(tl_i[33]),
    .o(net26));
 b15bfn001ah1n12x5 input27 (.a(tl_i[34]),
    .o(net27));
 b15bfn001ah1n12x5 input28 (.a(tl_i[35]),
    .o(net28));
 b15bfn001as1n12x5 input29 (.a(tl_i[36]),
    .o(net29));
 b15bfn001as1n12x5 input30 (.a(tl_i[37]),
    .o(net30));
 b15bfn001as1n12x5 input31 (.a(tl_i[38]),
    .o(net31));
 b15bfn001as1n12x5 input32 (.a(tl_i[39]),
    .o(net32));
 b15bfn001as1n12x5 input33 (.a(tl_i[40]),
    .o(net33));
 b15bfn001aq1n06x5 input34 (.a(tl_i[41]),
    .o(net34));
 b15bfn000ah1n06x5 input35 (.a(tl_i[42]),
    .o(net35));
 b15bfn001aq1n06x5 input36 (.a(tl_i[43]),
    .o(net36));
 b15bfn001ah1n08x5 input37 (.a(tl_i[44]),
    .o(net37));
 b15bfn001ah1n12x5 input38 (.a(tl_i[45]),
    .o(net38));
 b15bfn001ah1n12x5 input39 (.a(tl_i[46]),
    .o(net39));
 b15bfn001as1n08x5 input40 (.a(tl_i[47]),
    .o(net40));
 b15bfn001aq1n06x5 input41 (.a(tl_i[48]),
    .o(net41));
 b15bfn001aq1n06x5 input42 (.a(tl_i[49]),
    .o(net42));
 b15bfn001ah1n08x5 input43 (.a(tl_i[50]),
    .o(net43));
 b15bfn001as1n12x5 input44 (.a(tl_i[51]),
    .o(net44));
 b15bfn001ah1n12x5 input45 (.a(tl_i[52]),
    .o(net45));
 b15bfn001as1n12x5 input46 (.a(tl_i[53]),
    .o(net46));
 b15bfn001as1n08x5 input47 (.a(tl_i[54]),
    .o(net47));
 b15bfn001as1n08x5 input48 (.a(tl_i[55]),
    .o(net48));
 b15bfn001as1n32x5 input49 (.a(tl_i[56]),
    .o(net49));
 b15bfn001as1n32x5 input50 (.a(tl_i[57]),
    .o(net50));
 b15bfn001as1n32x5 input51 (.a(tl_i[58]),
    .o(net51));
 b15bfn001as1n32x5 input52 (.a(tl_i[59]),
    .o(net52));
 b15bfn001as1n16x5 input53 (.a(tl_i[60]),
    .o(net53));
 b15bfn001ah1n24x5 input54 (.a(tl_i[61]),
    .o(net54));
 b15bfn001as1n12x5 input55 (.a(tl_i[62]),
    .o(net55));
 b15bfn001as1n12x5 input56 (.a(tl_i[63]),
    .o(net56));
 b15bfn001as1n16x5 input57 (.a(tl_i[64]),
    .o(net57));
 b15bfn001ah1n16x5 input58 (.a(tl_i[65]),
    .o(net58));
 b15bfn001ah1n16x5 input59 (.a(tl_i[66]),
    .o(net59));
 b15bfn000ah1n04x5 input60 (.a(tl_i[67]),
    .o(net60));
 b15bfn001as1n24x5 input61 (.a(tl_i[68]),
    .o(net61));
 b15bfn001as1n08x5 input62 (.a(tl_i[69]),
    .o(net62));
 b15bfn000ah1n03x5 input63 (.a(tl_i[70]),
    .o(net63));
 b15bfn001as1n08x5 input64 (.a(tl_i[71]),
    .o(net64));
 b15bfn001ah1n32x5 input65 (.a(tl_i[72]),
    .o(net65));
 b15bfn001ah1n12x5 input66 (.a(tl_i[92]),
    .o(net66));
 b15bfn001ah1n12x5 input67 (.a(tl_i[93]),
    .o(net67));
 b15bfn001as1n12x5 input68 (.a(tl_i[94]),
    .o(net68));
 b15bfn001as1n12x5 input69 (.a(tl_i[95]),
    .o(net69));
 b15bfn001ah1n12x5 input70 (.a(tl_i[96]),
    .o(net70));
 b15bfn001ah1n12x5 input71 (.a(tl_i[97]),
    .o(net71));
 b15bfn001ah1n12x5 input72 (.a(tl_i[98]),
    .o(net72));
 b15bfn001ah1n12x5 input73 (.a(tl_i[99]),
    .o(net73));
 b15bfn000ah1n03x5 output74 (.a(net383),
    .o(net384));
 b15bfn000ah1n03x5 output75 (.a(net512),
    .o(tl_o[16]));
 b15bfn000ah1n03x5 output76 (.a(net434),
    .o(net435));
 b15bfn000ah1n03x5 output77 (.a(net505),
    .o(tl_o[18]));
 b15bfn000ah1n03x5 output78 (.a(net444),
    .o(net445));
 b15bfn000ah1n03x5 output79 (.a(net427),
    .o(net428));
 b15bfn000ah1n03x5 output80 (.a(net456),
    .o(net457));
 b15bfn000ah1n03x5 output81 (.a(net488),
    .o(net489));
 b15bfn000ah1n03x5 output82 (.a(net493),
    .o(tl_o[22]));
 b15bfn000ah1n03x5 output83 (.a(net462),
    .o(net463));
 b15bfn000ah1n03x5 output84 (.a(net478),
    .o(net479));
 b15bfn000ah1n03x5 output85 (.a(net439),
    .o(net440));
 b15bfn000ah1n03x5 output86 (.a(net564),
    .o(tl_o[26]));
 b15bfn000ah1n03x5 output87 (.a(net467),
    .o(net468));
 b15bfn000ah1n03x5 output88 (.a(net576),
    .o(tl_o[28]));
 b15bfn000ah1n03x5 output89 (.a(net579),
    .o(tl_o[29]));
 b15bfn000ah1n03x5 output90 (.a(net430),
    .o(tl_o[2]));
 b15bfn000ah1n03x5 output91 (.a(net508),
    .o(tl_o[30]));
 b15bfn000ah1n03x5 output92 (.a(net567),
    .o(tl_o[31]));
 b15bfn000ah1n03x5 output93 (.a(net546),
    .o(tl_o[32]));
 b15bfn000ah1n03x5 output94 (.a(net570),
    .o(tl_o[33]));
 b15bfn000ah1n03x5 output95 (.a(net537),
    .o(tl_o[34]));
 b15bfn000ah1n03x5 output96 (.a(net519),
    .o(tl_o[35]));
 b15bfn000ah1n03x5 output97 (.a(net573),
    .o(tl_o[36]));
 b15bfn000ah1n03x5 output98 (.a(net522),
    .o(tl_o[37]));
 b15bfn000ah1n03x5 output99 (.a(net582),
    .o(tl_o[38]));
 b15bfn000ah1n03x5 output100 (.a(net552),
    .o(tl_o[39]));
 b15bfn000ah1n03x5 output101 (.a(net415),
    .o(net416));
 b15bfn000ah1n03x5 output102 (.a(net534),
    .o(tl_o[40]));
 b15bfn000ah1n03x5 output103 (.a(net558),
    .o(tl_o[41]));
 b15bfn000ah1n03x5 output104 (.a(net549),
    .o(tl_o[42]));
 b15bfn000ah1n03x5 output105 (.a(net105),
    .o(tl_o[43]));
 b15bfn000ah1n03x5 output106 (.a(net472),
    .o(net473));
 b15bfn000ah1n03x5 output107 (.a(net498),
    .o(tl_o[45]));
 b15bfn000ah1n03x5 output108 (.a(net555),
    .o(tl_o[46]));
 b15bfn000ah1n03x5 output109 (.a(net501),
    .o(tl_o[47]));
 b15bfn000ah1n03x5 output110 (.a(net542),
    .o(net543));
 b15bfn000ah1n03x5 output111 (.a(net418),
    .o(net419));
 b15bfn000ah1n03x5 output112 (.a(net527),
    .o(net528));
 b15bfn000ah1n03x5 output113 (.a(net389),
    .o(net390));
 b15bfn000ah1n03x5 output114 (.a(net447),
    .o(net448));
 b15bfn000ah1n03x5 output115 (.a(net539),
    .o(net540));
 b15bfn000ah1n03x5 output116 (.a(net560),
    .o(net561));
 b15bfn000ah1n03x5 output117 (.a(net377),
    .o(net378));
 b15bfn000ah1n03x5 output118 (.a(net386),
    .o(net387));
 b15bfn000ah1n03x5 output119 (.a(net530),
    .o(net531));
 b15bfn000ah1n03x5 output120 (.a(net524),
    .o(net525));
 b15bfn000ah1n03x5 output121 (.a(net412),
    .o(net413));
 b15bfn000ah1n03x5 output122 (.a(net451),
    .o(net452));
 b15bfn000ah1n03x5 output123 (.a(net484),
    .o(tl_o[65]));
 b15bfn000ah1n03x5 output124 (.a(net403),
    .o(net404));
 b15bfn000ah1n03x5 output125 (.a(net396),
    .o(net397));
 b15bfn000ah1n03x5 output126 (.a(net421),
    .o(net422));
 b15bfn001ah1n48x5 fanout127 (.a(net487),
    .o(net127));
 b15bfn001as1n24x5 wire128 (.a(net127),
    .o(net128));
 b15bfn001as1n48x5 fanout129 (.a(net486),
    .o(net129));
 b15bfn001ah1n64x5 wire130 (.a(net129),
    .o(net130));
 b15bfn001as1n80x5 fanout131 (.a(net133),
    .o(net131));
 b15bfn001as1n64x5 fanout132 (.a(n383),
    .o(net132));
 b15bfn000as1n24x5 wire133 (.a(net132),
    .o(net133));
 b15bfn001as1n32x5 wire134 (.a(net132),
    .o(net134));
 b15bfn001as1n80x5 fanout135 (.a(net137),
    .o(net135));
 b15bfn001as1n64x5 fanout136 (.a(n381),
    .o(net136));
 b15bfn001ah1n32x5 wire137 (.a(net136),
    .o(net137));
 b15bfn001as1n32x5 wire138 (.a(net136),
    .o(net138));
 b15bfn001as1n32x5 wire139 (.a(n376),
    .o(net139));
 b15bfn001ah1n24x5 wire140 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .o(net140));
 b15bfn001ah1n48x5 wire141 (.a(u_tlul_adapter_sram_rdata_tlword[19]),
    .o(net141));
 b15bfn001ah1n48x5 wire142 (.a(u_tlul_adapter_sram_rdata_tlword[18]),
    .o(net142));
 b15bfn001ah1n48x5 wire143 (.a(u_tlul_adapter_sram_rdata_tlword[17]),
    .o(net143));
 b15bfn001as1n32x5 wire144 (.a(u_tlul_adapter_sram_rdata_tlword[16]),
    .o(net144));
 b15bfn001as1n24x5 wire145 (.a(u_tlul_adapter_sram_rdata_tlword[13]),
    .o(net145));
 b15bfn001as1n24x5 wire146 (.a(u_tlul_adapter_sram_rdata_tlword[10]),
    .o(net146));
 b15bfn001as1n48x5 wire147 (.a(u_tlul_adapter_sram_rdata_tlword[22]),
    .o(net147));
 b15bfn001ah1n48x5 wire148 (.a(u_tlul_adapter_sram_rdata_tlword[21]),
    .o(net148));
 b15bfn001ah1n48x5 wire149 (.a(u_tlul_adapter_sram_rdata_tlword[20]),
    .o(net149));
 b15bfn001as1n24x5 wire150 (.a(u_tlul_adapter_sram_rdata_tlword[25]),
    .o(net150));
 b15bfn001ah1n24x5 wire151 (.a(n434),
    .o(net151));
 b15bfn001ah1n48x5 max_length152 (.a(n434),
    .o(net152));
 b15bfn001ah1n48x5 wire153 (.a(net495),
    .o(net153));
 b15bfn001ah1n24x5 wire154 (.a(wdata[16]),
    .o(net154));
 b15bfn001as1n48x5 wire155 (.a(n418),
    .o(net155));
 b15bfn001ah1n32x5 wire156 (.a(n325),
    .o(net156));
 b15bfn001as1n16x5 wire157 (.a(n_0_net_),
    .o(net157));
 b15bfn001ah1n16x5 wire158 (.a(net431),
    .o(net158));
 b15bfn001as1n16x5 wire159 (.a(net509),
    .o(net159));
 b15bfn001ah1n16x5 wire160 (.a(net469),
    .o(net160));
 b15bfn001ah1n16x5 wire161 (.a(net513),
    .o(net161));
 b15bfn001as1n16x5 wire162 (.a(net516),
    .o(net162));
 b15bfn001as1n16x5 wire163 (.a(net464),
    .o(net163));
 b15bfn001as1n16x5 wire164 (.a(net436),
    .o(net164));
 b15bfn001ah1n24x5 wire165 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[16]),
    .o(net165));
 b15bfn001ah1n24x5 wire166 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[15]),
    .o(net166));
 b15bfn001ah1n24x5 wire167 (.a(net490),
    .o(net167));
 b15bfn001ah1n16x5 wire168 (.a(net453),
    .o(net168));
 b15bfn001ah1n16x5 wire169 (.a(net441),
    .o(net169));
 b15bfn001as1n16x5 wire170 (.a(net502),
    .o(net170));
 b15bfn001ah1n24x5 wire171 (.a(net424),
    .o(net171));
 b15bfn001ah1n12x5 wire172 (.a(net423),
    .o(net172));
 b15bfn001ah1n16x5 wire173 (.a(net398),
    .o(net173));
 b15bfn001ah1n48x5 wire174 (.a(wen),
    .o(net174));
 b15bfn001as1n16x5 wire175 (.a(addr[9]),
    .o(net175));
 b15bfn001as1n16x5 wire176 (.a(addr[10]),
    .o(net176));
 b15bfn001ah1n24x5 wire177 (.a(addr[2]),
    .o(net177));
 b15bfn001ah1n24x5 wire178 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst),
    .o(net178));
 b15bfn001as1n16x5 wire179 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_wptr_value_0_),
    .o(net179));
 b15bfn001as1n16x5 wire180 (.a(net379),
    .o(net180));
 b15bfn001ah1n16x5 wire181 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[3]),
    .o(net181));
 b15bfn001ah1n16x5 wire182 (.a(net391),
    .o(net182));
 b15bfn000ah1n24x5 wire183 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_wptr_value_0_),
    .o(net183));
 b15bfn001as1n16x5 wire184 (.a(net405),
    .o(net184));
 b15bfn001as1n16x5 wire185 (.a(net480),
    .o(net185));
 b15bfn001ah1n48x5 wire186 (.a(n328),
    .o(net186));
 b15bfn001as1n64x5 wire187 (.a(net188),
    .o(net187));
 b15bfn001as1n24x5 max_length188 (.a(n328),
    .o(net188));
 b15bfn001as1n32x5 wire189 (.a(net7),
    .o(net189));
 b15bfn001as1n32x5 wire190 (.a(net65),
    .o(net190));
 b15bfn001as1n24x5 wire191 (.a(net61),
    .o(net191));
 b15bfn001as1n32x5 wire192 (.a(net53),
    .o(net192));
 b15bfn001as1n24x5 wire193 (.a(net52),
    .o(net193));
 b15bfn000as1n32x5 wire194 (.a(net51),
    .o(net194));
 b15bfn001as1n32x5 wire195 (.a(net50),
    .o(net195));
 b15bfn001as1n32x5 wire196 (.a(net50),
    .o(net196));
 b15bfn001ah1n48x5 wire197 (.a(net5),
    .o(net197));
 b15bfn001as1n32x5 wire198 (.a(net49),
    .o(net198));
 b15bfn001ah1n32x5 wire199 (.a(net49),
    .o(net199));
 b15bfn001ah1n24x5 wire200 (.a(net33),
    .o(net200));
 b15bfn001ah1n32x5 wire201 (.a(rdata[31]),
    .o(net201));
 b15bfn001ah1n24x5 wire202 (.a(rdata[29]),
    .o(net202));
 b15bfn001ah1n24x5 wire203 (.a(rdata[22]),
    .o(net203));
 b15bfn001as1n16x5 wire204 (.a(rdata[21]),
    .o(net204));
 b15bfn001ah1n24x5 wire205 (.a(rdata[18]),
    .o(net205));
 b15bfn001ah1n24x5 wire206 (.a(rdata[17]),
    .o(net206));
 b15bfn001ah1n24x5 wire207 (.a(rdata[16]),
    .o(net207));
 b15tilo00an1n03x5 rvalid_reg_u_tlul_adapter_sram_intg_error_q_reg_208 (.o(net208));
 b15tilo00an1n03x5 rvalid_reg_u_tlul_adapter_sram_intg_error_q_reg_209 (.o(net209));
 b15tilo00an1n03x5 u_sram_210 (.o(net210));
 b15tilo00an1n03x5 u_sram_211 (.o(net211));
 b15tilo00an1n03x5 u_sram_212 (.o(net212));
 b15tilo00an1n03x5 u_sram_213 (.o(net213));
 b15tilo00an1n03x5 u_sram_214 (.o(net214));
 b15tilo00an1n03x5 u_sram_215 (.o(net215));
 b15tilo00an1n03x5 u_sram_216 (.o(net216));
 b15tilo00an1n03x5 u_sram_217 (.o(net217));
 b15tilo00an1n03x5 u_sram_218 (.o(net218));
 b15tilo00an1n03x5 u_sram_219 (.o(net219));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_clk_gate_gen_normal_fifo_storage_reg_0__0_latch_220 (.o(net220));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_clk_gate_gen_normal_fifo_storage_reg_0__latch_221 (.o(net221));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__1__222 (.o(net222));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__1__223 (.o(net223));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__11__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__12__224 (.o(net224));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__11__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__12__225 (.o(net225));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__13__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__14__226 (.o(net226));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__13__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__14__227 (.o(net227));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__15__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__16__228 (.o(net228));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__15__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__16__229 (.o(net229));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__15__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__16__230 (.o(net230));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__3__231 (.o(net231));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__3__232 (.o(net232));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__5__233 (.o(net233));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__5__234 (.o(net234));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__7__235 (.o(net235));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__7__236 (.o(net236));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__8__237 (.o(net237));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__9__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__10__238 (.o(net238));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__9__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__10__239 (.o(net239));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__240 (.o(net240));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__241 (.o(net241));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__242 (.o(net242));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__243 (.o(net243));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst_reg_244 (.o(net244));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst_reg_245 (.o(net245));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_clk_gate_gen_normal_fifo_storage_reg_0__0_latch_246 (.o(net246));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_clk_gate_gen_normal_fifo_storage_reg_0__latch_247 (.o(net247));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1__248 (.o(net248));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1__249 (.o(net249));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1__250 (.o(net250));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1__251 (.o(net251));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__10__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__11__252 (.o(net252));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__10__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__11__253 (.o(net253));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__12__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__13__254 (.o(net254));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__12__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__13__255 (.o(net255));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__14__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__15__256 (.o(net256));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__14__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__15__257 (.o(net257));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__16__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__17__258 (.o(net258));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__16__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__17__259 (.o(net259));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__18__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__19__260 (.o(net260));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__18__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__19__261 (.o(net261));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__20__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__21__262 (.o(net262));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__20__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__21__263 (.o(net263));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__22__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__23__264 (.o(net264));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__22__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__23__265 (.o(net265));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__24__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__25__266 (.o(net266));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__24__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__25__267 (.o(net267));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__26__268 (.o(net268));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__27__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__28__269 (.o(net269));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__27__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__28__270 (.o(net270));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__29__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__30__271 (.o(net271));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__29__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__30__272 (.o(net272));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3__273 (.o(net273));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3__274 (.o(net274));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3__275 (.o(net275));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3__276 (.o(net276));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__31__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__32__277 (.o(net277));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__31__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__32__278 (.o(net278));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__33__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__34__279 (.o(net279));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__33__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__34__280 (.o(net280));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__35__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__36__281 (.o(net281));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__35__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__36__282 (.o(net282));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__37__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__38__283 (.o(net283));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__37__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__38__284 (.o(net284));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__39__285 (.o(net285));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5__286 (.o(net286));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5__287 (.o(net287));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5__288 (.o(net288));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5__289 (.o(net289));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7__290 (.o(net290));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7__291 (.o(net291));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7__292 (.o(net292));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7__293 (.o(net293));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__8__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__9__294 (.o(net294));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__8__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__9__295 (.o(net295));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__296 (.o(net296));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__297 (.o(net297));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__298 (.o(net298));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__299 (.o(net299));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst_reg_300 (.o(net300));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst_reg_301 (.o(net301));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__0__302 (.o(net302));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__1__303 (.o(net303));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__2__304 (.o(net304));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__3__305 (.o(net305));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__4__306 (.o(net306));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__307 (.o(net307));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__308 (.o(net308));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__309 (.o(net309));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__310 (.o(net310));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst_reg_311 (.o(net311));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst_reg_312 (.o(net312));
 b15tihi00an1n03x5 U588_314 (.o(net314));
 b15tihi00an1n03x5 U594_315 (.o(net315));
 b15tihi00an1n03x5 U602_316 (.o(net316));
 b15tihi00an1n03x5 U622_317 (.o(net317));
 b15tihi00an1n03x5 U637_318 (.o(net318));
 b15tihi00an1n03x5 U702_319 (.o(net319));
 b15tihi00an1n03x5 U704_320 (.o(net320));
 b15tihi00an1n03x5 U706_321 (.o(net321));
 b15tihi00an1n03x5 U708_322 (.o(net322));
 b15tihi00an1n03x5 U710_323 (.o(net323));
 b15tihi00an1n03x5 U712_324 (.o(net324));
 b15tihi00an1n03x5 U714_325 (.o(net325));
 b15tihi00an1n03x5 rvalid_reg_u_tlul_adapter_sram_intg_error_q_reg_326 (.o(net326));
 b15tihi00an1n03x5 u_sram_327 (.o(net327));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__1__328 (.o(net328));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__11__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__12__329 (.o(net329));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__13__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__14__330 (.o(net330));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__15__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__16__331 (.o(net331));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__3__332 (.o(net332));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__5__333 (.o(net333));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__7__334 (.o(net334));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__8__335 (.o(net335));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__9__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__10__336 (.o(net336));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__337 (.o(net337));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__338 (.o(net338));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__339 (.o(net339));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst_reg_340 (.o(net340));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1__341 (.o(net341));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__10__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__11__342 (.o(net342));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__12__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__13__343 (.o(net343));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__14__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__15__344 (.o(net344));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__16__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__17__345 (.o(net345));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__18__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__19__346 (.o(net346));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__20__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__21__347 (.o(net347));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__22__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__23__348 (.o(net348));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__24__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__25__349 (.o(net349));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__26__350 (.o(net350));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__27__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__28__351 (.o(net351));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__29__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__30__352 (.o(net352));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3__353 (.o(net353));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__31__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__32__354 (.o(net354));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__33__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__34__355 (.o(net355));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__35__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__36__356 (.o(net356));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__37__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__38__357 (.o(net357));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__39__358 (.o(net358));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5__359 (.o(net359));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7__360 (.o(net360));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__8__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__9__361 (.o(net361));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__362 (.o(net362));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__363 (.o(net363));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__364 (.o(net364));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst_reg_365 (.o(net365));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__0__366 (.o(net366));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__1__367 (.o(net367));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__2__368 (.o(net368));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__3__369 (.o(net369));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__4__370 (.o(net370));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__371 (.o(net371));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__372 (.o(net372));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__373 (.o(net373));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst_reg_374 (.o(net374));
 b15cbf000an1n16x5 clkbuf_1_0__f_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_1_0__leaf_clk_i));
 b15cbf000an1n16x5 clkbuf_1_1__f_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_1_1__leaf_clk_i));
 b15cbf000an1n16x5 clkbuf_0_u_tlul_adapter_sram_u_rspfifo_net616 (.clk(u_tlul_adapter_sram_u_rspfifo_net616),
    .clkout(clknet_0_u_tlul_adapter_sram_u_rspfifo_net616));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_tlul_adapter_sram_u_rspfifo_net616 (.clk(clknet_0_u_tlul_adapter_sram_u_rspfifo_net616),
    .clkout(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net616));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_tlul_adapter_sram_u_rspfifo_net616 (.clk(clknet_0_u_tlul_adapter_sram_u_rspfifo_net616),
    .clkout(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net616));
 b15cbf000an1n16x5 clkbuf_0_u_tlul_adapter_sram_u_rspfifo_net622 (.clk(u_tlul_adapter_sram_u_rspfifo_net622),
    .clkout(clknet_0_u_tlul_adapter_sram_u_rspfifo_net622));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_tlul_adapter_sram_u_rspfifo_net622 (.clk(clknet_0_u_tlul_adapter_sram_u_rspfifo_net622),
    .clkout(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_tlul_adapter_sram_u_rspfifo_net622 (.clk(clknet_0_u_tlul_adapter_sram_u_rspfifo_net622),
    .clkout(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622));
 b15cbf000an1n16x5 clkbuf_0_u_tlul_adapter_sram_u_reqfifo_net644 (.clk(u_tlul_adapter_sram_u_reqfifo_net644),
    .clkout(clknet_0_u_tlul_adapter_sram_u_reqfifo_net644));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_tlul_adapter_sram_u_reqfifo_net644 (.clk(clknet_0_u_tlul_adapter_sram_u_reqfifo_net644),
    .clkout(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net644));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_tlul_adapter_sram_u_reqfifo_net644 (.clk(clknet_0_u_tlul_adapter_sram_u_reqfifo_net644),
    .clkout(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net644));
 b15cbf000an1n16x5 clkbuf_0_u_tlul_adapter_sram_u_reqfifo_net650 (.clk(u_tlul_adapter_sram_u_reqfifo_net650),
    .clkout(clknet_0_u_tlul_adapter_sram_u_reqfifo_net650));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_tlul_adapter_sram_u_reqfifo_net650 (.clk(clknet_0_u_tlul_adapter_sram_u_reqfifo_net650),
    .clkout(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net650));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_tlul_adapter_sram_u_reqfifo_net650 (.clk(clknet_0_u_tlul_adapter_sram_u_reqfifo_net650),
    .clkout(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net650));
 b15bfn001as1n16x5 wire1 (.a(clk_i),
    .o(net375));
 b15cbf034ar1n64x5 hold2 (.clk(net586),
    .clkout(net376));
 b15cbf034ar1n64x5 hold3 (.clk(net117),
    .clkout(net377));
 b15cbf034ar1n64x5 hold4 (.clk(net378),
    .clkout(tl_o[55]));
 b15cbf034ar1n64x5 hold5 (.clk(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_rptr_value_0_),
    .clkout(net379));
 b15cbf034ar1n64x5 hold6 (.clk(net180),
    .clkout(net380));
 b15cbf034ar1n64x5 hold7 (.clk(n359),
    .clkout(net381));
 b15cbf034ar1n64x5 hold8 (.clk(n362),
    .clkout(net382));
 b15cbf034ar1n64x5 hold9 (.clk(net74),
    .clkout(net383));
 b15cbf034ar1n64x5 hold10 (.clk(net384),
    .clkout(tl_o[0]));
 b15cbf034ar1n64x5 hold11 (.clk(net587),
    .clkout(net385));
 b15cbf034ar1n64x5 hold12 (.clk(net118),
    .clkout(net386));
 b15cbf034ar1n64x5 hold13 (.clk(net387),
    .clkout(tl_o[56]));
 b15cbf034ar1n64x5 hold14 (.clk(net588),
    .clkout(net388));
 b15cbf034ar1n64x5 hold15 (.clk(net113),
    .clkout(net389));
 b15cbf034ar1n64x5 hold16 (.clk(net390),
    .clkout(tl_o[51]));
 b15cbf034ar1n64x5 hold17 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_rptr_value_0_),
    .clkout(net391));
 b15cbf034ar1n64x5 hold18 (.clk(net182),
    .clkout(net392));
 b15cbf034ar1n64x5 hold19 (.clk(n368),
    .clkout(net393));
 b15cbf034ar1n64x5 hold20 (.clk(n380),
    .clkout(net394));
 b15cbf034ar1n64x5 hold21 (.clk(n386),
    .clkout(net395));
 b15cbf034ar1n64x5 hold22 (.clk(net125),
    .clkout(net396));
 b15cbf034ar1n64x5 hold23 (.clk(net397),
    .clkout(tl_o[7]));
 b15cbf034ar1n64x5 hold24 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[14]),
    .clkout(net398));
 b15cbf034ar1n64x5 hold25 (.clk(net173),
    .clkout(net399));
 b15cbf034ar1n64x5 hold26 (.clk(net410),
    .clkout(net400));
 b15cbf034ar1n64x5 hold27 (.clk(n382),
    .clkout(net401));
 b15cbf034ar1n64x5 hold28 (.clk(n371),
    .clkout(net402));
 b15cbf034ar1n64x5 hold29 (.clk(net124),
    .clkout(net403));
 b15cbf034ar1n64x5 hold30 (.clk(net404),
    .clkout(tl_o[6]));
 b15cbf034ar1n64x5 hold31 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_rptr_value_0_),
    .clkout(net405));
 b15cbf034ar1n64x5 hold32 (.clk(net184),
    .clkout(net406));
 b15cbf034ar1n64x5 hold33 (.clk(n358),
    .clkout(net407));
 b15cbf034ar1n64x5 hold34 (.clk(n384),
    .clkout(net408));
 b15cbf034ar1n64x5 hold35 (.clk(n374),
    .clkout(net409));
 b15cbf034ar1n64x5 hold36 (.clk(n385),
    .clkout(net410));
 b15cbf034ar1n64x5 hold37 (.clk(net400),
    .clkout(net411));
 b15cbf034ar1n64x5 hold38 (.clk(net121),
    .clkout(net412));
 b15cbf034ar1n64x5 hold39 (.clk(net413),
    .clkout(tl_o[5]));
 b15cbf034ar1n64x5 hold40 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[2]),
    .clkout(net414));
 b15cbf034ar1n64x5 hold41 (.clk(net101),
    .clkout(net415));
 b15cbf034ar1n64x5 hold42 (.clk(net416),
    .clkout(tl_o[3]));
 b15cbf034ar1n64x5 hold43 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[3]),
    .clkout(net417));
 b15cbf034ar1n64x5 hold44 (.clk(net111),
    .clkout(net418));
 b15cbf034ar1n64x5 hold45 (.clk(net419),
    .clkout(tl_o[4]));
 b15cbf034ar1n64x5 hold46 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[7]),
    .clkout(net420));
 b15cbf034ar1n64x5 hold47 (.clk(net126),
    .clkout(net421));
 b15cbf034ar1n64x5 hold48 (.clk(net422),
    .clkout(tl_o[8]));
 b15cbf034ar1n64x5 hold49 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[0]),
    .clkout(net423));
 b15cbf034ar1n64x5 hold50 (.clk(net172),
    .clkout(net424));
 b15cbf034ar1n64x5 hold51 (.clk(net171),
    .clkout(net425));
 b15cbf034ar1n64x5 hold52 (.clk(n378),
    .clkout(net426));
 b15cbf034ar1n64x5 hold53 (.clk(net79),
    .clkout(net427));
 b15cbf034ar1n64x5 hold54 (.clk(net428),
    .clkout(tl_o[1]));
 b15cbf034ar1n64x5 hold55 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[1]),
    .clkout(net429));
 b15cbf034ar1n64x5 hold56 (.clk(net90),
    .clkout(net430));
 b15cbf034ar1n64x5 hold57 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[9]),
    .clkout(net431));
 b15cbf034ar1n64x5 hold58 (.clk(net158),
    .clkout(net432));
 b15cbf034ar1n64x5 hold59 (.clk(n410),
    .clkout(net433));
 b15cbf034ar1n64x5 hold60 (.clk(net76),
    .clkout(net434));
 b15cbf034ar1n64x5 hold61 (.clk(net435),
    .clkout(tl_o[17]));
 b15cbf034ar1n64x5 hold62 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[17]),
    .clkout(net436));
 b15cbf034ar1n64x5 hold63 (.clk(net164),
    .clkout(net437));
 b15cbf034ar1n64x5 hold64 (.clk(n420),
    .clkout(net438));
 b15cbf034ar1n64x5 hold65 (.clk(net85),
    .clkout(net439));
 b15cbf034ar1n64x5 hold66 (.clk(net440),
    .clkout(tl_o[25]));
 b15cbf034ar1n64x5 hold67 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[11]),
    .clkout(net441));
 b15cbf034ar1n64x5 hold68 (.clk(net169),
    .clkout(net442));
 b15cbf034ar1n64x5 hold69 (.clk(n412),
    .clkout(net443));
 b15cbf034ar1n64x5 hold70 (.clk(net78),
    .clkout(net444));
 b15cbf034ar1n64x5 hold71 (.clk(net445),
    .clkout(tl_o[19]));
 b15cbf034ar1n64x5 hold72 (.clk(net589),
    .clkout(net446));
 b15cbf034ar1n64x5 hold73 (.clk(net114),
    .clkout(net447));
 b15cbf034ar1n64x5 hold74 (.clk(net448),
    .clkout(tl_o[52]));
 b15cbf034ar1n64x5 hold75 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[15]),
    .clkout(net449));
 b15cbf034ar1n64x5 hold76 (.clk(n379),
    .clkout(net450));
 b15cbf034ar1n64x5 hold77 (.clk(net122),
    .clkout(net451));
 b15cbf034ar1n64x5 hold78 (.clk(net452),
    .clkout(tl_o[62]));
 b15cbf034ar1n64x5 hold79 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[12]),
    .clkout(net453));
 b15cbf034ar1n64x5 hold80 (.clk(net168),
    .clkout(net454));
 b15cbf034ar1n64x5 hold81 (.clk(n413),
    .clkout(net455));
 b15cbf034ar1n64x5 hold82 (.clk(net80),
    .clkout(net456));
 b15cbf034ar1n64x5 hold83 (.clk(net457),
    .clkout(tl_o[20]));
 b15cbf034ar1n64x5 hold84 (.clk(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[1]),
    .clkout(net458));
 b15cbf034ar1n64x5 hold85 (.clk(n416),
    .clkout(net459));
 b15cbf034ar1n64x5 hold86 (.clk(u_tlul_adapter_sram_rdata_tlword[7]),
    .clkout(net460));
 b15cbf034ar1n64x5 hold87 (.clk(n417),
    .clkout(net461));
 b15cbf034ar1n64x5 hold88 (.clk(net83),
    .clkout(net462));
 b15cbf034ar1n64x5 hold89 (.clk(net463),
    .clkout(tl_o[23]));
 b15cbf034ar1n64x5 hold90 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[19]),
    .clkout(net464));
 b15cbf034ar1n64x5 hold91 (.clk(net163),
    .clkout(net465));
 b15cbf034ar1n64x5 hold92 (.clk(n424),
    .clkout(net466));
 b15cbf034ar1n64x5 hold93 (.clk(net87),
    .clkout(net467));
 b15cbf034ar1n64x5 hold94 (.clk(net468),
    .clkout(tl_o[27]));
 b15cbf034ar1n64x5 hold95 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[36]),
    .clkout(net469));
 b15cbf034ar1n64x5 hold96 (.clk(net160),
    .clkout(net470));
 b15cbf034ar1n64x5 hold97 (.clk(n396),
    .clkout(net471));
 b15cbf034ar1n64x5 hold98 (.clk(net106),
    .clkout(net472));
 b15cbf034ar1n64x5 hold99 (.clk(net473),
    .clkout(tl_o[44]));
 b15cbf034ar1n64x5 hold100 (.clk(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[2]),
    .clkout(net474));
 b15cbf034ar1n64x5 hold101 (.clk(n429),
    .clkout(net475));
 b15cbf034ar1n64x5 hold102 (.clk(u_tlul_adapter_sram_rdata_tlword[8]),
    .clkout(net476));
 b15cbf034ar1n64x5 hold103 (.clk(n419),
    .clkout(net477));
 b15cbf034ar1n64x5 hold104 (.clk(net84),
    .clkout(net478));
 b15cbf034ar1n64x5 hold105 (.clk(net479),
    .clkout(tl_o[24]));
 b15cbf034ar1n64x5 hold106 (.clk(rvalid),
    .clkout(net480));
 b15cbf034ar1n64x5 hold107 (.clk(net185),
    .clkout(net481));
 b15cbf034ar1n64x5 hold108 (.clk(n369),
    .clkout(net482));
 b15cbf034ar1n64x5 hold109 (.clk(n375),
    .clkout(net483));
 b15cbf034ar1n64x5 hold110 (.clk(net123),
    .clkout(net484));
 b15cbf034ar1n64x5 hold111 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[10]),
    .clkout(net485));
 b15cbf034ar1n64x5 hold112 (.clk(n389),
    .clkout(net486));
 b15cbf034ar1n64x5 hold113 (.clk(net129),
    .clkout(net487));
 b15cbf034ar1n64x5 hold114 (.clk(net81),
    .clkout(net488));
 b15cbf034ar1n64x5 hold115 (.clk(net489),
    .clkout(tl_o[21]));
 b15cbf034ar1n64x5 hold116 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[14]),
    .clkout(net490));
 b15cbf034ar1n64x5 hold117 (.clk(net167),
    .clkout(net491));
 b15cbf034ar1n64x5 hold118 (.clk(n415),
    .clkout(net492));
 b15cbf034ar1n64x5 hold119 (.clk(net82),
    .clkout(net493));
 b15cbf034ar1n64x5 hold120 (.clk(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[4]),
    .clkout(net494));
 b15cbf034ar1n64x5 hold121 (.clk(n397),
    .clkout(net495));
 b15cbf034ar1n64x5 hold122 (.clk(u_tlul_adapter_sram_rdata_tlword[29]),
    .clkout(net496));
 b15cbf034ar1n64x5 hold123 (.clk(n401),
    .clkout(net497));
 b15cbf034ar1n64x5 hold124 (.clk(net107),
    .clkout(net498));
 b15cbf034ar1n64x5 hold125 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[39]),
    .clkout(net499));
 b15cbf034ar1n64x5 hold126 (.clk(n395),
    .clkout(net500));
 b15cbf034ar1n64x5 hold127 (.clk(net109),
    .clkout(net501));
 b15cbf034ar1n64x5 hold128 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[10]),
    .clkout(net502));
 b15cbf034ar1n64x5 hold129 (.clk(net170),
    .clkout(net503));
 b15cbf034ar1n64x5 hold130 (.clk(n411),
    .clkout(net504));
 b15cbf034ar1n64x5 hold131 (.clk(net77),
    .clkout(net505));
 b15cbf034ar1n64x5 hold132 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[22]),
    .clkout(net506));
 b15cbf034ar1n64x5 hold133 (.clk(n428),
    .clkout(net507));
 b15cbf034ar1n64x5 hold134 (.clk(net91),
    .clkout(net508));
 b15cbf034ar1n64x5 hold135 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[8]),
    .clkout(net509));
 b15cbf034ar1n64x5 hold136 (.clk(net159),
    .clkout(net510));
 b15cbf034ar1n64x5 hold137 (.clk(n409),
    .clkout(net511));
 b15cbf034ar1n64x5 hold138 (.clk(net75),
    .clkout(net512));
 b15cbf034ar1n64x5 hold139 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[35]),
    .clkout(net513));
 b15cbf034ar1n64x5 hold140 (.clk(net161),
    .clkout(net514));
 b15cbf034ar1n64x5 hold141 (.clk(n391),
    .clkout(net515));
 b15cbf034ar1n64x5 hold142 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[27]),
    .clkout(net516));
 b15cbf034ar1n64x5 hold143 (.clk(net162),
    .clkout(net517));
 b15cbf034ar1n64x5 hold144 (.clk(n438),
    .clkout(net518));
 b15cbf034ar1n64x5 hold145 (.clk(net96),
    .clkout(net519));
 b15cbf034ar1n64x5 hold146 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[29]),
    .clkout(net520));
 b15cbf034ar1n64x5 hold147 (.clk(n403),
    .clkout(net521));
 b15cbf034ar1n64x5 hold148 (.clk(net98),
    .clkout(net522));
 b15cbf034ar1n64x5 hold149 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[9]),
    .clkout(net523));
 b15cbf034ar1n64x5 hold150 (.clk(net120),
    .clkout(net524));
 b15cbf034ar1n64x5 hold151 (.clk(net525),
    .clkout(tl_o[58]));
 b15cbf034ar1n64x5 hold152 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[1]),
    .clkout(net526));
 b15cbf034ar1n64x5 hold153 (.clk(net112),
    .clkout(net527));
 b15cbf034ar1n64x5 hold154 (.clk(net528),
    .clkout(tl_o[50]));
 b15cbf034ar1n64x5 hold155 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[8]),
    .clkout(net529));
 b15cbf034ar1n64x5 hold156 (.clk(net119),
    .clkout(net530));
 b15cbf034ar1n64x5 hold157 (.clk(net531),
    .clkout(tl_o[57]));
 b15cbf034ar1n64x5 hold158 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[32]),
    .clkout(net532));
 b15cbf034ar1n64x5 hold159 (.clk(n392),
    .clkout(net533));
 b15cbf034ar1n64x5 hold160 (.clk(net102),
    .clkout(net534));
 b15cbf034ar1n64x5 hold161 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[26]),
    .clkout(net535));
 b15cbf034ar1n64x5 hold162 (.clk(n433),
    .clkout(net536));
 b15cbf034ar1n64x5 hold163 (.clk(net95),
    .clkout(net537));
 b15cbf034ar1n64x5 hold164 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[4]),
    .clkout(net538));
 b15cbf034ar1n64x5 hold165 (.clk(net115),
    .clkout(net539));
 b15cbf034ar1n64x5 hold166 (.clk(net540),
    .clkout(tl_o[53]));
 b15cbf034ar1n64x5 hold167 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[0]),
    .clkout(net541));
 b15cbf034ar1n64x5 hold168 (.clk(net110),
    .clkout(net542));
 b15cbf034ar1n64x5 hold169 (.clk(net543),
    .clkout(tl_o[49]));
 b15cbf034ar1n64x5 hold170 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[24]),
    .clkout(net544));
 b15cbf034ar1n64x5 hold171 (.clk(n431),
    .clkout(net545));
 b15cbf034ar1n64x5 hold172 (.clk(net93),
    .clkout(net546));
 b15cbf034ar1n64x5 hold173 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[34]),
    .clkout(net547));
 b15cbf034ar1n64x5 hold174 (.clk(n390),
    .clkout(net548));
 b15cbf034ar1n64x5 hold175 (.clk(net104),
    .clkout(net549));
 b15cbf034ar1n64x5 hold176 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[31]),
    .clkout(net550));
 b15cbf034ar1n64x5 hold177 (.clk(n405),
    .clkout(net551));
 b15cbf034ar1n64x5 hold178 (.clk(net100),
    .clkout(net552));
 b15cbf034ar1n64x5 hold179 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[38]),
    .clkout(net553));
 b15cbf034ar1n64x5 hold180 (.clk(n394),
    .clkout(net554));
 b15cbf034ar1n64x5 hold181 (.clk(net108),
    .clkout(net555));
 b15cbf034ar1n64x5 hold182 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[33]),
    .clkout(net556));
 b15cbf034ar1n64x5 hold183 (.clk(n393),
    .clkout(net557));
 b15cbf034ar1n64x5 hold184 (.clk(net103),
    .clkout(net558));
 b15cbf034ar1n64x5 hold185 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[5]),
    .clkout(net559));
 b15cbf034ar1n64x5 hold186 (.clk(net116),
    .clkout(net560));
 b15cbf034ar1n64x5 hold187 (.clk(net561),
    .clkout(tl_o[54]));
 b15cbf034ar1n64x5 hold188 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[18]),
    .clkout(net562));
 b15cbf034ar1n64x5 hold189 (.clk(n421),
    .clkout(net563));
 b15cbf034ar1n64x5 hold190 (.clk(net86),
    .clkout(net564));
 b15cbf034ar1n64x5 hold191 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[23]),
    .clkout(net565));
 b15cbf034ar1n64x5 hold192 (.clk(n430),
    .clkout(net566));
 b15cbf034ar1n64x5 hold193 (.clk(net92),
    .clkout(net567));
 b15cbf034ar1n64x5 hold194 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[25]),
    .clkout(net568));
 b15cbf034ar1n64x5 hold195 (.clk(n432),
    .clkout(net569));
 b15cbf034ar1n64x5 hold196 (.clk(net94),
    .clkout(net570));
 b15cbf034ar1n64x5 hold197 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[28]),
    .clkout(net571));
 b15cbf034ar1n64x5 hold198 (.clk(n402),
    .clkout(net572));
 b15cbf034ar1n64x5 hold199 (.clk(net97),
    .clkout(net573));
 b15cbf034ar1n64x5 hold200 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[20]),
    .clkout(net574));
 b15cbf034ar1n64x5 hold201 (.clk(n426),
    .clkout(net575));
 b15cbf034ar1n64x5 hold202 (.clk(net88),
    .clkout(net576));
 b15cbf034ar1n64x5 hold203 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[21]),
    .clkout(net577));
 b15cbf034ar1n64x5 hold204 (.clk(n427),
    .clkout(net578));
 b15cbf034ar1n64x5 hold205 (.clk(net89),
    .clkout(net579));
 b15cbf034ar1n64x5 hold206 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[30]),
    .clkout(net580));
 b15cbf034ar1n64x5 hold207 (.clk(n404),
    .clkout(net581));
 b15cbf034ar1n64x5 hold208 (.clk(net99),
    .clkout(net582));
 b15cbf034ar1n64x5 hold209 (.clk(n211),
    .clkout(net583));
 b15cbf034ar1n64x5 hold210 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_wptr_1_),
    .clkout(net584));
 b15cbf034ar1n64x5 hold211 (.clk(n357),
    .clkout(net585));
 b15cbf034ar1n64x5 hold212 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[6]),
    .clkout(net586));
 b15cbf034ar1n64x5 hold213 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[7]),
    .clkout(net587));
 b15cbf034ar1n64x5 hold214 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[2]),
    .clkout(net588));
 b15cbf034ar1n64x5 hold215 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[3]),
    .clkout(net589));
 b15zdnd11an1n64x5 FILLER_0_8 ();
 b15zdnd11an1n64x5 FILLER_0_72 ();
 b15zdnd11an1n64x5 FILLER_0_136 ();
 b15zdnd11an1n64x5 FILLER_0_200 ();
 b15zdnd11an1n64x5 FILLER_0_264 ();
 b15zdnd11an1n64x5 FILLER_0_328 ();
 b15zdnd11an1n64x5 FILLER_0_392 ();
 b15zdnd11an1n64x5 FILLER_0_456 ();
 b15zdnd11an1n64x5 FILLER_0_520 ();
 b15zdnd11an1n64x5 FILLER_0_584 ();
 b15zdnd11an1n04x5 FILLER_0_648 ();
 b15zdnd00an1n01x5 FILLER_0_652 ();
 b15zdnd11an1n04x5 FILLER_0_657 ();
 b15zdnd11an1n04x5 FILLER_0_665 ();
 b15zdnd11an1n04x5 FILLER_0_711 ();
 b15zdnd00an1n02x5 FILLER_0_715 ();
 b15zdnd00an1n01x5 FILLER_0_717 ();
 b15zdnd00an1n02x5 FILLER_0_726 ();
 b15zdnd11an1n64x5 FILLER_0_770 ();
 b15zdnd11an1n32x5 FILLER_0_834 ();
 b15zdnd00an1n02x5 FILLER_0_866 ();
 b15zdnd00an1n01x5 FILLER_0_868 ();
 b15zdnd11an1n04x5 FILLER_0_880 ();
 b15zdnd11an1n04x5 FILLER_0_888 ();
 b15zdnd11an1n08x5 FILLER_0_896 ();
 b15zdnd00an1n02x5 FILLER_0_904 ();
 b15zdnd00an1n01x5 FILLER_0_906 ();
 b15zdnd11an1n32x5 FILLER_0_911 ();
 b15zdnd00an1n02x5 FILLER_0_943 ();
 b15zdnd00an1n01x5 FILLER_0_945 ();
 b15zdnd11an1n08x5 FILLER_0_950 ();
 b15zdnd11an1n04x5 FILLER_0_962 ();
 b15zdnd11an1n04x5 FILLER_0_970 ();
 b15zdnd11an1n08x5 FILLER_0_988 ();
 b15zdnd00an1n02x5 FILLER_0_996 ();
 b15zdnd00an1n01x5 FILLER_0_998 ();
 b15zdnd11an1n64x5 FILLER_0_1013 ();
 b15zdnd11an1n64x5 FILLER_0_1077 ();
 b15zdnd11an1n04x5 FILLER_0_1141 ();
 b15zdnd00an1n02x5 FILLER_0_1145 ();
 b15zdnd00an1n01x5 FILLER_0_1147 ();
 b15zdnd11an1n16x5 FILLER_0_1152 ();
 b15zdnd11an1n08x5 FILLER_0_1168 ();
 b15zdnd11an1n08x5 FILLER_0_1180 ();
 b15zdnd11an1n04x5 FILLER_0_1188 ();
 b15zdnd11an1n08x5 FILLER_0_1196 ();
 b15zdnd11an1n04x5 FILLER_0_1204 ();
 b15zdnd11an1n04x5 FILLER_0_1212 ();
 b15zdnd11an1n04x5 FILLER_0_1220 ();
 b15zdnd11an1n08x5 FILLER_0_1228 ();
 b15zdnd11an1n04x5 FILLER_0_1236 ();
 b15zdnd11an1n08x5 FILLER_0_1244 ();
 b15zdnd11an1n04x5 FILLER_0_1252 ();
 b15zdnd11an1n08x5 FILLER_0_1260 ();
 b15zdnd00an1n02x5 FILLER_0_1268 ();
 b15zdnd11an1n16x5 FILLER_0_1312 ();
 b15zdnd00an1n02x5 FILLER_0_1328 ();
 b15zdnd00an1n01x5 FILLER_0_1330 ();
 b15zdnd11an1n08x5 FILLER_0_1345 ();
 b15zdnd11an1n04x5 FILLER_0_1358 ();
 b15zdnd11an1n04x5 FILLER_0_1368 ();
 b15zdnd11an1n04x5 FILLER_0_1376 ();
 b15zdnd00an1n01x5 FILLER_0_1380 ();
 b15zdnd11an1n04x5 FILLER_0_1386 ();
 b15zdnd11an1n04x5 FILLER_0_1396 ();
 b15zdnd11an1n16x5 FILLER_0_1407 ();
 b15zdnd11an1n04x5 FILLER_0_1423 ();
 b15zdnd00an1n02x5 FILLER_0_1434 ();
 b15zdnd11an1n16x5 FILLER_0_1444 ();
 b15zdnd11an1n08x5 FILLER_0_1460 ();
 b15zdnd11an1n04x5 FILLER_0_1468 ();
 b15zdnd00an1n02x5 FILLER_0_1472 ();
 b15zdnd00an1n01x5 FILLER_0_1474 ();
 b15zdnd11an1n64x5 FILLER_0_1486 ();
 b15zdnd11an1n16x5 FILLER_0_1550 ();
 b15zdnd00an1n01x5 FILLER_0_1566 ();
 b15zdnd11an1n04x5 FILLER_0_1572 ();
 b15zdnd11an1n04x5 FILLER_0_1581 ();
 b15zdnd11an1n04x5 FILLER_0_1590 ();
 b15zdnd11an1n16x5 FILLER_0_1600 ();
 b15zdnd11an1n16x5 FILLER_0_1623 ();
 b15zdnd11an1n04x5 FILLER_0_1639 ();
 b15zdnd00an1n02x5 FILLER_0_1643 ();
 b15zdnd00an1n01x5 FILLER_0_1645 ();
 b15zdnd11an1n64x5 FILLER_0_1652 ();
 b15zdnd11an1n64x5 FILLER_0_1716 ();
 b15zdnd11an1n64x5 FILLER_0_1780 ();
 b15zdnd11an1n64x5 FILLER_0_1844 ();
 b15zdnd11an1n64x5 FILLER_0_1908 ();
 b15zdnd11an1n64x5 FILLER_0_1972 ();
 b15zdnd11an1n64x5 FILLER_0_2036 ();
 b15zdnd11an1n32x5 FILLER_0_2100 ();
 b15zdnd11an1n16x5 FILLER_0_2132 ();
 b15zdnd11an1n04x5 FILLER_0_2148 ();
 b15zdnd00an1n02x5 FILLER_0_2152 ();
 b15zdnd11an1n64x5 FILLER_0_2162 ();
 b15zdnd11an1n32x5 FILLER_0_2226 ();
 b15zdnd11an1n16x5 FILLER_0_2258 ();
 b15zdnd00an1n02x5 FILLER_0_2274 ();
 b15zdnd11an1n64x5 FILLER_1_0 ();
 b15zdnd11an1n64x5 FILLER_1_64 ();
 b15zdnd11an1n64x5 FILLER_1_128 ();
 b15zdnd11an1n64x5 FILLER_1_192 ();
 b15zdnd11an1n64x5 FILLER_1_256 ();
 b15zdnd11an1n64x5 FILLER_1_320 ();
 b15zdnd11an1n64x5 FILLER_1_384 ();
 b15zdnd11an1n64x5 FILLER_1_448 ();
 b15zdnd11an1n64x5 FILLER_1_512 ();
 b15zdnd11an1n64x5 FILLER_1_576 ();
 b15zdnd11an1n16x5 FILLER_1_640 ();
 b15zdnd00an1n02x5 FILLER_1_656 ();
 b15zdnd00an1n01x5 FILLER_1_658 ();
 b15zdnd11an1n04x5 FILLER_1_666 ();
 b15zdnd11an1n04x5 FILLER_1_677 ();
 b15zdnd11an1n04x5 FILLER_1_695 ();
 b15zdnd11an1n04x5 FILLER_1_703 ();
 b15zdnd11an1n08x5 FILLER_1_749 ();
 b15zdnd11an1n64x5 FILLER_1_765 ();
 b15zdnd11an1n64x5 FILLER_1_829 ();
 b15zdnd11an1n64x5 FILLER_1_893 ();
 b15zdnd11an1n16x5 FILLER_1_957 ();
 b15zdnd11an1n08x5 FILLER_1_973 ();
 b15zdnd00an1n01x5 FILLER_1_981 ();
 b15zdnd11an1n04x5 FILLER_1_986 ();
 b15zdnd00an1n02x5 FILLER_1_990 ();
 b15zdnd11an1n08x5 FILLER_1_1006 ();
 b15zdnd00an1n01x5 FILLER_1_1014 ();
 b15zdnd11an1n64x5 FILLER_1_1029 ();
 b15zdnd11an1n64x5 FILLER_1_1093 ();
 b15zdnd11an1n32x5 FILLER_1_1157 ();
 b15zdnd11an1n16x5 FILLER_1_1189 ();
 b15zdnd11an1n08x5 FILLER_1_1205 ();
 b15zdnd00an1n02x5 FILLER_1_1213 ();
 b15zdnd00an1n01x5 FILLER_1_1215 ();
 b15zdnd11an1n16x5 FILLER_1_1220 ();
 b15zdnd11an1n08x5 FILLER_1_1236 ();
 b15zdnd11an1n04x5 FILLER_1_1244 ();
 b15zdnd00an1n02x5 FILLER_1_1248 ();
 b15zdnd11an1n08x5 FILLER_1_1254 ();
 b15zdnd00an1n02x5 FILLER_1_1262 ();
 b15zdnd11an1n04x5 FILLER_1_1268 ();
 b15zdnd00an1n01x5 FILLER_1_1272 ();
 b15zdnd11an1n04x5 FILLER_1_1277 ();
 b15zdnd11an1n08x5 FILLER_1_1289 ();
 b15zdnd11an1n04x5 FILLER_1_1297 ();
 b15zdnd00an1n01x5 FILLER_1_1301 ();
 b15zdnd11an1n32x5 FILLER_1_1308 ();
 b15zdnd11an1n16x5 FILLER_1_1340 ();
 b15zdnd11an1n08x5 FILLER_1_1356 ();
 b15zdnd11an1n04x5 FILLER_1_1364 ();
 b15zdnd11an1n04x5 FILLER_1_1374 ();
 b15zdnd00an1n02x5 FILLER_1_1378 ();
 b15zdnd00an1n01x5 FILLER_1_1380 ();
 b15zdnd11an1n04x5 FILLER_1_1388 ();
 b15zdnd11an1n04x5 FILLER_1_1399 ();
 b15zdnd11an1n64x5 FILLER_1_1408 ();
 b15zdnd11an1n64x5 FILLER_1_1472 ();
 b15zdnd11an1n64x5 FILLER_1_1536 ();
 b15zdnd11an1n16x5 FILLER_1_1600 ();
 b15zdnd11an1n04x5 FILLER_1_1616 ();
 b15zdnd00an1n02x5 FILLER_1_1620 ();
 b15zdnd00an1n01x5 FILLER_1_1622 ();
 b15zdnd11an1n64x5 FILLER_1_1630 ();
 b15zdnd11an1n64x5 FILLER_1_1694 ();
 b15zdnd11an1n64x5 FILLER_1_1758 ();
 b15zdnd11an1n64x5 FILLER_1_1822 ();
 b15zdnd11an1n64x5 FILLER_1_1886 ();
 b15zdnd11an1n64x5 FILLER_1_1950 ();
 b15zdnd11an1n64x5 FILLER_1_2014 ();
 b15zdnd11an1n64x5 FILLER_1_2078 ();
 b15zdnd11an1n64x5 FILLER_1_2142 ();
 b15zdnd11an1n64x5 FILLER_1_2206 ();
 b15zdnd11an1n08x5 FILLER_1_2270 ();
 b15zdnd11an1n04x5 FILLER_1_2278 ();
 b15zdnd00an1n02x5 FILLER_1_2282 ();
 b15zdnd11an1n64x5 FILLER_2_8 ();
 b15zdnd11an1n64x5 FILLER_2_72 ();
 b15zdnd11an1n64x5 FILLER_2_136 ();
 b15zdnd11an1n64x5 FILLER_2_200 ();
 b15zdnd11an1n64x5 FILLER_2_264 ();
 b15zdnd11an1n64x5 FILLER_2_328 ();
 b15zdnd11an1n64x5 FILLER_2_392 ();
 b15zdnd11an1n64x5 FILLER_2_456 ();
 b15zdnd11an1n64x5 FILLER_2_520 ();
 b15zdnd11an1n64x5 FILLER_2_584 ();
 b15zdnd11an1n16x5 FILLER_2_648 ();
 b15zdnd00an1n02x5 FILLER_2_664 ();
 b15zdnd00an1n01x5 FILLER_2_666 ();
 b15zdnd11an1n08x5 FILLER_2_709 ();
 b15zdnd00an1n01x5 FILLER_2_717 ();
 b15zdnd00an1n02x5 FILLER_2_726 ();
 b15zdnd11an1n16x5 FILLER_2_732 ();
 b15zdnd11an1n08x5 FILLER_2_748 ();
 b15zdnd00an1n02x5 FILLER_2_756 ();
 b15zdnd11an1n64x5 FILLER_2_772 ();
 b15zdnd11an1n64x5 FILLER_2_836 ();
 b15zdnd11an1n64x5 FILLER_2_900 ();
 b15zdnd00an1n01x5 FILLER_2_964 ();
 b15zdnd11an1n32x5 FILLER_2_979 ();
 b15zdnd11an1n04x5 FILLER_2_1011 ();
 b15zdnd00an1n01x5 FILLER_2_1015 ();
 b15zdnd11an1n64x5 FILLER_2_1030 ();
 b15zdnd11an1n64x5 FILLER_2_1094 ();
 b15zdnd11an1n32x5 FILLER_2_1158 ();
 b15zdnd11an1n08x5 FILLER_2_1190 ();
 b15zdnd11an1n04x5 FILLER_2_1198 ();
 b15zdnd00an1n01x5 FILLER_2_1202 ();
 b15zdnd11an1n64x5 FILLER_2_1207 ();
 b15zdnd11an1n32x5 FILLER_2_1271 ();
 b15zdnd11an1n16x5 FILLER_2_1303 ();
 b15zdnd11an1n08x5 FILLER_2_1319 ();
 b15zdnd00an1n02x5 FILLER_2_1327 ();
 b15zdnd11an1n64x5 FILLER_2_1340 ();
 b15zdnd11an1n64x5 FILLER_2_1404 ();
 b15zdnd11an1n64x5 FILLER_2_1468 ();
 b15zdnd11an1n64x5 FILLER_2_1532 ();
 b15zdnd11an1n64x5 FILLER_2_1596 ();
 b15zdnd11an1n64x5 FILLER_2_1660 ();
 b15zdnd11an1n64x5 FILLER_2_1724 ();
 b15zdnd11an1n64x5 FILLER_2_1788 ();
 b15zdnd11an1n64x5 FILLER_2_1852 ();
 b15zdnd11an1n64x5 FILLER_2_1916 ();
 b15zdnd11an1n64x5 FILLER_2_1980 ();
 b15zdnd11an1n64x5 FILLER_2_2044 ();
 b15zdnd11an1n32x5 FILLER_2_2108 ();
 b15zdnd11an1n08x5 FILLER_2_2140 ();
 b15zdnd11an1n04x5 FILLER_2_2148 ();
 b15zdnd00an1n02x5 FILLER_2_2152 ();
 b15zdnd11an1n64x5 FILLER_2_2162 ();
 b15zdnd11an1n32x5 FILLER_2_2226 ();
 b15zdnd11an1n16x5 FILLER_2_2258 ();
 b15zdnd00an1n02x5 FILLER_2_2274 ();
 b15zdnd11an1n64x5 FILLER_3_0 ();
 b15zdnd11an1n64x5 FILLER_3_64 ();
 b15zdnd11an1n64x5 FILLER_3_128 ();
 b15zdnd11an1n64x5 FILLER_3_192 ();
 b15zdnd11an1n64x5 FILLER_3_256 ();
 b15zdnd11an1n64x5 FILLER_3_320 ();
 b15zdnd11an1n64x5 FILLER_3_384 ();
 b15zdnd11an1n64x5 FILLER_3_448 ();
 b15zdnd11an1n64x5 FILLER_3_512 ();
 b15zdnd11an1n64x5 FILLER_3_576 ();
 b15zdnd11an1n32x5 FILLER_3_640 ();
 b15zdnd11an1n08x5 FILLER_3_672 ();
 b15zdnd00an1n01x5 FILLER_3_680 ();
 b15zdnd11an1n08x5 FILLER_3_689 ();
 b15zdnd11an1n04x5 FILLER_3_697 ();
 b15zdnd00an1n01x5 FILLER_3_701 ();
 b15zdnd11an1n64x5 FILLER_3_744 ();
 b15zdnd11an1n64x5 FILLER_3_808 ();
 b15zdnd11an1n64x5 FILLER_3_872 ();
 b15zdnd11an1n32x5 FILLER_3_936 ();
 b15zdnd11an1n04x5 FILLER_3_968 ();
 b15zdnd00an1n01x5 FILLER_3_972 ();
 b15zdnd11an1n08x5 FILLER_3_985 ();
 b15zdnd11an1n04x5 FILLER_3_993 ();
 b15zdnd00an1n02x5 FILLER_3_997 ();
 b15zdnd00an1n01x5 FILLER_3_999 ();
 b15zdnd11an1n64x5 FILLER_3_1004 ();
 b15zdnd11an1n64x5 FILLER_3_1068 ();
 b15zdnd11an1n64x5 FILLER_3_1132 ();
 b15zdnd11an1n64x5 FILLER_3_1196 ();
 b15zdnd11an1n64x5 FILLER_3_1260 ();
 b15zdnd11an1n64x5 FILLER_3_1324 ();
 b15zdnd11an1n04x5 FILLER_3_1388 ();
 b15zdnd00an1n02x5 FILLER_3_1392 ();
 b15zdnd11an1n64x5 FILLER_3_1400 ();
 b15zdnd11an1n64x5 FILLER_3_1464 ();
 b15zdnd11an1n64x5 FILLER_3_1528 ();
 b15zdnd11an1n64x5 FILLER_3_1592 ();
 b15zdnd11an1n64x5 FILLER_3_1656 ();
 b15zdnd11an1n64x5 FILLER_3_1720 ();
 b15zdnd11an1n64x5 FILLER_3_1784 ();
 b15zdnd11an1n64x5 FILLER_3_1848 ();
 b15zdnd11an1n64x5 FILLER_3_1912 ();
 b15zdnd11an1n64x5 FILLER_3_1976 ();
 b15zdnd11an1n64x5 FILLER_3_2040 ();
 b15zdnd11an1n64x5 FILLER_3_2104 ();
 b15zdnd11an1n64x5 FILLER_3_2168 ();
 b15zdnd11an1n32x5 FILLER_3_2232 ();
 b15zdnd11an1n16x5 FILLER_3_2264 ();
 b15zdnd11an1n04x5 FILLER_3_2280 ();
 b15zdnd11an1n64x5 FILLER_4_8 ();
 b15zdnd11an1n64x5 FILLER_4_72 ();
 b15zdnd11an1n64x5 FILLER_4_136 ();
 b15zdnd11an1n64x5 FILLER_4_200 ();
 b15zdnd11an1n64x5 FILLER_4_264 ();
 b15zdnd11an1n64x5 FILLER_4_328 ();
 b15zdnd11an1n64x5 FILLER_4_392 ();
 b15zdnd11an1n64x5 FILLER_4_456 ();
 b15zdnd11an1n64x5 FILLER_4_520 ();
 b15zdnd11an1n64x5 FILLER_4_584 ();
 b15zdnd11an1n32x5 FILLER_4_648 ();
 b15zdnd11an1n08x5 FILLER_4_687 ();
 b15zdnd11an1n04x5 FILLER_4_695 ();
 b15zdnd11an1n04x5 FILLER_4_706 ();
 b15zdnd11an1n04x5 FILLER_4_714 ();
 b15zdnd11an1n64x5 FILLER_4_726 ();
 b15zdnd11an1n64x5 FILLER_4_790 ();
 b15zdnd11an1n64x5 FILLER_4_854 ();
 b15zdnd11an1n32x5 FILLER_4_918 ();
 b15zdnd11an1n04x5 FILLER_4_950 ();
 b15zdnd11an1n64x5 FILLER_4_965 ();
 b15zdnd11an1n64x5 FILLER_4_1029 ();
 b15zdnd11an1n64x5 FILLER_4_1093 ();
 b15zdnd11an1n64x5 FILLER_4_1157 ();
 b15zdnd11an1n64x5 FILLER_4_1221 ();
 b15zdnd11an1n64x5 FILLER_4_1285 ();
 b15zdnd11an1n64x5 FILLER_4_1349 ();
 b15zdnd11an1n64x5 FILLER_4_1413 ();
 b15zdnd00an1n01x5 FILLER_4_1477 ();
 b15zdnd11an1n08x5 FILLER_4_2265 ();
 b15zdnd00an1n02x5 FILLER_4_2273 ();
 b15zdnd00an1n01x5 FILLER_4_2275 ();
 b15zdnd11an1n64x5 FILLER_5_0 ();
 b15zdnd11an1n64x5 FILLER_5_64 ();
 b15zdnd11an1n64x5 FILLER_5_128 ();
 b15zdnd11an1n64x5 FILLER_5_192 ();
 b15zdnd11an1n64x5 FILLER_5_256 ();
 b15zdnd11an1n64x5 FILLER_5_320 ();
 b15zdnd11an1n64x5 FILLER_5_384 ();
 b15zdnd11an1n64x5 FILLER_5_448 ();
 b15zdnd11an1n64x5 FILLER_5_512 ();
 b15zdnd11an1n64x5 FILLER_5_576 ();
 b15zdnd11an1n64x5 FILLER_5_640 ();
 b15zdnd11an1n64x5 FILLER_5_704 ();
 b15zdnd11an1n64x5 FILLER_5_768 ();
 b15zdnd11an1n64x5 FILLER_5_832 ();
 b15zdnd11an1n64x5 FILLER_5_896 ();
 b15zdnd11an1n64x5 FILLER_5_960 ();
 b15zdnd11an1n64x5 FILLER_5_1024 ();
 b15zdnd11an1n64x5 FILLER_5_1088 ();
 b15zdnd11an1n64x5 FILLER_5_1152 ();
 b15zdnd11an1n64x5 FILLER_5_1216 ();
 b15zdnd11an1n64x5 FILLER_5_1280 ();
 b15zdnd11an1n64x5 FILLER_5_1344 ();
 b15zdnd11an1n64x5 FILLER_5_1408 ();
 b15zdnd11an1n08x5 FILLER_5_1472 ();
 b15zdnd11an1n04x5 FILLER_5_1480 ();
 b15zdnd00an1n02x5 FILLER_5_1484 ();
 b15zdnd11an1n16x5 FILLER_5_2257 ();
 b15zdnd11an1n08x5 FILLER_5_2273 ();
 b15zdnd00an1n02x5 FILLER_5_2281 ();
 b15zdnd00an1n01x5 FILLER_5_2283 ();
 b15zdnd11an1n64x5 FILLER_6_8 ();
 b15zdnd11an1n64x5 FILLER_6_72 ();
 b15zdnd11an1n64x5 FILLER_6_136 ();
 b15zdnd11an1n64x5 FILLER_6_200 ();
 b15zdnd11an1n64x5 FILLER_6_264 ();
 b15zdnd11an1n64x5 FILLER_6_328 ();
 b15zdnd11an1n64x5 FILLER_6_392 ();
 b15zdnd11an1n64x5 FILLER_6_456 ();
 b15zdnd11an1n64x5 FILLER_6_520 ();
 b15zdnd11an1n64x5 FILLER_6_584 ();
 b15zdnd11an1n64x5 FILLER_6_648 ();
 b15zdnd11an1n04x5 FILLER_6_712 ();
 b15zdnd00an1n02x5 FILLER_6_716 ();
 b15zdnd11an1n64x5 FILLER_6_726 ();
 b15zdnd11an1n64x5 FILLER_6_790 ();
 b15zdnd11an1n64x5 FILLER_6_854 ();
 b15zdnd11an1n64x5 FILLER_6_918 ();
 b15zdnd11an1n64x5 FILLER_6_982 ();
 b15zdnd11an1n64x5 FILLER_6_1046 ();
 b15zdnd11an1n64x5 FILLER_6_1110 ();
 b15zdnd11an1n64x5 FILLER_6_1174 ();
 b15zdnd11an1n64x5 FILLER_6_1238 ();
 b15zdnd11an1n64x5 FILLER_6_1302 ();
 b15zdnd11an1n64x5 FILLER_6_1366 ();
 b15zdnd11an1n32x5 FILLER_6_1430 ();
 b15zdnd11an1n16x5 FILLER_6_1462 ();
 b15zdnd11an1n08x5 FILLER_6_2265 ();
 b15zdnd00an1n02x5 FILLER_6_2273 ();
 b15zdnd00an1n01x5 FILLER_6_2275 ();
 b15zdnd11an1n64x5 FILLER_7_0 ();
 b15zdnd11an1n64x5 FILLER_7_64 ();
 b15zdnd11an1n64x5 FILLER_7_128 ();
 b15zdnd11an1n64x5 FILLER_7_192 ();
 b15zdnd11an1n64x5 FILLER_7_256 ();
 b15zdnd11an1n64x5 FILLER_7_320 ();
 b15zdnd11an1n64x5 FILLER_7_384 ();
 b15zdnd11an1n64x5 FILLER_7_448 ();
 b15zdnd11an1n64x5 FILLER_7_512 ();
 b15zdnd11an1n64x5 FILLER_7_576 ();
 b15zdnd11an1n64x5 FILLER_7_640 ();
 b15zdnd11an1n64x5 FILLER_7_704 ();
 b15zdnd11an1n64x5 FILLER_7_768 ();
 b15zdnd11an1n64x5 FILLER_7_832 ();
 b15zdnd11an1n64x5 FILLER_7_896 ();
 b15zdnd11an1n64x5 FILLER_7_960 ();
 b15zdnd11an1n64x5 FILLER_7_1024 ();
 b15zdnd11an1n64x5 FILLER_7_1088 ();
 b15zdnd11an1n64x5 FILLER_7_1152 ();
 b15zdnd11an1n64x5 FILLER_7_1216 ();
 b15zdnd11an1n64x5 FILLER_7_1280 ();
 b15zdnd11an1n64x5 FILLER_7_1344 ();
 b15zdnd11an1n64x5 FILLER_7_1408 ();
 b15zdnd11an1n08x5 FILLER_7_1472 ();
 b15zdnd11an1n04x5 FILLER_7_1480 ();
 b15zdnd00an1n02x5 FILLER_7_1484 ();
 b15zdnd11an1n16x5 FILLER_7_2257 ();
 b15zdnd11an1n08x5 FILLER_7_2273 ();
 b15zdnd00an1n02x5 FILLER_7_2281 ();
 b15zdnd00an1n01x5 FILLER_7_2283 ();
 b15zdnd11an1n64x5 FILLER_8_8 ();
 b15zdnd11an1n64x5 FILLER_8_72 ();
 b15zdnd11an1n64x5 FILLER_8_136 ();
 b15zdnd11an1n64x5 FILLER_8_200 ();
 b15zdnd11an1n64x5 FILLER_8_264 ();
 b15zdnd11an1n64x5 FILLER_8_328 ();
 b15zdnd11an1n64x5 FILLER_8_392 ();
 b15zdnd11an1n64x5 FILLER_8_456 ();
 b15zdnd11an1n64x5 FILLER_8_520 ();
 b15zdnd11an1n64x5 FILLER_8_584 ();
 b15zdnd11an1n64x5 FILLER_8_648 ();
 b15zdnd11an1n04x5 FILLER_8_712 ();
 b15zdnd00an1n02x5 FILLER_8_716 ();
 b15zdnd11an1n64x5 FILLER_8_726 ();
 b15zdnd11an1n64x5 FILLER_8_790 ();
 b15zdnd11an1n64x5 FILLER_8_854 ();
 b15zdnd11an1n04x5 FILLER_8_918 ();
 b15zdnd11an1n64x5 FILLER_8_964 ();
 b15zdnd11an1n16x5 FILLER_8_1028 ();
 b15zdnd00an1n01x5 FILLER_8_1044 ();
 b15zdnd11an1n64x5 FILLER_8_1087 ();
 b15zdnd11an1n64x5 FILLER_8_1151 ();
 b15zdnd11an1n64x5 FILLER_8_1215 ();
 b15zdnd11an1n64x5 FILLER_8_1279 ();
 b15zdnd11an1n64x5 FILLER_8_1343 ();
 b15zdnd11an1n64x5 FILLER_8_1407 ();
 b15zdnd11an1n04x5 FILLER_8_1471 ();
 b15zdnd00an1n02x5 FILLER_8_1475 ();
 b15zdnd00an1n01x5 FILLER_8_1477 ();
 b15zdnd11an1n08x5 FILLER_8_2265 ();
 b15zdnd00an1n02x5 FILLER_8_2273 ();
 b15zdnd00an1n01x5 FILLER_8_2275 ();
 b15zdnd11an1n64x5 FILLER_9_0 ();
 b15zdnd11an1n64x5 FILLER_9_64 ();
 b15zdnd11an1n64x5 FILLER_9_128 ();
 b15zdnd11an1n64x5 FILLER_9_192 ();
 b15zdnd11an1n64x5 FILLER_9_256 ();
 b15zdnd11an1n64x5 FILLER_9_320 ();
 b15zdnd11an1n64x5 FILLER_9_384 ();
 b15zdnd11an1n64x5 FILLER_9_448 ();
 b15zdnd11an1n64x5 FILLER_9_512 ();
 b15zdnd11an1n64x5 FILLER_9_576 ();
 b15zdnd11an1n64x5 FILLER_9_640 ();
 b15zdnd11an1n32x5 FILLER_9_704 ();
 b15zdnd11an1n16x5 FILLER_9_736 ();
 b15zdnd11an1n04x5 FILLER_9_752 ();
 b15zdnd00an1n02x5 FILLER_9_756 ();
 b15zdnd11an1n32x5 FILLER_9_800 ();
 b15zdnd11an1n08x5 FILLER_9_832 ();
 b15zdnd00an1n02x5 FILLER_9_840 ();
 b15zdnd00an1n01x5 FILLER_9_842 ();
 b15zdnd11an1n08x5 FILLER_9_885 ();
 b15zdnd00an1n02x5 FILLER_9_893 ();
 b15zdnd00an1n01x5 FILLER_9_895 ();
 b15zdnd11an1n04x5 FILLER_9_938 ();
 b15zdnd11an1n32x5 FILLER_9_984 ();
 b15zdnd11an1n16x5 FILLER_9_1016 ();
 b15zdnd11an1n08x5 FILLER_9_1032 ();
 b15zdnd11an1n04x5 FILLER_9_1040 ();
 b15zdnd00an1n02x5 FILLER_9_1044 ();
 b15zdnd11an1n64x5 FILLER_9_1088 ();
 b15zdnd11an1n32x5 FILLER_9_1152 ();
 b15zdnd11an1n16x5 FILLER_9_1184 ();
 b15zdnd11an1n08x5 FILLER_9_1200 ();
 b15zdnd00an1n02x5 FILLER_9_1208 ();
 b15zdnd00an1n01x5 FILLER_9_1210 ();
 b15zdnd11an1n16x5 FILLER_9_1253 ();
 b15zdnd11an1n08x5 FILLER_9_1269 ();
 b15zdnd11an1n04x5 FILLER_9_1277 ();
 b15zdnd11an1n64x5 FILLER_9_1323 ();
 b15zdnd11an1n64x5 FILLER_9_1387 ();
 b15zdnd11an1n32x5 FILLER_9_1451 ();
 b15zdnd00an1n02x5 FILLER_9_1483 ();
 b15zdnd00an1n01x5 FILLER_9_1485 ();
 b15zdnd11an1n16x5 FILLER_9_2257 ();
 b15zdnd11an1n08x5 FILLER_9_2273 ();
 b15zdnd00an1n02x5 FILLER_9_2281 ();
 b15zdnd00an1n01x5 FILLER_9_2283 ();
 b15zdnd11an1n64x5 FILLER_10_8 ();
 b15zdnd11an1n64x5 FILLER_10_72 ();
 b15zdnd11an1n64x5 FILLER_10_136 ();
 b15zdnd11an1n64x5 FILLER_10_200 ();
 b15zdnd11an1n64x5 FILLER_10_264 ();
 b15zdnd11an1n64x5 FILLER_10_328 ();
 b15zdnd11an1n64x5 FILLER_10_392 ();
 b15zdnd11an1n64x5 FILLER_10_456 ();
 b15zdnd11an1n64x5 FILLER_10_520 ();
 b15zdnd11an1n64x5 FILLER_10_584 ();
 b15zdnd11an1n64x5 FILLER_10_648 ();
 b15zdnd11an1n04x5 FILLER_10_712 ();
 b15zdnd00an1n02x5 FILLER_10_716 ();
 b15zdnd11an1n64x5 FILLER_10_726 ();
 b15zdnd11an1n64x5 FILLER_10_790 ();
 b15zdnd11an1n04x5 FILLER_10_854 ();
 b15zdnd00an1n01x5 FILLER_10_858 ();
 b15zdnd11an1n32x5 FILLER_10_901 ();
 b15zdnd11an1n08x5 FILLER_10_933 ();
 b15zdnd11an1n04x5 FILLER_10_941 ();
 b15zdnd00an1n02x5 FILLER_10_945 ();
 b15zdnd00an1n01x5 FILLER_10_947 ();
 b15zdnd11an1n32x5 FILLER_10_990 ();
 b15zdnd11an1n64x5 FILLER_10_1064 ();
 b15zdnd11an1n32x5 FILLER_10_1128 ();
 b15zdnd11an1n16x5 FILLER_10_1160 ();
 b15zdnd11an1n08x5 FILLER_10_1176 ();
 b15zdnd11an1n32x5 FILLER_10_1226 ();
 b15zdnd11an1n16x5 FILLER_10_1258 ();
 b15zdnd00an1n01x5 FILLER_10_1274 ();
 b15zdnd11an1n64x5 FILLER_10_1317 ();
 b15zdnd11an1n64x5 FILLER_10_1381 ();
 b15zdnd11an1n32x5 FILLER_10_1445 ();
 b15zdnd00an1n01x5 FILLER_10_1477 ();
 b15zdnd11an1n08x5 FILLER_10_2265 ();
 b15zdnd00an1n02x5 FILLER_10_2273 ();
 b15zdnd00an1n01x5 FILLER_10_2275 ();
 b15zdnd11an1n64x5 FILLER_11_0 ();
 b15zdnd11an1n64x5 FILLER_11_64 ();
 b15zdnd11an1n64x5 FILLER_11_128 ();
 b15zdnd11an1n64x5 FILLER_11_192 ();
 b15zdnd11an1n64x5 FILLER_11_256 ();
 b15zdnd11an1n64x5 FILLER_11_320 ();
 b15zdnd11an1n64x5 FILLER_11_384 ();
 b15zdnd11an1n64x5 FILLER_11_448 ();
 b15zdnd11an1n64x5 FILLER_11_512 ();
 b15zdnd11an1n64x5 FILLER_11_576 ();
 b15zdnd11an1n64x5 FILLER_11_640 ();
 b15zdnd11an1n64x5 FILLER_11_704 ();
 b15zdnd11an1n64x5 FILLER_11_768 ();
 b15zdnd11an1n16x5 FILLER_11_832 ();
 b15zdnd11an1n08x5 FILLER_11_848 ();
 b15zdnd11an1n04x5 FILLER_11_856 ();
 b15zdnd00an1n02x5 FILLER_11_860 ();
 b15zdnd00an1n01x5 FILLER_11_862 ();
 b15zdnd11an1n16x5 FILLER_11_905 ();
 b15zdnd11an1n08x5 FILLER_11_921 ();
 b15zdnd11an1n04x5 FILLER_11_929 ();
 b15zdnd11an1n16x5 FILLER_11_975 ();
 b15zdnd00an1n02x5 FILLER_11_991 ();
 b15zdnd11an1n64x5 FILLER_11_1035 ();
 b15zdnd11an1n64x5 FILLER_11_1099 ();
 b15zdnd11an1n64x5 FILLER_11_1163 ();
 b15zdnd11an1n04x5 FILLER_11_1227 ();
 b15zdnd00an1n01x5 FILLER_11_1231 ();
 b15zdnd11an1n64x5 FILLER_11_1274 ();
 b15zdnd11an1n64x5 FILLER_11_1338 ();
 b15zdnd11an1n64x5 FILLER_11_1402 ();
 b15zdnd11an1n16x5 FILLER_11_1466 ();
 b15zdnd11an1n04x5 FILLER_11_1482 ();
 b15zdnd11an1n16x5 FILLER_11_2257 ();
 b15zdnd11an1n08x5 FILLER_11_2273 ();
 b15zdnd00an1n02x5 FILLER_11_2281 ();
 b15zdnd00an1n01x5 FILLER_11_2283 ();
 b15zdnd11an1n64x5 FILLER_12_8 ();
 b15zdnd11an1n64x5 FILLER_12_72 ();
 b15zdnd11an1n64x5 FILLER_12_136 ();
 b15zdnd11an1n64x5 FILLER_12_200 ();
 b15zdnd11an1n64x5 FILLER_12_264 ();
 b15zdnd11an1n64x5 FILLER_12_328 ();
 b15zdnd11an1n64x5 FILLER_12_392 ();
 b15zdnd11an1n64x5 FILLER_12_456 ();
 b15zdnd11an1n64x5 FILLER_12_520 ();
 b15zdnd11an1n64x5 FILLER_12_584 ();
 b15zdnd11an1n64x5 FILLER_12_648 ();
 b15zdnd11an1n04x5 FILLER_12_712 ();
 b15zdnd00an1n02x5 FILLER_12_716 ();
 b15zdnd11an1n64x5 FILLER_12_726 ();
 b15zdnd11an1n64x5 FILLER_12_790 ();
 b15zdnd00an1n01x5 FILLER_12_854 ();
 b15zdnd11an1n64x5 FILLER_12_897 ();
 b15zdnd11an1n64x5 FILLER_12_961 ();
 b15zdnd11an1n64x5 FILLER_12_1067 ();
 b15zdnd11an1n64x5 FILLER_12_1131 ();
 b15zdnd11an1n04x5 FILLER_12_1195 ();
 b15zdnd00an1n01x5 FILLER_12_1199 ();
 b15zdnd11an1n04x5 FILLER_12_1242 ();
 b15zdnd11an1n64x5 FILLER_12_1288 ();
 b15zdnd11an1n64x5 FILLER_12_1352 ();
 b15zdnd11an1n32x5 FILLER_12_1416 ();
 b15zdnd11an1n16x5 FILLER_12_1448 ();
 b15zdnd11an1n08x5 FILLER_12_1464 ();
 b15zdnd11an1n04x5 FILLER_12_1472 ();
 b15zdnd00an1n02x5 FILLER_12_1476 ();
 b15zdnd11an1n08x5 FILLER_12_2265 ();
 b15zdnd00an1n02x5 FILLER_12_2273 ();
 b15zdnd00an1n01x5 FILLER_12_2275 ();
 b15zdnd11an1n64x5 FILLER_13_0 ();
 b15zdnd11an1n64x5 FILLER_13_64 ();
 b15zdnd11an1n64x5 FILLER_13_128 ();
 b15zdnd11an1n64x5 FILLER_13_192 ();
 b15zdnd11an1n64x5 FILLER_13_256 ();
 b15zdnd11an1n64x5 FILLER_13_320 ();
 b15zdnd11an1n64x5 FILLER_13_384 ();
 b15zdnd11an1n64x5 FILLER_13_448 ();
 b15zdnd11an1n64x5 FILLER_13_512 ();
 b15zdnd11an1n64x5 FILLER_13_576 ();
 b15zdnd11an1n64x5 FILLER_13_640 ();
 b15zdnd11an1n64x5 FILLER_13_704 ();
 b15zdnd11an1n64x5 FILLER_13_768 ();
 b15zdnd11an1n08x5 FILLER_13_832 ();
 b15zdnd11an1n04x5 FILLER_13_840 ();
 b15zdnd11an1n64x5 FILLER_13_886 ();
 b15zdnd11an1n64x5 FILLER_13_950 ();
 b15zdnd11an1n64x5 FILLER_13_1014 ();
 b15zdnd11an1n64x5 FILLER_13_1078 ();
 b15zdnd11an1n08x5 FILLER_13_1142 ();
 b15zdnd11an1n64x5 FILLER_13_1192 ();
 b15zdnd11an1n64x5 FILLER_13_1256 ();
 b15zdnd11an1n64x5 FILLER_13_1320 ();
 b15zdnd11an1n64x5 FILLER_13_1384 ();
 b15zdnd11an1n32x5 FILLER_13_1448 ();
 b15zdnd11an1n04x5 FILLER_13_1480 ();
 b15zdnd00an1n02x5 FILLER_13_1484 ();
 b15zdnd11an1n16x5 FILLER_13_2257 ();
 b15zdnd11an1n08x5 FILLER_13_2273 ();
 b15zdnd00an1n02x5 FILLER_13_2281 ();
 b15zdnd00an1n01x5 FILLER_13_2283 ();
 b15zdnd11an1n64x5 FILLER_14_8 ();
 b15zdnd11an1n64x5 FILLER_14_72 ();
 b15zdnd11an1n64x5 FILLER_14_136 ();
 b15zdnd11an1n64x5 FILLER_14_200 ();
 b15zdnd11an1n64x5 FILLER_14_264 ();
 b15zdnd11an1n64x5 FILLER_14_328 ();
 b15zdnd11an1n64x5 FILLER_14_392 ();
 b15zdnd11an1n64x5 FILLER_14_456 ();
 b15zdnd11an1n64x5 FILLER_14_520 ();
 b15zdnd11an1n64x5 FILLER_14_584 ();
 b15zdnd11an1n32x5 FILLER_14_648 ();
 b15zdnd11an1n04x5 FILLER_14_680 ();
 b15zdnd11an1n04x5 FILLER_14_687 ();
 b15zdnd11an1n16x5 FILLER_14_694 ();
 b15zdnd11an1n08x5 FILLER_14_710 ();
 b15zdnd11an1n64x5 FILLER_14_726 ();
 b15zdnd11an1n64x5 FILLER_14_790 ();
 b15zdnd11an1n64x5 FILLER_14_854 ();
 b15zdnd11an1n64x5 FILLER_14_918 ();
 b15zdnd11an1n64x5 FILLER_14_982 ();
 b15zdnd11an1n64x5 FILLER_14_1046 ();
 b15zdnd11an1n64x5 FILLER_14_1110 ();
 b15zdnd11an1n64x5 FILLER_14_1174 ();
 b15zdnd11an1n64x5 FILLER_14_1238 ();
 b15zdnd11an1n64x5 FILLER_14_1302 ();
 b15zdnd11an1n64x5 FILLER_14_1366 ();
 b15zdnd11an1n32x5 FILLER_14_1430 ();
 b15zdnd11an1n16x5 FILLER_14_1462 ();
 b15zdnd11an1n08x5 FILLER_14_2265 ();
 b15zdnd00an1n02x5 FILLER_14_2273 ();
 b15zdnd00an1n01x5 FILLER_14_2275 ();
 b15zdnd11an1n64x5 FILLER_15_0 ();
 b15zdnd11an1n64x5 FILLER_15_64 ();
 b15zdnd11an1n64x5 FILLER_15_128 ();
 b15zdnd11an1n64x5 FILLER_15_192 ();
 b15zdnd11an1n64x5 FILLER_15_256 ();
 b15zdnd11an1n64x5 FILLER_15_320 ();
 b15zdnd11an1n64x5 FILLER_15_384 ();
 b15zdnd11an1n64x5 FILLER_15_448 ();
 b15zdnd11an1n64x5 FILLER_15_512 ();
 b15zdnd11an1n64x5 FILLER_15_576 ();
 b15zdnd11an1n32x5 FILLER_15_640 ();
 b15zdnd11an1n08x5 FILLER_15_672 ();
 b15zdnd00an1n02x5 FILLER_15_680 ();
 b15zdnd00an1n01x5 FILLER_15_682 ();
 b15zdnd11an1n16x5 FILLER_15_686 ();
 b15zdnd11an1n08x5 FILLER_15_702 ();
 b15zdnd00an1n01x5 FILLER_15_710 ();
 b15zdnd11an1n04x5 FILLER_15_714 ();
 b15zdnd00an1n02x5 FILLER_15_718 ();
 b15zdnd11an1n64x5 FILLER_15_723 ();
 b15zdnd11an1n64x5 FILLER_15_787 ();
 b15zdnd11an1n64x5 FILLER_15_851 ();
 b15zdnd11an1n64x5 FILLER_15_915 ();
 b15zdnd11an1n64x5 FILLER_15_979 ();
 b15zdnd11an1n64x5 FILLER_15_1043 ();
 b15zdnd11an1n64x5 FILLER_15_1107 ();
 b15zdnd11an1n64x5 FILLER_15_1171 ();
 b15zdnd11an1n64x5 FILLER_15_1235 ();
 b15zdnd11an1n64x5 FILLER_15_1299 ();
 b15zdnd11an1n64x5 FILLER_15_1363 ();
 b15zdnd11an1n32x5 FILLER_15_1427 ();
 b15zdnd11an1n16x5 FILLER_15_1459 ();
 b15zdnd11an1n08x5 FILLER_15_1475 ();
 b15zdnd00an1n02x5 FILLER_15_1483 ();
 b15zdnd00an1n01x5 FILLER_15_1485 ();
 b15zdnd11an1n16x5 FILLER_15_2257 ();
 b15zdnd11an1n08x5 FILLER_15_2273 ();
 b15zdnd00an1n02x5 FILLER_15_2281 ();
 b15zdnd00an1n01x5 FILLER_15_2283 ();
 b15zdnd11an1n64x5 FILLER_16_8 ();
 b15zdnd11an1n64x5 FILLER_16_72 ();
 b15zdnd11an1n64x5 FILLER_16_136 ();
 b15zdnd11an1n64x5 FILLER_16_200 ();
 b15zdnd11an1n64x5 FILLER_16_264 ();
 b15zdnd11an1n64x5 FILLER_16_328 ();
 b15zdnd11an1n32x5 FILLER_16_392 ();
 b15zdnd11an1n04x5 FILLER_16_424 ();
 b15zdnd00an1n02x5 FILLER_16_428 ();
 b15zdnd00an1n01x5 FILLER_16_430 ();
 b15zdnd11an1n64x5 FILLER_16_476 ();
 b15zdnd11an1n64x5 FILLER_16_540 ();
 b15zdnd11an1n32x5 FILLER_16_604 ();
 b15zdnd11an1n16x5 FILLER_16_636 ();
 b15zdnd11an1n08x5 FILLER_16_652 ();
 b15zdnd11an1n04x5 FILLER_16_663 ();
 b15zdnd11an1n04x5 FILLER_16_670 ();
 b15zdnd11an1n04x5 FILLER_16_677 ();
 b15zdnd00an1n02x5 FILLER_16_681 ();
 b15zdnd11an1n04x5 FILLER_16_686 ();
 b15zdnd11an1n08x5 FILLER_16_693 ();
 b15zdnd00an1n02x5 FILLER_16_701 ();
 b15zdnd00an1n01x5 FILLER_16_703 ();
 b15zdnd11an1n04x5 FILLER_16_707 ();
 b15zdnd00an1n02x5 FILLER_16_711 ();
 b15zdnd00an1n02x5 FILLER_16_716 ();
 b15zdnd11an1n64x5 FILLER_16_726 ();
 b15zdnd11an1n64x5 FILLER_16_790 ();
 b15zdnd11an1n04x5 FILLER_16_854 ();
 b15zdnd00an1n02x5 FILLER_16_858 ();
 b15zdnd00an1n01x5 FILLER_16_860 ();
 b15zdnd11an1n08x5 FILLER_16_869 ();
 b15zdnd00an1n01x5 FILLER_16_877 ();
 b15zdnd11an1n32x5 FILLER_16_891 ();
 b15zdnd00an1n02x5 FILLER_16_923 ();
 b15zdnd00an1n01x5 FILLER_16_925 ();
 b15zdnd11an1n16x5 FILLER_16_939 ();
 b15zdnd11an1n64x5 FILLER_16_961 ();
 b15zdnd11an1n08x5 FILLER_16_1025 ();
 b15zdnd11an1n04x5 FILLER_16_1033 ();
 b15zdnd00an1n02x5 FILLER_16_1037 ();
 b15zdnd00an1n01x5 FILLER_16_1039 ();
 b15zdnd11an1n64x5 FILLER_16_1050 ();
 b15zdnd11an1n64x5 FILLER_16_1114 ();
 b15zdnd11an1n64x5 FILLER_16_1178 ();
 b15zdnd11an1n64x5 FILLER_16_1242 ();
 b15zdnd11an1n64x5 FILLER_16_1306 ();
 b15zdnd11an1n64x5 FILLER_16_1370 ();
 b15zdnd11an1n32x5 FILLER_16_1434 ();
 b15zdnd11an1n08x5 FILLER_16_1466 ();
 b15zdnd11an1n04x5 FILLER_16_1474 ();
 b15zdnd11an1n08x5 FILLER_16_2265 ();
 b15zdnd00an1n02x5 FILLER_16_2273 ();
 b15zdnd00an1n01x5 FILLER_16_2275 ();
 b15zdnd11an1n64x5 FILLER_17_0 ();
 b15zdnd11an1n64x5 FILLER_17_64 ();
 b15zdnd11an1n64x5 FILLER_17_128 ();
 b15zdnd11an1n64x5 FILLER_17_192 ();
 b15zdnd11an1n64x5 FILLER_17_256 ();
 b15zdnd11an1n64x5 FILLER_17_320 ();
 b15zdnd11an1n64x5 FILLER_17_384 ();
 b15zdnd11an1n64x5 FILLER_17_448 ();
 b15zdnd11an1n64x5 FILLER_17_512 ();
 b15zdnd11an1n16x5 FILLER_17_588 ();
 b15zdnd11an1n08x5 FILLER_17_604 ();
 b15zdnd11an1n04x5 FILLER_17_612 ();
 b15zdnd00an1n01x5 FILLER_17_616 ();
 b15zdnd11an1n16x5 FILLER_17_625 ();
 b15zdnd11an1n04x5 FILLER_17_644 ();
 b15zdnd00an1n02x5 FILLER_17_648 ();
 b15zdnd00an1n01x5 FILLER_17_650 ();
 b15zdnd11an1n04x5 FILLER_17_654 ();
 b15zdnd11an1n04x5 FILLER_17_661 ();
 b15zdnd11an1n04x5 FILLER_17_668 ();
 b15zdnd11an1n04x5 FILLER_17_675 ();
 b15zdnd00an1n02x5 FILLER_17_679 ();
 b15zdnd00an1n01x5 FILLER_17_681 ();
 b15zdnd11an1n04x5 FILLER_17_685 ();
 b15zdnd00an1n01x5 FILLER_17_689 ();
 b15zdnd11an1n04x5 FILLER_17_693 ();
 b15zdnd11an1n04x5 FILLER_17_700 ();
 b15zdnd00an1n01x5 FILLER_17_704 ();
 b15zdnd11an1n64x5 FILLER_17_721 ();
 b15zdnd11an1n32x5 FILLER_17_785 ();
 b15zdnd00an1n02x5 FILLER_17_817 ();
 b15zdnd00an1n01x5 FILLER_17_819 ();
 b15zdnd11an1n04x5 FILLER_17_832 ();
 b15zdnd11an1n08x5 FILLER_17_847 ();
 b15zdnd11an1n04x5 FILLER_17_855 ();
 b15zdnd00an1n01x5 FILLER_17_859 ();
 b15zdnd11an1n64x5 FILLER_17_876 ();
 b15zdnd11an1n08x5 FILLER_17_940 ();
 b15zdnd11an1n08x5 FILLER_17_964 ();
 b15zdnd11an1n64x5 FILLER_17_978 ();
 b15zdnd11an1n64x5 FILLER_17_1042 ();
 b15zdnd11an1n64x5 FILLER_17_1106 ();
 b15zdnd11an1n16x5 FILLER_17_1170 ();
 b15zdnd11an1n08x5 FILLER_17_1186 ();
 b15zdnd00an1n02x5 FILLER_17_1194 ();
 b15zdnd00an1n01x5 FILLER_17_1196 ();
 b15zdnd11an1n04x5 FILLER_17_1207 ();
 b15zdnd11an1n64x5 FILLER_17_1215 ();
 b15zdnd11an1n16x5 FILLER_17_1279 ();
 b15zdnd11an1n04x5 FILLER_17_1295 ();
 b15zdnd00an1n02x5 FILLER_17_1299 ();
 b15zdnd00an1n01x5 FILLER_17_1301 ();
 b15zdnd11an1n64x5 FILLER_17_1306 ();
 b15zdnd11an1n16x5 FILLER_17_1370 ();
 b15zdnd11an1n08x5 FILLER_17_1386 ();
 b15zdnd00an1n01x5 FILLER_17_1394 ();
 b15zdnd11an1n64x5 FILLER_17_1405 ();
 b15zdnd11an1n16x5 FILLER_17_1469 ();
 b15zdnd00an1n01x5 FILLER_17_1485 ();
 b15zdnd11an1n16x5 FILLER_17_2257 ();
 b15zdnd11an1n08x5 FILLER_17_2273 ();
 b15zdnd00an1n02x5 FILLER_17_2281 ();
 b15zdnd00an1n01x5 FILLER_17_2283 ();
 b15zdnd11an1n64x5 FILLER_18_8 ();
 b15zdnd11an1n64x5 FILLER_18_72 ();
 b15zdnd11an1n64x5 FILLER_18_136 ();
 b15zdnd11an1n64x5 FILLER_18_200 ();
 b15zdnd11an1n64x5 FILLER_18_264 ();
 b15zdnd11an1n64x5 FILLER_18_328 ();
 b15zdnd11an1n64x5 FILLER_18_392 ();
 b15zdnd11an1n32x5 FILLER_18_456 ();
 b15zdnd11an1n16x5 FILLER_18_488 ();
 b15zdnd11an1n08x5 FILLER_18_504 ();
 b15zdnd11an1n04x5 FILLER_18_512 ();
 b15zdnd11an1n64x5 FILLER_18_547 ();
 b15zdnd11an1n32x5 FILLER_18_611 ();
 b15zdnd11an1n16x5 FILLER_18_643 ();
 b15zdnd11an1n08x5 FILLER_18_659 ();
 b15zdnd11an1n04x5 FILLER_18_667 ();
 b15zdnd00an1n02x5 FILLER_18_671 ();
 b15zdnd00an1n01x5 FILLER_18_673 ();
 b15zdnd11an1n04x5 FILLER_18_686 ();
 b15zdnd11an1n04x5 FILLER_18_693 ();
 b15zdnd11an1n04x5 FILLER_18_700 ();
 b15zdnd11an1n04x5 FILLER_18_707 ();
 b15zdnd00an1n02x5 FILLER_18_711 ();
 b15zdnd00an1n02x5 FILLER_18_716 ();
 b15zdnd11an1n08x5 FILLER_18_726 ();
 b15zdnd11an1n04x5 FILLER_18_734 ();
 b15zdnd00an1n02x5 FILLER_18_738 ();
 b15zdnd11an1n16x5 FILLER_18_753 ();
 b15zdnd11an1n04x5 FILLER_18_769 ();
 b15zdnd00an1n01x5 FILLER_18_773 ();
 b15zdnd11an1n64x5 FILLER_18_784 ();
 b15zdnd11an1n08x5 FILLER_18_848 ();
 b15zdnd11an1n04x5 FILLER_18_856 ();
 b15zdnd11an1n64x5 FILLER_18_876 ();
 b15zdnd00an1n02x5 FILLER_18_940 ();
 b15zdnd11an1n32x5 FILLER_18_984 ();
 b15zdnd11an1n16x5 FILLER_18_1016 ();
 b15zdnd11an1n04x5 FILLER_18_1032 ();
 b15zdnd00an1n01x5 FILLER_18_1036 ();
 b15zdnd11an1n08x5 FILLER_18_1047 ();
 b15zdnd00an1n02x5 FILLER_18_1055 ();
 b15zdnd11an1n64x5 FILLER_18_1063 ();
 b15zdnd11an1n32x5 FILLER_18_1127 ();
 b15zdnd11an1n16x5 FILLER_18_1159 ();
 b15zdnd11an1n08x5 FILLER_18_1175 ();
 b15zdnd11an1n04x5 FILLER_18_1183 ();
 b15zdnd00an1n01x5 FILLER_18_1187 ();
 b15zdnd11an1n04x5 FILLER_18_1219 ();
 b15zdnd11an1n64x5 FILLER_18_1233 ();
 b15zdnd11an1n16x5 FILLER_18_1297 ();
 b15zdnd11an1n04x5 FILLER_18_1313 ();
 b15zdnd00an1n02x5 FILLER_18_1317 ();
 b15zdnd00an1n01x5 FILLER_18_1319 ();
 b15zdnd11an1n32x5 FILLER_18_1332 ();
 b15zdnd11an1n16x5 FILLER_18_1364 ();
 b15zdnd11an1n08x5 FILLER_18_1380 ();
 b15zdnd11an1n04x5 FILLER_18_1388 ();
 b15zdnd00an1n01x5 FILLER_18_1392 ();
 b15zdnd11an1n04x5 FILLER_18_1406 ();
 b15zdnd11an1n32x5 FILLER_18_1423 ();
 b15zdnd11an1n16x5 FILLER_18_1455 ();
 b15zdnd11an1n04x5 FILLER_18_1471 ();
 b15zdnd00an1n02x5 FILLER_18_1475 ();
 b15zdnd00an1n01x5 FILLER_18_1477 ();
 b15zdnd11an1n08x5 FILLER_18_2265 ();
 b15zdnd00an1n02x5 FILLER_18_2273 ();
 b15zdnd00an1n01x5 FILLER_18_2275 ();
 b15zdnd11an1n64x5 FILLER_19_0 ();
 b15zdnd11an1n64x5 FILLER_19_64 ();
 b15zdnd11an1n64x5 FILLER_19_128 ();
 b15zdnd11an1n16x5 FILLER_19_192 ();
 b15zdnd11an1n04x5 FILLER_19_208 ();
 b15zdnd00an1n02x5 FILLER_19_212 ();
 b15zdnd00an1n01x5 FILLER_19_214 ();
 b15zdnd11an1n64x5 FILLER_19_231 ();
 b15zdnd11an1n64x5 FILLER_19_295 ();
 b15zdnd11an1n64x5 FILLER_19_359 ();
 b15zdnd11an1n64x5 FILLER_19_423 ();
 b15zdnd11an1n64x5 FILLER_19_487 ();
 b15zdnd11an1n64x5 FILLER_19_551 ();
 b15zdnd11an1n64x5 FILLER_19_615 ();
 b15zdnd11an1n16x5 FILLER_19_679 ();
 b15zdnd11an1n08x5 FILLER_19_695 ();
 b15zdnd11an1n04x5 FILLER_19_706 ();
 b15zdnd11an1n64x5 FILLER_19_713 ();
 b15zdnd11an1n16x5 FILLER_19_777 ();
 b15zdnd11an1n08x5 FILLER_19_793 ();
 b15zdnd00an1n02x5 FILLER_19_801 ();
 b15zdnd11an1n16x5 FILLER_19_845 ();
 b15zdnd00an1n02x5 FILLER_19_861 ();
 b15zdnd11an1n64x5 FILLER_19_905 ();
 b15zdnd11an1n32x5 FILLER_19_969 ();
 b15zdnd11an1n16x5 FILLER_19_1001 ();
 b15zdnd11an1n04x5 FILLER_19_1017 ();
 b15zdnd11an1n64x5 FILLER_19_1063 ();
 b15zdnd11an1n32x5 FILLER_19_1127 ();
 b15zdnd11an1n16x5 FILLER_19_1159 ();
 b15zdnd11an1n08x5 FILLER_19_1175 ();
 b15zdnd11an1n04x5 FILLER_19_1183 ();
 b15zdnd00an1n02x5 FILLER_19_1187 ();
 b15zdnd11an1n04x5 FILLER_19_1193 ();
 b15zdnd00an1n02x5 FILLER_19_1197 ();
 b15zdnd00an1n01x5 FILLER_19_1199 ();
 b15zdnd11an1n32x5 FILLER_19_1231 ();
 b15zdnd11an1n08x5 FILLER_19_1263 ();
 b15zdnd00an1n02x5 FILLER_19_1271 ();
 b15zdnd00an1n01x5 FILLER_19_1273 ();
 b15zdnd11an1n16x5 FILLER_19_1278 ();
 b15zdnd11an1n04x5 FILLER_19_1294 ();
 b15zdnd00an1n02x5 FILLER_19_1298 ();
 b15zdnd00an1n01x5 FILLER_19_1300 ();
 b15zdnd11an1n08x5 FILLER_19_1343 ();
 b15zdnd11an1n04x5 FILLER_19_1351 ();
 b15zdnd00an1n02x5 FILLER_19_1355 ();
 b15zdnd11an1n64x5 FILLER_19_1373 ();
 b15zdnd11an1n32x5 FILLER_19_1437 ();
 b15zdnd11an1n16x5 FILLER_19_1469 ();
 b15zdnd00an1n01x5 FILLER_19_1485 ();
 b15zdnd11an1n16x5 FILLER_19_2257 ();
 b15zdnd11an1n08x5 FILLER_19_2273 ();
 b15zdnd00an1n02x5 FILLER_19_2281 ();
 b15zdnd00an1n01x5 FILLER_19_2283 ();
 b15zdnd11an1n64x5 FILLER_20_8 ();
 b15zdnd11an1n64x5 FILLER_20_72 ();
 b15zdnd11an1n64x5 FILLER_20_136 ();
 b15zdnd11an1n64x5 FILLER_20_200 ();
 b15zdnd11an1n64x5 FILLER_20_264 ();
 b15zdnd11an1n64x5 FILLER_20_328 ();
 b15zdnd11an1n64x5 FILLER_20_392 ();
 b15zdnd11an1n64x5 FILLER_20_456 ();
 b15zdnd11an1n64x5 FILLER_20_520 ();
 b15zdnd11an1n64x5 FILLER_20_584 ();
 b15zdnd11an1n64x5 FILLER_20_648 ();
 b15zdnd11an1n04x5 FILLER_20_712 ();
 b15zdnd00an1n02x5 FILLER_20_716 ();
 b15zdnd11an1n64x5 FILLER_20_726 ();
 b15zdnd11an1n64x5 FILLER_20_790 ();
 b15zdnd11an1n16x5 FILLER_20_854 ();
 b15zdnd11an1n08x5 FILLER_20_870 ();
 b15zdnd11an1n04x5 FILLER_20_878 ();
 b15zdnd00an1n01x5 FILLER_20_882 ();
 b15zdnd11an1n32x5 FILLER_20_925 ();
 b15zdnd11an1n08x5 FILLER_20_957 ();
 b15zdnd11an1n04x5 FILLER_20_965 ();
 b15zdnd00an1n02x5 FILLER_20_969 ();
 b15zdnd00an1n01x5 FILLER_20_971 ();
 b15zdnd11an1n32x5 FILLER_20_984 ();
 b15zdnd11an1n16x5 FILLER_20_1016 ();
 b15zdnd11an1n04x5 FILLER_20_1032 ();
 b15zdnd00an1n01x5 FILLER_20_1036 ();
 b15zdnd11an1n16x5 FILLER_20_1047 ();
 b15zdnd11an1n04x5 FILLER_20_1063 ();
 b15zdnd00an1n02x5 FILLER_20_1067 ();
 b15zdnd00an1n01x5 FILLER_20_1069 ();
 b15zdnd11an1n64x5 FILLER_20_1112 ();
 b15zdnd11an1n64x5 FILLER_20_1176 ();
 b15zdnd11an1n64x5 FILLER_20_1240 ();
 b15zdnd00an1n02x5 FILLER_20_1304 ();
 b15zdnd11an1n16x5 FILLER_20_1322 ();
 b15zdnd00an1n02x5 FILLER_20_1338 ();
 b15zdnd11an1n64x5 FILLER_20_1356 ();
 b15zdnd11an1n32x5 FILLER_20_1420 ();
 b15zdnd11an1n16x5 FILLER_20_1452 ();
 b15zdnd11an1n08x5 FILLER_20_1468 ();
 b15zdnd00an1n02x5 FILLER_20_1476 ();
 b15zdnd11an1n08x5 FILLER_20_2265 ();
 b15zdnd00an1n02x5 FILLER_20_2273 ();
 b15zdnd00an1n01x5 FILLER_20_2275 ();
 b15zdnd11an1n64x5 FILLER_21_0 ();
 b15zdnd11an1n64x5 FILLER_21_64 ();
 b15zdnd11an1n64x5 FILLER_21_128 ();
 b15zdnd11an1n64x5 FILLER_21_192 ();
 b15zdnd11an1n64x5 FILLER_21_256 ();
 b15zdnd11an1n64x5 FILLER_21_320 ();
 b15zdnd11an1n64x5 FILLER_21_384 ();
 b15zdnd11an1n64x5 FILLER_21_448 ();
 b15zdnd11an1n64x5 FILLER_21_512 ();
 b15zdnd11an1n08x5 FILLER_21_576 ();
 b15zdnd00an1n01x5 FILLER_21_584 ();
 b15zdnd11an1n64x5 FILLER_21_601 ();
 b15zdnd11an1n64x5 FILLER_21_665 ();
 b15zdnd11an1n64x5 FILLER_21_729 ();
 b15zdnd11an1n64x5 FILLER_21_793 ();
 b15zdnd11an1n64x5 FILLER_21_857 ();
 b15zdnd11an1n32x5 FILLER_21_921 ();
 b15zdnd11an1n08x5 FILLER_21_953 ();
 b15zdnd11an1n04x5 FILLER_21_961 ();
 b15zdnd00an1n01x5 FILLER_21_965 ();
 b15zdnd11an1n32x5 FILLER_21_986 ();
 b15zdnd11an1n04x5 FILLER_21_1034 ();
 b15zdnd00an1n02x5 FILLER_21_1038 ();
 b15zdnd11an1n64x5 FILLER_21_1053 ();
 b15zdnd11an1n16x5 FILLER_21_1117 ();
 b15zdnd11an1n08x5 FILLER_21_1133 ();
 b15zdnd11an1n04x5 FILLER_21_1141 ();
 b15zdnd11an1n64x5 FILLER_21_1151 ();
 b15zdnd11an1n16x5 FILLER_21_1215 ();
 b15zdnd11an1n04x5 FILLER_21_1231 ();
 b15zdnd00an1n01x5 FILLER_21_1235 ();
 b15zdnd11an1n64x5 FILLER_21_1240 ();
 b15zdnd11an1n32x5 FILLER_21_1304 ();
 b15zdnd11an1n08x5 FILLER_21_1336 ();
 b15zdnd00an1n02x5 FILLER_21_1344 ();
 b15zdnd11an1n64x5 FILLER_21_1362 ();
 b15zdnd11an1n32x5 FILLER_21_1426 ();
 b15zdnd11an1n16x5 FILLER_21_1458 ();
 b15zdnd11an1n08x5 FILLER_21_1474 ();
 b15zdnd11an1n04x5 FILLER_21_1482 ();
 b15zdnd11an1n16x5 FILLER_21_2257 ();
 b15zdnd11an1n08x5 FILLER_21_2273 ();
 b15zdnd00an1n02x5 FILLER_21_2281 ();
 b15zdnd00an1n01x5 FILLER_21_2283 ();
 b15zdnd11an1n64x5 FILLER_22_8 ();
 b15zdnd11an1n64x5 FILLER_22_72 ();
 b15zdnd11an1n64x5 FILLER_22_136 ();
 b15zdnd11an1n64x5 FILLER_22_200 ();
 b15zdnd11an1n64x5 FILLER_22_264 ();
 b15zdnd11an1n64x5 FILLER_22_328 ();
 b15zdnd11an1n64x5 FILLER_22_392 ();
 b15zdnd11an1n64x5 FILLER_22_456 ();
 b15zdnd11an1n64x5 FILLER_22_520 ();
 b15zdnd11an1n64x5 FILLER_22_584 ();
 b15zdnd11an1n64x5 FILLER_22_648 ();
 b15zdnd11an1n04x5 FILLER_22_712 ();
 b15zdnd00an1n02x5 FILLER_22_716 ();
 b15zdnd11an1n64x5 FILLER_22_726 ();
 b15zdnd11an1n64x5 FILLER_22_790 ();
 b15zdnd11an1n64x5 FILLER_22_854 ();
 b15zdnd11an1n32x5 FILLER_22_918 ();
 b15zdnd11an1n16x5 FILLER_22_950 ();
 b15zdnd00an1n01x5 FILLER_22_966 ();
 b15zdnd11an1n32x5 FILLER_22_977 ();
 b15zdnd00an1n01x5 FILLER_22_1009 ();
 b15zdnd11an1n08x5 FILLER_22_1022 ();
 b15zdnd11an1n04x5 FILLER_22_1030 ();
 b15zdnd00an1n02x5 FILLER_22_1034 ();
 b15zdnd00an1n01x5 FILLER_22_1036 ();
 b15zdnd11an1n64x5 FILLER_22_1041 ();
 b15zdnd11an1n16x5 FILLER_22_1147 ();
 b15zdnd00an1n02x5 FILLER_22_1163 ();
 b15zdnd00an1n01x5 FILLER_22_1165 ();
 b15zdnd11an1n64x5 FILLER_22_1197 ();
 b15zdnd11an1n16x5 FILLER_22_1261 ();
 b15zdnd11an1n08x5 FILLER_22_1277 ();
 b15zdnd00an1n02x5 FILLER_22_1285 ();
 b15zdnd00an1n01x5 FILLER_22_1287 ();
 b15zdnd11an1n32x5 FILLER_22_1312 ();
 b15zdnd11an1n16x5 FILLER_22_1344 ();
 b15zdnd11an1n04x5 FILLER_22_1360 ();
 b15zdnd00an1n01x5 FILLER_22_1364 ();
 b15zdnd11an1n64x5 FILLER_22_1374 ();
 b15zdnd11an1n32x5 FILLER_22_1438 ();
 b15zdnd11an1n08x5 FILLER_22_1470 ();
 b15zdnd11an1n08x5 FILLER_22_2265 ();
 b15zdnd00an1n02x5 FILLER_22_2273 ();
 b15zdnd00an1n01x5 FILLER_22_2275 ();
 b15zdnd11an1n64x5 FILLER_23_0 ();
 b15zdnd11an1n64x5 FILLER_23_64 ();
 b15zdnd11an1n64x5 FILLER_23_128 ();
 b15zdnd11an1n64x5 FILLER_23_192 ();
 b15zdnd11an1n64x5 FILLER_23_256 ();
 b15zdnd11an1n16x5 FILLER_23_320 ();
 b15zdnd11an1n08x5 FILLER_23_336 ();
 b15zdnd11an1n04x5 FILLER_23_344 ();
 b15zdnd11an1n64x5 FILLER_23_352 ();
 b15zdnd11an1n64x5 FILLER_23_416 ();
 b15zdnd11an1n64x5 FILLER_23_480 ();
 b15zdnd11an1n64x5 FILLER_23_544 ();
 b15zdnd11an1n64x5 FILLER_23_608 ();
 b15zdnd11an1n64x5 FILLER_23_672 ();
 b15zdnd11an1n64x5 FILLER_23_736 ();
 b15zdnd11an1n64x5 FILLER_23_800 ();
 b15zdnd11an1n64x5 FILLER_23_864 ();
 b15zdnd11an1n64x5 FILLER_23_928 ();
 b15zdnd11an1n64x5 FILLER_23_992 ();
 b15zdnd11an1n64x5 FILLER_23_1056 ();
 b15zdnd11an1n64x5 FILLER_23_1120 ();
 b15zdnd11an1n16x5 FILLER_23_1184 ();
 b15zdnd11an1n04x5 FILLER_23_1200 ();
 b15zdnd11an1n16x5 FILLER_23_1212 ();
 b15zdnd11an1n08x5 FILLER_23_1228 ();
 b15zdnd00an1n02x5 FILLER_23_1236 ();
 b15zdnd11an1n64x5 FILLER_23_1242 ();
 b15zdnd11an1n32x5 FILLER_23_1306 ();
 b15zdnd11an1n16x5 FILLER_23_1338 ();
 b15zdnd00an1n02x5 FILLER_23_1354 ();
 b15zdnd00an1n01x5 FILLER_23_1356 ();
 b15zdnd11an1n64x5 FILLER_23_1368 ();
 b15zdnd11an1n32x5 FILLER_23_1432 ();
 b15zdnd11an1n16x5 FILLER_23_1464 ();
 b15zdnd11an1n04x5 FILLER_23_1480 ();
 b15zdnd00an1n02x5 FILLER_23_1484 ();
 b15zdnd11an1n16x5 FILLER_23_2257 ();
 b15zdnd11an1n08x5 FILLER_23_2273 ();
 b15zdnd00an1n02x5 FILLER_23_2281 ();
 b15zdnd00an1n01x5 FILLER_23_2283 ();
 b15zdnd11an1n64x5 FILLER_24_8 ();
 b15zdnd11an1n64x5 FILLER_24_72 ();
 b15zdnd11an1n08x5 FILLER_24_136 ();
 b15zdnd00an1n01x5 FILLER_24_144 ();
 b15zdnd11an1n64x5 FILLER_24_155 ();
 b15zdnd11an1n64x5 FILLER_24_219 ();
 b15zdnd11an1n64x5 FILLER_24_283 ();
 b15zdnd11an1n64x5 FILLER_24_347 ();
 b15zdnd11an1n64x5 FILLER_24_411 ();
 b15zdnd11an1n64x5 FILLER_24_475 ();
 b15zdnd11an1n64x5 FILLER_24_539 ();
 b15zdnd11an1n64x5 FILLER_24_603 ();
 b15zdnd11an1n32x5 FILLER_24_667 ();
 b15zdnd11an1n16x5 FILLER_24_699 ();
 b15zdnd00an1n02x5 FILLER_24_715 ();
 b15zdnd00an1n01x5 FILLER_24_717 ();
 b15zdnd11an1n64x5 FILLER_24_726 ();
 b15zdnd11an1n64x5 FILLER_24_790 ();
 b15zdnd11an1n64x5 FILLER_24_854 ();
 b15zdnd11an1n64x5 FILLER_24_918 ();
 b15zdnd11an1n64x5 FILLER_24_982 ();
 b15zdnd11an1n32x5 FILLER_24_1046 ();
 b15zdnd11an1n32x5 FILLER_24_1086 ();
 b15zdnd11an1n16x5 FILLER_24_1118 ();
 b15zdnd11an1n08x5 FILLER_24_1134 ();
 b15zdnd11an1n04x5 FILLER_24_1142 ();
 b15zdnd00an1n01x5 FILLER_24_1146 ();
 b15zdnd11an1n64x5 FILLER_24_1155 ();
 b15zdnd11an1n64x5 FILLER_24_1219 ();
 b15zdnd11an1n64x5 FILLER_24_1283 ();
 b15zdnd11an1n64x5 FILLER_24_1347 ();
 b15zdnd11an1n64x5 FILLER_24_1411 ();
 b15zdnd00an1n02x5 FILLER_24_1475 ();
 b15zdnd00an1n01x5 FILLER_24_1477 ();
 b15zdnd11an1n08x5 FILLER_24_2265 ();
 b15zdnd00an1n02x5 FILLER_24_2273 ();
 b15zdnd00an1n01x5 FILLER_24_2275 ();
 b15zdnd11an1n64x5 FILLER_25_0 ();
 b15zdnd11an1n64x5 FILLER_25_64 ();
 b15zdnd11an1n64x5 FILLER_25_128 ();
 b15zdnd11an1n64x5 FILLER_25_192 ();
 b15zdnd11an1n64x5 FILLER_25_256 ();
 b15zdnd11an1n64x5 FILLER_25_320 ();
 b15zdnd11an1n64x5 FILLER_25_384 ();
 b15zdnd11an1n64x5 FILLER_25_448 ();
 b15zdnd11an1n64x5 FILLER_25_512 ();
 b15zdnd11an1n64x5 FILLER_25_576 ();
 b15zdnd11an1n32x5 FILLER_25_640 ();
 b15zdnd11an1n08x5 FILLER_25_672 ();
 b15zdnd00an1n02x5 FILLER_25_680 ();
 b15zdnd00an1n01x5 FILLER_25_682 ();
 b15zdnd11an1n64x5 FILLER_25_725 ();
 b15zdnd11an1n64x5 FILLER_25_789 ();
 b15zdnd11an1n64x5 FILLER_25_853 ();
 b15zdnd11an1n64x5 FILLER_25_917 ();
 b15zdnd11an1n64x5 FILLER_25_981 ();
 b15zdnd11an1n64x5 FILLER_25_1045 ();
 b15zdnd11an1n64x5 FILLER_25_1109 ();
 b15zdnd11an1n64x5 FILLER_25_1173 ();
 b15zdnd11an1n64x5 FILLER_25_1237 ();
 b15zdnd11an1n64x5 FILLER_25_1301 ();
 b15zdnd11an1n64x5 FILLER_25_1365 ();
 b15zdnd11an1n32x5 FILLER_25_1429 ();
 b15zdnd11an1n16x5 FILLER_25_1461 ();
 b15zdnd11an1n08x5 FILLER_25_1477 ();
 b15zdnd00an1n01x5 FILLER_25_1485 ();
 b15zdnd11an1n16x5 FILLER_25_2257 ();
 b15zdnd11an1n08x5 FILLER_25_2273 ();
 b15zdnd00an1n02x5 FILLER_25_2281 ();
 b15zdnd00an1n01x5 FILLER_25_2283 ();
 b15zdnd11an1n64x5 FILLER_26_8 ();
 b15zdnd11an1n64x5 FILLER_26_72 ();
 b15zdnd11an1n64x5 FILLER_26_136 ();
 b15zdnd11an1n64x5 FILLER_26_200 ();
 b15zdnd11an1n64x5 FILLER_26_264 ();
 b15zdnd11an1n64x5 FILLER_26_328 ();
 b15zdnd11an1n64x5 FILLER_26_392 ();
 b15zdnd11an1n64x5 FILLER_26_456 ();
 b15zdnd11an1n64x5 FILLER_26_520 ();
 b15zdnd11an1n64x5 FILLER_26_584 ();
 b15zdnd11an1n64x5 FILLER_26_648 ();
 b15zdnd11an1n04x5 FILLER_26_712 ();
 b15zdnd00an1n02x5 FILLER_26_716 ();
 b15zdnd11an1n64x5 FILLER_26_726 ();
 b15zdnd11an1n64x5 FILLER_26_790 ();
 b15zdnd11an1n64x5 FILLER_26_854 ();
 b15zdnd11an1n64x5 FILLER_26_918 ();
 b15zdnd11an1n64x5 FILLER_26_982 ();
 b15zdnd11an1n64x5 FILLER_26_1046 ();
 b15zdnd11an1n64x5 FILLER_26_1110 ();
 b15zdnd11an1n64x5 FILLER_26_1174 ();
 b15zdnd11an1n16x5 FILLER_26_1238 ();
 b15zdnd11an1n04x5 FILLER_26_1254 ();
 b15zdnd00an1n02x5 FILLER_26_1258 ();
 b15zdnd11an1n64x5 FILLER_26_1273 ();
 b15zdnd11an1n64x5 FILLER_26_1337 ();
 b15zdnd11an1n64x5 FILLER_26_1401 ();
 b15zdnd11an1n08x5 FILLER_26_1465 ();
 b15zdnd11an1n04x5 FILLER_26_1473 ();
 b15zdnd00an1n01x5 FILLER_26_1477 ();
 b15zdnd11an1n08x5 FILLER_26_2265 ();
 b15zdnd00an1n02x5 FILLER_26_2273 ();
 b15zdnd00an1n01x5 FILLER_26_2275 ();
 b15zdnd11an1n64x5 FILLER_27_0 ();
 b15zdnd11an1n64x5 FILLER_27_64 ();
 b15zdnd11an1n64x5 FILLER_27_128 ();
 b15zdnd11an1n64x5 FILLER_27_192 ();
 b15zdnd11an1n64x5 FILLER_27_256 ();
 b15zdnd11an1n64x5 FILLER_27_320 ();
 b15zdnd11an1n64x5 FILLER_27_384 ();
 b15zdnd11an1n64x5 FILLER_27_448 ();
 b15zdnd11an1n64x5 FILLER_27_512 ();
 b15zdnd11an1n64x5 FILLER_27_576 ();
 b15zdnd11an1n64x5 FILLER_27_640 ();
 b15zdnd11an1n64x5 FILLER_27_704 ();
 b15zdnd11an1n64x5 FILLER_27_768 ();
 b15zdnd11an1n64x5 FILLER_27_832 ();
 b15zdnd11an1n64x5 FILLER_27_896 ();
 b15zdnd11an1n64x5 FILLER_27_960 ();
 b15zdnd11an1n32x5 FILLER_27_1024 ();
 b15zdnd11an1n16x5 FILLER_27_1056 ();
 b15zdnd11an1n04x5 FILLER_27_1072 ();
 b15zdnd00an1n02x5 FILLER_27_1076 ();
 b15zdnd00an1n01x5 FILLER_27_1078 ();
 b15zdnd11an1n64x5 FILLER_27_1095 ();
 b15zdnd11an1n16x5 FILLER_27_1159 ();
 b15zdnd11an1n08x5 FILLER_27_1175 ();
 b15zdnd11an1n04x5 FILLER_27_1183 ();
 b15zdnd00an1n01x5 FILLER_27_1187 ();
 b15zdnd11an1n64x5 FILLER_27_1201 ();
 b15zdnd11an1n64x5 FILLER_27_1265 ();
 b15zdnd11an1n64x5 FILLER_27_1329 ();
 b15zdnd11an1n64x5 FILLER_27_1393 ();
 b15zdnd11an1n16x5 FILLER_27_1457 ();
 b15zdnd11an1n08x5 FILLER_27_1473 ();
 b15zdnd11an1n04x5 FILLER_27_1481 ();
 b15zdnd00an1n01x5 FILLER_27_1485 ();
 b15zdnd11an1n16x5 FILLER_27_2257 ();
 b15zdnd11an1n08x5 FILLER_27_2273 ();
 b15zdnd00an1n02x5 FILLER_27_2281 ();
 b15zdnd00an1n01x5 FILLER_27_2283 ();
 b15zdnd11an1n64x5 FILLER_28_8 ();
 b15zdnd11an1n64x5 FILLER_28_72 ();
 b15zdnd11an1n64x5 FILLER_28_136 ();
 b15zdnd11an1n64x5 FILLER_28_200 ();
 b15zdnd11an1n64x5 FILLER_28_264 ();
 b15zdnd11an1n64x5 FILLER_28_328 ();
 b15zdnd11an1n64x5 FILLER_28_392 ();
 b15zdnd11an1n64x5 FILLER_28_456 ();
 b15zdnd11an1n64x5 FILLER_28_520 ();
 b15zdnd11an1n64x5 FILLER_28_584 ();
 b15zdnd11an1n64x5 FILLER_28_648 ();
 b15zdnd11an1n04x5 FILLER_28_712 ();
 b15zdnd00an1n02x5 FILLER_28_716 ();
 b15zdnd11an1n64x5 FILLER_28_726 ();
 b15zdnd11an1n64x5 FILLER_28_790 ();
 b15zdnd11an1n64x5 FILLER_28_854 ();
 b15zdnd11an1n64x5 FILLER_28_918 ();
 b15zdnd11an1n64x5 FILLER_28_982 ();
 b15zdnd11an1n64x5 FILLER_28_1046 ();
 b15zdnd11an1n64x5 FILLER_28_1110 ();
 b15zdnd11an1n64x5 FILLER_28_1174 ();
 b15zdnd11an1n64x5 FILLER_28_1238 ();
 b15zdnd11an1n64x5 FILLER_28_1302 ();
 b15zdnd11an1n64x5 FILLER_28_1366 ();
 b15zdnd11an1n32x5 FILLER_28_1430 ();
 b15zdnd11an1n16x5 FILLER_28_1462 ();
 b15zdnd11an1n08x5 FILLER_28_2265 ();
 b15zdnd00an1n02x5 FILLER_28_2273 ();
 b15zdnd00an1n01x5 FILLER_28_2275 ();
 b15zdnd11an1n64x5 FILLER_29_0 ();
 b15zdnd11an1n64x5 FILLER_29_64 ();
 b15zdnd11an1n64x5 FILLER_29_128 ();
 b15zdnd11an1n64x5 FILLER_29_192 ();
 b15zdnd11an1n64x5 FILLER_29_256 ();
 b15zdnd11an1n64x5 FILLER_29_320 ();
 b15zdnd11an1n64x5 FILLER_29_384 ();
 b15zdnd11an1n64x5 FILLER_29_448 ();
 b15zdnd11an1n64x5 FILLER_29_512 ();
 b15zdnd11an1n64x5 FILLER_29_576 ();
 b15zdnd11an1n64x5 FILLER_29_640 ();
 b15zdnd11an1n64x5 FILLER_29_704 ();
 b15zdnd11an1n32x5 FILLER_29_768 ();
 b15zdnd11an1n16x5 FILLER_29_800 ();
 b15zdnd11an1n08x5 FILLER_29_816 ();
 b15zdnd11an1n04x5 FILLER_29_824 ();
 b15zdnd00an1n01x5 FILLER_29_828 ();
 b15zdnd11an1n64x5 FILLER_29_871 ();
 b15zdnd11an1n64x5 FILLER_29_935 ();
 b15zdnd11an1n64x5 FILLER_29_999 ();
 b15zdnd11an1n64x5 FILLER_29_1063 ();
 b15zdnd11an1n64x5 FILLER_29_1127 ();
 b15zdnd11an1n64x5 FILLER_29_1191 ();
 b15zdnd11an1n64x5 FILLER_29_1255 ();
 b15zdnd11an1n64x5 FILLER_29_1319 ();
 b15zdnd11an1n64x5 FILLER_29_1383 ();
 b15zdnd11an1n32x5 FILLER_29_1447 ();
 b15zdnd11an1n04x5 FILLER_29_1479 ();
 b15zdnd00an1n02x5 FILLER_29_1483 ();
 b15zdnd00an1n01x5 FILLER_29_1485 ();
 b15zdnd11an1n16x5 FILLER_29_2257 ();
 b15zdnd11an1n08x5 FILLER_29_2273 ();
 b15zdnd00an1n02x5 FILLER_29_2281 ();
 b15zdnd00an1n01x5 FILLER_29_2283 ();
 b15zdnd11an1n64x5 FILLER_30_8 ();
 b15zdnd11an1n64x5 FILLER_30_72 ();
 b15zdnd11an1n64x5 FILLER_30_136 ();
 b15zdnd11an1n64x5 FILLER_30_200 ();
 b15zdnd11an1n64x5 FILLER_30_264 ();
 b15zdnd11an1n64x5 FILLER_30_328 ();
 b15zdnd11an1n64x5 FILLER_30_392 ();
 b15zdnd11an1n64x5 FILLER_30_456 ();
 b15zdnd11an1n64x5 FILLER_30_520 ();
 b15zdnd11an1n64x5 FILLER_30_584 ();
 b15zdnd11an1n64x5 FILLER_30_648 ();
 b15zdnd11an1n04x5 FILLER_30_712 ();
 b15zdnd00an1n02x5 FILLER_30_716 ();
 b15zdnd11an1n64x5 FILLER_30_726 ();
 b15zdnd11an1n64x5 FILLER_30_790 ();
 b15zdnd11an1n32x5 FILLER_30_854 ();
 b15zdnd11an1n16x5 FILLER_30_886 ();
 b15zdnd11an1n04x5 FILLER_30_902 ();
 b15zdnd00an1n02x5 FILLER_30_906 ();
 b15zdnd00an1n01x5 FILLER_30_908 ();
 b15zdnd11an1n64x5 FILLER_30_917 ();
 b15zdnd11an1n64x5 FILLER_30_981 ();
 b15zdnd11an1n64x5 FILLER_30_1045 ();
 b15zdnd11an1n64x5 FILLER_30_1109 ();
 b15zdnd11an1n64x5 FILLER_30_1173 ();
 b15zdnd11an1n64x5 FILLER_30_1237 ();
 b15zdnd11an1n64x5 FILLER_30_1301 ();
 b15zdnd11an1n64x5 FILLER_30_1365 ();
 b15zdnd11an1n32x5 FILLER_30_1429 ();
 b15zdnd11an1n16x5 FILLER_30_1461 ();
 b15zdnd00an1n01x5 FILLER_30_1477 ();
 b15zdnd11an1n08x5 FILLER_30_2265 ();
 b15zdnd00an1n02x5 FILLER_30_2273 ();
 b15zdnd00an1n01x5 FILLER_30_2275 ();
 b15zdnd11an1n64x5 FILLER_31_0 ();
 b15zdnd11an1n64x5 FILLER_31_64 ();
 b15zdnd11an1n64x5 FILLER_31_128 ();
 b15zdnd11an1n64x5 FILLER_31_192 ();
 b15zdnd11an1n64x5 FILLER_31_256 ();
 b15zdnd11an1n64x5 FILLER_31_320 ();
 b15zdnd11an1n64x5 FILLER_31_384 ();
 b15zdnd11an1n64x5 FILLER_31_448 ();
 b15zdnd11an1n64x5 FILLER_31_512 ();
 b15zdnd11an1n64x5 FILLER_31_576 ();
 b15zdnd11an1n64x5 FILLER_31_640 ();
 b15zdnd11an1n64x5 FILLER_31_704 ();
 b15zdnd11an1n64x5 FILLER_31_768 ();
 b15zdnd11an1n64x5 FILLER_31_832 ();
 b15zdnd11an1n64x5 FILLER_31_896 ();
 b15zdnd11an1n64x5 FILLER_31_960 ();
 b15zdnd11an1n64x5 FILLER_31_1024 ();
 b15zdnd11an1n64x5 FILLER_31_1088 ();
 b15zdnd11an1n64x5 FILLER_31_1152 ();
 b15zdnd11an1n64x5 FILLER_31_1216 ();
 b15zdnd11an1n64x5 FILLER_31_1280 ();
 b15zdnd11an1n64x5 FILLER_31_1344 ();
 b15zdnd11an1n64x5 FILLER_31_1408 ();
 b15zdnd11an1n08x5 FILLER_31_1472 ();
 b15zdnd11an1n04x5 FILLER_31_1480 ();
 b15zdnd00an1n02x5 FILLER_31_1484 ();
 b15zdnd11an1n16x5 FILLER_31_2257 ();
 b15zdnd11an1n08x5 FILLER_31_2273 ();
 b15zdnd00an1n02x5 FILLER_31_2281 ();
 b15zdnd00an1n01x5 FILLER_31_2283 ();
 b15zdnd11an1n64x5 FILLER_32_8 ();
 b15zdnd11an1n64x5 FILLER_32_72 ();
 b15zdnd11an1n64x5 FILLER_32_136 ();
 b15zdnd11an1n64x5 FILLER_32_200 ();
 b15zdnd11an1n64x5 FILLER_32_264 ();
 b15zdnd11an1n64x5 FILLER_32_328 ();
 b15zdnd11an1n64x5 FILLER_32_392 ();
 b15zdnd11an1n64x5 FILLER_32_456 ();
 b15zdnd11an1n16x5 FILLER_32_520 ();
 b15zdnd11an1n64x5 FILLER_32_578 ();
 b15zdnd11an1n64x5 FILLER_32_642 ();
 b15zdnd11an1n08x5 FILLER_32_706 ();
 b15zdnd11an1n04x5 FILLER_32_714 ();
 b15zdnd00an1n02x5 FILLER_32_726 ();
 b15zdnd11an1n64x5 FILLER_32_770 ();
 b15zdnd11an1n64x5 FILLER_32_834 ();
 b15zdnd11an1n64x5 FILLER_32_898 ();
 b15zdnd11an1n64x5 FILLER_32_962 ();
 b15zdnd11an1n64x5 FILLER_32_1026 ();
 b15zdnd11an1n64x5 FILLER_32_1090 ();
 b15zdnd11an1n64x5 FILLER_32_1154 ();
 b15zdnd11an1n64x5 FILLER_32_1218 ();
 b15zdnd11an1n64x5 FILLER_32_1282 ();
 b15zdnd11an1n64x5 FILLER_32_1346 ();
 b15zdnd11an1n64x5 FILLER_32_1410 ();
 b15zdnd11an1n04x5 FILLER_32_1474 ();
 b15zdnd11an1n08x5 FILLER_32_2265 ();
 b15zdnd00an1n02x5 FILLER_32_2273 ();
 b15zdnd00an1n01x5 FILLER_32_2275 ();
 b15zdnd11an1n64x5 FILLER_33_0 ();
 b15zdnd11an1n64x5 FILLER_33_64 ();
 b15zdnd11an1n64x5 FILLER_33_128 ();
 b15zdnd11an1n64x5 FILLER_33_192 ();
 b15zdnd11an1n64x5 FILLER_33_256 ();
 b15zdnd11an1n64x5 FILLER_33_320 ();
 b15zdnd11an1n32x5 FILLER_33_384 ();
 b15zdnd11an1n16x5 FILLER_33_416 ();
 b15zdnd11an1n64x5 FILLER_33_463 ();
 b15zdnd11an1n64x5 FILLER_33_527 ();
 b15zdnd11an1n08x5 FILLER_33_591 ();
 b15zdnd00an1n02x5 FILLER_33_599 ();
 b15zdnd11an1n64x5 FILLER_33_617 ();
 b15zdnd11an1n64x5 FILLER_33_681 ();
 b15zdnd11an1n64x5 FILLER_33_745 ();
 b15zdnd11an1n64x5 FILLER_33_809 ();
 b15zdnd11an1n64x5 FILLER_33_873 ();
 b15zdnd11an1n64x5 FILLER_33_937 ();
 b15zdnd11an1n64x5 FILLER_33_1001 ();
 b15zdnd11an1n64x5 FILLER_33_1065 ();
 b15zdnd11an1n64x5 FILLER_33_1129 ();
 b15zdnd11an1n64x5 FILLER_33_1193 ();
 b15zdnd11an1n64x5 FILLER_33_1257 ();
 b15zdnd11an1n64x5 FILLER_33_1321 ();
 b15zdnd11an1n64x5 FILLER_33_1385 ();
 b15zdnd11an1n32x5 FILLER_33_1449 ();
 b15zdnd11an1n04x5 FILLER_33_1481 ();
 b15zdnd00an1n01x5 FILLER_33_1485 ();
 b15zdnd11an1n16x5 FILLER_33_2257 ();
 b15zdnd11an1n08x5 FILLER_33_2273 ();
 b15zdnd00an1n02x5 FILLER_33_2281 ();
 b15zdnd00an1n01x5 FILLER_33_2283 ();
 b15zdnd11an1n64x5 FILLER_34_8 ();
 b15zdnd11an1n64x5 FILLER_34_72 ();
 b15zdnd11an1n64x5 FILLER_34_136 ();
 b15zdnd11an1n64x5 FILLER_34_200 ();
 b15zdnd11an1n64x5 FILLER_34_264 ();
 b15zdnd11an1n64x5 FILLER_34_328 ();
 b15zdnd11an1n64x5 FILLER_34_392 ();
 b15zdnd11an1n64x5 FILLER_34_456 ();
 b15zdnd11an1n64x5 FILLER_34_520 ();
 b15zdnd11an1n64x5 FILLER_34_584 ();
 b15zdnd11an1n64x5 FILLER_34_648 ();
 b15zdnd11an1n04x5 FILLER_34_712 ();
 b15zdnd00an1n02x5 FILLER_34_716 ();
 b15zdnd11an1n64x5 FILLER_34_726 ();
 b15zdnd11an1n64x5 FILLER_34_790 ();
 b15zdnd11an1n64x5 FILLER_34_854 ();
 b15zdnd11an1n64x5 FILLER_34_918 ();
 b15zdnd11an1n64x5 FILLER_34_982 ();
 b15zdnd11an1n64x5 FILLER_34_1046 ();
 b15zdnd11an1n64x5 FILLER_34_1110 ();
 b15zdnd11an1n64x5 FILLER_34_1174 ();
 b15zdnd11an1n64x5 FILLER_34_1238 ();
 b15zdnd11an1n64x5 FILLER_34_1302 ();
 b15zdnd11an1n64x5 FILLER_34_1366 ();
 b15zdnd11an1n32x5 FILLER_34_1430 ();
 b15zdnd11an1n16x5 FILLER_34_1462 ();
 b15zdnd11an1n08x5 FILLER_34_2265 ();
 b15zdnd00an1n02x5 FILLER_34_2273 ();
 b15zdnd00an1n01x5 FILLER_34_2275 ();
 b15zdnd11an1n64x5 FILLER_35_0 ();
 b15zdnd11an1n64x5 FILLER_35_64 ();
 b15zdnd11an1n64x5 FILLER_35_128 ();
 b15zdnd11an1n64x5 FILLER_35_192 ();
 b15zdnd11an1n64x5 FILLER_35_256 ();
 b15zdnd11an1n64x5 FILLER_35_320 ();
 b15zdnd11an1n64x5 FILLER_35_384 ();
 b15zdnd11an1n64x5 FILLER_35_448 ();
 b15zdnd11an1n64x5 FILLER_35_512 ();
 b15zdnd11an1n64x5 FILLER_35_576 ();
 b15zdnd11an1n64x5 FILLER_35_640 ();
 b15zdnd11an1n64x5 FILLER_35_704 ();
 b15zdnd11an1n64x5 FILLER_35_768 ();
 b15zdnd11an1n64x5 FILLER_35_832 ();
 b15zdnd11an1n64x5 FILLER_35_896 ();
 b15zdnd11an1n64x5 FILLER_35_960 ();
 b15zdnd11an1n64x5 FILLER_35_1024 ();
 b15zdnd11an1n64x5 FILLER_35_1088 ();
 b15zdnd11an1n64x5 FILLER_35_1152 ();
 b15zdnd11an1n64x5 FILLER_35_1216 ();
 b15zdnd11an1n64x5 FILLER_35_1280 ();
 b15zdnd11an1n64x5 FILLER_35_1344 ();
 b15zdnd11an1n64x5 FILLER_35_1408 ();
 b15zdnd11an1n08x5 FILLER_35_1472 ();
 b15zdnd11an1n04x5 FILLER_35_1480 ();
 b15zdnd00an1n02x5 FILLER_35_1484 ();
 b15zdnd11an1n16x5 FILLER_35_2257 ();
 b15zdnd11an1n08x5 FILLER_35_2273 ();
 b15zdnd00an1n02x5 FILLER_35_2281 ();
 b15zdnd00an1n01x5 FILLER_35_2283 ();
 b15zdnd11an1n64x5 FILLER_36_8 ();
 b15zdnd11an1n64x5 FILLER_36_72 ();
 b15zdnd11an1n64x5 FILLER_36_136 ();
 b15zdnd11an1n64x5 FILLER_36_200 ();
 b15zdnd11an1n64x5 FILLER_36_264 ();
 b15zdnd11an1n64x5 FILLER_36_328 ();
 b15zdnd11an1n64x5 FILLER_36_392 ();
 b15zdnd11an1n64x5 FILLER_36_456 ();
 b15zdnd11an1n64x5 FILLER_36_520 ();
 b15zdnd11an1n32x5 FILLER_36_584 ();
 b15zdnd11an1n08x5 FILLER_36_616 ();
 b15zdnd11an1n04x5 FILLER_36_624 ();
 b15zdnd11an1n32x5 FILLER_36_670 ();
 b15zdnd11an1n16x5 FILLER_36_702 ();
 b15zdnd11an1n64x5 FILLER_36_726 ();
 b15zdnd11an1n64x5 FILLER_36_790 ();
 b15zdnd11an1n64x5 FILLER_36_854 ();
 b15zdnd11an1n64x5 FILLER_36_918 ();
 b15zdnd11an1n64x5 FILLER_36_982 ();
 b15zdnd11an1n64x5 FILLER_36_1046 ();
 b15zdnd11an1n64x5 FILLER_36_1110 ();
 b15zdnd11an1n64x5 FILLER_36_1174 ();
 b15zdnd11an1n64x5 FILLER_36_1238 ();
 b15zdnd11an1n64x5 FILLER_36_1302 ();
 b15zdnd11an1n64x5 FILLER_36_1366 ();
 b15zdnd11an1n32x5 FILLER_36_1430 ();
 b15zdnd11an1n16x5 FILLER_36_1462 ();
 b15zdnd11an1n08x5 FILLER_36_2265 ();
 b15zdnd00an1n02x5 FILLER_36_2273 ();
 b15zdnd00an1n01x5 FILLER_36_2275 ();
 b15zdnd11an1n64x5 FILLER_37_0 ();
 b15zdnd11an1n64x5 FILLER_37_64 ();
 b15zdnd11an1n64x5 FILLER_37_128 ();
 b15zdnd11an1n64x5 FILLER_37_192 ();
 b15zdnd11an1n64x5 FILLER_37_256 ();
 b15zdnd11an1n64x5 FILLER_37_320 ();
 b15zdnd11an1n64x5 FILLER_37_384 ();
 b15zdnd11an1n64x5 FILLER_37_448 ();
 b15zdnd11an1n64x5 FILLER_37_512 ();
 b15zdnd11an1n64x5 FILLER_37_576 ();
 b15zdnd11an1n64x5 FILLER_37_640 ();
 b15zdnd11an1n64x5 FILLER_37_704 ();
 b15zdnd11an1n64x5 FILLER_37_768 ();
 b15zdnd11an1n64x5 FILLER_37_832 ();
 b15zdnd11an1n64x5 FILLER_37_896 ();
 b15zdnd11an1n64x5 FILLER_37_960 ();
 b15zdnd11an1n64x5 FILLER_37_1024 ();
 b15zdnd11an1n64x5 FILLER_37_1088 ();
 b15zdnd11an1n64x5 FILLER_37_1152 ();
 b15zdnd11an1n64x5 FILLER_37_1216 ();
 b15zdnd11an1n64x5 FILLER_37_1280 ();
 b15zdnd11an1n64x5 FILLER_37_1344 ();
 b15zdnd11an1n64x5 FILLER_37_1408 ();
 b15zdnd11an1n08x5 FILLER_37_1472 ();
 b15zdnd11an1n04x5 FILLER_37_1480 ();
 b15zdnd00an1n02x5 FILLER_37_1484 ();
 b15zdnd11an1n16x5 FILLER_37_2257 ();
 b15zdnd11an1n08x5 FILLER_37_2273 ();
 b15zdnd00an1n02x5 FILLER_37_2281 ();
 b15zdnd00an1n01x5 FILLER_37_2283 ();
 b15zdnd11an1n64x5 FILLER_38_8 ();
 b15zdnd11an1n64x5 FILLER_38_72 ();
 b15zdnd11an1n64x5 FILLER_38_136 ();
 b15zdnd11an1n64x5 FILLER_38_200 ();
 b15zdnd11an1n64x5 FILLER_38_264 ();
 b15zdnd11an1n64x5 FILLER_38_328 ();
 b15zdnd11an1n64x5 FILLER_38_392 ();
 b15zdnd11an1n64x5 FILLER_38_456 ();
 b15zdnd11an1n64x5 FILLER_38_520 ();
 b15zdnd11an1n64x5 FILLER_38_584 ();
 b15zdnd11an1n64x5 FILLER_38_648 ();
 b15zdnd11an1n04x5 FILLER_38_712 ();
 b15zdnd00an1n02x5 FILLER_38_716 ();
 b15zdnd11an1n64x5 FILLER_38_726 ();
 b15zdnd11an1n64x5 FILLER_38_790 ();
 b15zdnd11an1n04x5 FILLER_38_854 ();
 b15zdnd11an1n64x5 FILLER_38_900 ();
 b15zdnd11an1n64x5 FILLER_38_964 ();
 b15zdnd11an1n64x5 FILLER_38_1028 ();
 b15zdnd11an1n64x5 FILLER_38_1092 ();
 b15zdnd11an1n64x5 FILLER_38_1156 ();
 b15zdnd11an1n64x5 FILLER_38_1220 ();
 b15zdnd11an1n64x5 FILLER_38_1284 ();
 b15zdnd11an1n64x5 FILLER_38_1348 ();
 b15zdnd11an1n64x5 FILLER_38_1412 ();
 b15zdnd00an1n02x5 FILLER_38_1476 ();
 b15zdnd11an1n08x5 FILLER_38_2265 ();
 b15zdnd00an1n02x5 FILLER_38_2273 ();
 b15zdnd00an1n01x5 FILLER_38_2275 ();
 b15zdnd11an1n64x5 FILLER_39_0 ();
 b15zdnd11an1n64x5 FILLER_39_64 ();
 b15zdnd11an1n64x5 FILLER_39_128 ();
 b15zdnd11an1n64x5 FILLER_39_192 ();
 b15zdnd11an1n64x5 FILLER_39_256 ();
 b15zdnd11an1n64x5 FILLER_39_320 ();
 b15zdnd11an1n64x5 FILLER_39_384 ();
 b15zdnd11an1n64x5 FILLER_39_448 ();
 b15zdnd11an1n64x5 FILLER_39_512 ();
 b15zdnd11an1n64x5 FILLER_39_576 ();
 b15zdnd11an1n32x5 FILLER_39_640 ();
 b15zdnd11an1n16x5 FILLER_39_672 ();
 b15zdnd11an1n04x5 FILLER_39_688 ();
 b15zdnd00an1n02x5 FILLER_39_692 ();
 b15zdnd00an1n01x5 FILLER_39_694 ();
 b15zdnd11an1n64x5 FILLER_39_737 ();
 b15zdnd11an1n64x5 FILLER_39_801 ();
 b15zdnd11an1n64x5 FILLER_39_865 ();
 b15zdnd11an1n64x5 FILLER_39_929 ();
 b15zdnd11an1n64x5 FILLER_39_993 ();
 b15zdnd11an1n64x5 FILLER_39_1057 ();
 b15zdnd11an1n16x5 FILLER_39_1121 ();
 b15zdnd11an1n64x5 FILLER_39_1151 ();
 b15zdnd11an1n64x5 FILLER_39_1215 ();
 b15zdnd11an1n64x5 FILLER_39_1279 ();
 b15zdnd11an1n64x5 FILLER_39_1343 ();
 b15zdnd11an1n64x5 FILLER_39_1407 ();
 b15zdnd11an1n08x5 FILLER_39_1471 ();
 b15zdnd11an1n04x5 FILLER_39_1479 ();
 b15zdnd00an1n02x5 FILLER_39_1483 ();
 b15zdnd00an1n01x5 FILLER_39_1485 ();
 b15zdnd11an1n16x5 FILLER_39_2257 ();
 b15zdnd11an1n08x5 FILLER_39_2273 ();
 b15zdnd00an1n02x5 FILLER_39_2281 ();
 b15zdnd00an1n01x5 FILLER_39_2283 ();
 b15zdnd11an1n64x5 FILLER_40_8 ();
 b15zdnd11an1n64x5 FILLER_40_72 ();
 b15zdnd11an1n64x5 FILLER_40_136 ();
 b15zdnd11an1n64x5 FILLER_40_200 ();
 b15zdnd11an1n64x5 FILLER_40_264 ();
 b15zdnd11an1n64x5 FILLER_40_328 ();
 b15zdnd11an1n64x5 FILLER_40_392 ();
 b15zdnd11an1n64x5 FILLER_40_456 ();
 b15zdnd11an1n64x5 FILLER_40_520 ();
 b15zdnd11an1n64x5 FILLER_40_584 ();
 b15zdnd11an1n64x5 FILLER_40_648 ();
 b15zdnd11an1n04x5 FILLER_40_712 ();
 b15zdnd00an1n02x5 FILLER_40_716 ();
 b15zdnd11an1n32x5 FILLER_40_726 ();
 b15zdnd11an1n08x5 FILLER_40_758 ();
 b15zdnd00an1n02x5 FILLER_40_766 ();
 b15zdnd00an1n01x5 FILLER_40_768 ();
 b15zdnd11an1n64x5 FILLER_40_811 ();
 b15zdnd11an1n64x5 FILLER_40_875 ();
 b15zdnd11an1n64x5 FILLER_40_939 ();
 b15zdnd11an1n64x5 FILLER_40_1003 ();
 b15zdnd11an1n64x5 FILLER_40_1067 ();
 b15zdnd11an1n64x5 FILLER_40_1131 ();
 b15zdnd11an1n64x5 FILLER_40_1195 ();
 b15zdnd11an1n64x5 FILLER_40_1259 ();
 b15zdnd11an1n64x5 FILLER_40_1323 ();
 b15zdnd11an1n64x5 FILLER_40_1387 ();
 b15zdnd11an1n16x5 FILLER_40_1451 ();
 b15zdnd11an1n08x5 FILLER_40_1467 ();
 b15zdnd00an1n02x5 FILLER_40_1475 ();
 b15zdnd00an1n01x5 FILLER_40_1477 ();
 b15zdnd11an1n08x5 FILLER_40_2265 ();
 b15zdnd00an1n02x5 FILLER_40_2273 ();
 b15zdnd00an1n01x5 FILLER_40_2275 ();
 b15zdnd11an1n64x5 FILLER_41_0 ();
 b15zdnd11an1n64x5 FILLER_41_64 ();
 b15zdnd11an1n64x5 FILLER_41_128 ();
 b15zdnd11an1n64x5 FILLER_41_192 ();
 b15zdnd11an1n64x5 FILLER_41_256 ();
 b15zdnd11an1n32x5 FILLER_41_320 ();
 b15zdnd11an1n16x5 FILLER_41_352 ();
 b15zdnd11an1n08x5 FILLER_41_368 ();
 b15zdnd11an1n04x5 FILLER_41_376 ();
 b15zdnd00an1n02x5 FILLER_41_380 ();
 b15zdnd11an1n64x5 FILLER_41_413 ();
 b15zdnd11an1n64x5 FILLER_41_477 ();
 b15zdnd11an1n64x5 FILLER_41_541 ();
 b15zdnd11an1n64x5 FILLER_41_605 ();
 b15zdnd11an1n64x5 FILLER_41_669 ();
 b15zdnd11an1n64x5 FILLER_41_733 ();
 b15zdnd11an1n32x5 FILLER_41_797 ();
 b15zdnd11an1n08x5 FILLER_41_829 ();
 b15zdnd11an1n04x5 FILLER_41_837 ();
 b15zdnd11an1n64x5 FILLER_41_883 ();
 b15zdnd11an1n64x5 FILLER_41_947 ();
 b15zdnd11an1n64x5 FILLER_41_1011 ();
 b15zdnd11an1n64x5 FILLER_41_1075 ();
 b15zdnd11an1n64x5 FILLER_41_1139 ();
 b15zdnd11an1n64x5 FILLER_41_1203 ();
 b15zdnd11an1n64x5 FILLER_41_1267 ();
 b15zdnd11an1n64x5 FILLER_41_1331 ();
 b15zdnd11an1n64x5 FILLER_41_1395 ();
 b15zdnd11an1n16x5 FILLER_41_1459 ();
 b15zdnd11an1n08x5 FILLER_41_1475 ();
 b15zdnd00an1n02x5 FILLER_41_1483 ();
 b15zdnd00an1n01x5 FILLER_41_1485 ();
 b15zdnd11an1n16x5 FILLER_41_2257 ();
 b15zdnd11an1n08x5 FILLER_41_2273 ();
 b15zdnd00an1n02x5 FILLER_41_2281 ();
 b15zdnd00an1n01x5 FILLER_41_2283 ();
 b15zdnd11an1n64x5 FILLER_42_8 ();
 b15zdnd11an1n64x5 FILLER_42_72 ();
 b15zdnd11an1n64x5 FILLER_42_136 ();
 b15zdnd11an1n64x5 FILLER_42_200 ();
 b15zdnd11an1n64x5 FILLER_42_264 ();
 b15zdnd11an1n64x5 FILLER_42_328 ();
 b15zdnd11an1n64x5 FILLER_42_392 ();
 b15zdnd11an1n64x5 FILLER_42_456 ();
 b15zdnd11an1n64x5 FILLER_42_520 ();
 b15zdnd11an1n64x5 FILLER_42_584 ();
 b15zdnd11an1n64x5 FILLER_42_648 ();
 b15zdnd11an1n04x5 FILLER_42_712 ();
 b15zdnd00an1n02x5 FILLER_42_716 ();
 b15zdnd11an1n64x5 FILLER_42_726 ();
 b15zdnd11an1n64x5 FILLER_42_790 ();
 b15zdnd11an1n64x5 FILLER_42_854 ();
 b15zdnd11an1n32x5 FILLER_42_918 ();
 b15zdnd11an1n16x5 FILLER_42_950 ();
 b15zdnd00an1n01x5 FILLER_42_966 ();
 b15zdnd11an1n64x5 FILLER_42_1009 ();
 b15zdnd11an1n16x5 FILLER_42_1073 ();
 b15zdnd11an1n08x5 FILLER_42_1089 ();
 b15zdnd00an1n02x5 FILLER_42_1097 ();
 b15zdnd11an1n64x5 FILLER_42_1141 ();
 b15zdnd11an1n64x5 FILLER_42_1205 ();
 b15zdnd11an1n64x5 FILLER_42_1269 ();
 b15zdnd11an1n64x5 FILLER_42_1333 ();
 b15zdnd11an1n64x5 FILLER_42_1397 ();
 b15zdnd11an1n16x5 FILLER_42_1461 ();
 b15zdnd00an1n01x5 FILLER_42_1477 ();
 b15zdnd11an1n08x5 FILLER_42_2265 ();
 b15zdnd00an1n02x5 FILLER_42_2273 ();
 b15zdnd00an1n01x5 FILLER_42_2275 ();
 b15zdnd11an1n64x5 FILLER_43_0 ();
 b15zdnd11an1n64x5 FILLER_43_64 ();
 b15zdnd11an1n64x5 FILLER_43_128 ();
 b15zdnd11an1n64x5 FILLER_43_192 ();
 b15zdnd11an1n64x5 FILLER_43_256 ();
 b15zdnd11an1n64x5 FILLER_43_320 ();
 b15zdnd11an1n64x5 FILLER_43_384 ();
 b15zdnd11an1n64x5 FILLER_43_448 ();
 b15zdnd11an1n64x5 FILLER_43_512 ();
 b15zdnd11an1n64x5 FILLER_43_576 ();
 b15zdnd11an1n64x5 FILLER_43_640 ();
 b15zdnd11an1n64x5 FILLER_43_704 ();
 b15zdnd11an1n64x5 FILLER_43_768 ();
 b15zdnd11an1n64x5 FILLER_43_832 ();
 b15zdnd11an1n64x5 FILLER_43_896 ();
 b15zdnd11an1n64x5 FILLER_43_960 ();
 b15zdnd11an1n64x5 FILLER_43_1024 ();
 b15zdnd11an1n16x5 FILLER_43_1088 ();
 b15zdnd11an1n04x5 FILLER_43_1104 ();
 b15zdnd00an1n01x5 FILLER_43_1108 ();
 b15zdnd11an1n32x5 FILLER_43_1151 ();
 b15zdnd00an1n02x5 FILLER_43_1183 ();
 b15zdnd11an1n64x5 FILLER_43_1199 ();
 b15zdnd11an1n64x5 FILLER_43_1263 ();
 b15zdnd11an1n64x5 FILLER_43_1327 ();
 b15zdnd11an1n64x5 FILLER_43_1391 ();
 b15zdnd11an1n16x5 FILLER_43_1455 ();
 b15zdnd11an1n08x5 FILLER_43_1471 ();
 b15zdnd11an1n04x5 FILLER_43_1479 ();
 b15zdnd00an1n02x5 FILLER_43_1483 ();
 b15zdnd00an1n01x5 FILLER_43_1485 ();
 b15zdnd11an1n16x5 FILLER_43_2257 ();
 b15zdnd11an1n08x5 FILLER_43_2273 ();
 b15zdnd00an1n02x5 FILLER_43_2281 ();
 b15zdnd00an1n01x5 FILLER_43_2283 ();
 b15zdnd11an1n64x5 FILLER_44_8 ();
 b15zdnd11an1n64x5 FILLER_44_72 ();
 b15zdnd11an1n64x5 FILLER_44_136 ();
 b15zdnd11an1n64x5 FILLER_44_200 ();
 b15zdnd11an1n64x5 FILLER_44_264 ();
 b15zdnd11an1n64x5 FILLER_44_328 ();
 b15zdnd11an1n64x5 FILLER_44_392 ();
 b15zdnd11an1n64x5 FILLER_44_456 ();
 b15zdnd11an1n64x5 FILLER_44_520 ();
 b15zdnd11an1n64x5 FILLER_44_584 ();
 b15zdnd11an1n64x5 FILLER_44_648 ();
 b15zdnd11an1n04x5 FILLER_44_712 ();
 b15zdnd00an1n02x5 FILLER_44_716 ();
 b15zdnd11an1n64x5 FILLER_44_726 ();
 b15zdnd11an1n64x5 FILLER_44_790 ();
 b15zdnd11an1n64x5 FILLER_44_854 ();
 b15zdnd11an1n64x5 FILLER_44_918 ();
 b15zdnd11an1n64x5 FILLER_44_982 ();
 b15zdnd11an1n32x5 FILLER_44_1046 ();
 b15zdnd11an1n04x5 FILLER_44_1078 ();
 b15zdnd11an1n08x5 FILLER_44_1124 ();
 b15zdnd11an1n04x5 FILLER_44_1132 ();
 b15zdnd00an1n02x5 FILLER_44_1136 ();
 b15zdnd11an1n64x5 FILLER_44_1180 ();
 b15zdnd11an1n64x5 FILLER_44_1244 ();
 b15zdnd11an1n64x5 FILLER_44_1308 ();
 b15zdnd11an1n64x5 FILLER_44_1372 ();
 b15zdnd11an1n32x5 FILLER_44_1436 ();
 b15zdnd11an1n08x5 FILLER_44_1468 ();
 b15zdnd00an1n02x5 FILLER_44_1476 ();
 b15zdnd11an1n08x5 FILLER_44_2265 ();
 b15zdnd00an1n02x5 FILLER_44_2273 ();
 b15zdnd00an1n01x5 FILLER_44_2275 ();
 b15zdnd11an1n64x5 FILLER_45_0 ();
 b15zdnd11an1n64x5 FILLER_45_64 ();
 b15zdnd11an1n64x5 FILLER_45_128 ();
 b15zdnd11an1n64x5 FILLER_45_192 ();
 b15zdnd11an1n64x5 FILLER_45_256 ();
 b15zdnd11an1n64x5 FILLER_45_320 ();
 b15zdnd11an1n64x5 FILLER_45_384 ();
 b15zdnd11an1n64x5 FILLER_45_448 ();
 b15zdnd11an1n64x5 FILLER_45_512 ();
 b15zdnd11an1n64x5 FILLER_45_576 ();
 b15zdnd11an1n64x5 FILLER_45_640 ();
 b15zdnd11an1n64x5 FILLER_45_704 ();
 b15zdnd11an1n64x5 FILLER_45_768 ();
 b15zdnd11an1n64x5 FILLER_45_832 ();
 b15zdnd11an1n64x5 FILLER_45_896 ();
 b15zdnd11an1n64x5 FILLER_45_960 ();
 b15zdnd11an1n64x5 FILLER_45_1024 ();
 b15zdnd11an1n64x5 FILLER_45_1088 ();
 b15zdnd11an1n64x5 FILLER_45_1152 ();
 b15zdnd11an1n64x5 FILLER_45_1216 ();
 b15zdnd11an1n64x5 FILLER_45_1280 ();
 b15zdnd11an1n64x5 FILLER_45_1344 ();
 b15zdnd11an1n64x5 FILLER_45_1408 ();
 b15zdnd11an1n08x5 FILLER_45_1472 ();
 b15zdnd11an1n04x5 FILLER_45_1480 ();
 b15zdnd00an1n02x5 FILLER_45_1484 ();
 b15zdnd11an1n16x5 FILLER_45_2257 ();
 b15zdnd11an1n08x5 FILLER_45_2273 ();
 b15zdnd00an1n02x5 FILLER_45_2281 ();
 b15zdnd00an1n01x5 FILLER_45_2283 ();
 b15zdnd11an1n64x5 FILLER_46_8 ();
 b15zdnd11an1n64x5 FILLER_46_72 ();
 b15zdnd11an1n64x5 FILLER_46_136 ();
 b15zdnd11an1n64x5 FILLER_46_200 ();
 b15zdnd11an1n64x5 FILLER_46_264 ();
 b15zdnd11an1n32x5 FILLER_46_328 ();
 b15zdnd11an1n08x5 FILLER_46_360 ();
 b15zdnd11an1n04x5 FILLER_46_368 ();
 b15zdnd00an1n02x5 FILLER_46_372 ();
 b15zdnd00an1n01x5 FILLER_46_374 ();
 b15zdnd11an1n32x5 FILLER_46_391 ();
 b15zdnd11an1n04x5 FILLER_46_423 ();
 b15zdnd00an1n02x5 FILLER_46_427 ();
 b15zdnd00an1n01x5 FILLER_46_429 ();
 b15zdnd11an1n64x5 FILLER_46_461 ();
 b15zdnd11an1n64x5 FILLER_46_525 ();
 b15zdnd11an1n64x5 FILLER_46_589 ();
 b15zdnd11an1n64x5 FILLER_46_653 ();
 b15zdnd00an1n01x5 FILLER_46_717 ();
 b15zdnd00an1n02x5 FILLER_46_726 ();
 b15zdnd11an1n32x5 FILLER_46_739 ();
 b15zdnd11an1n08x5 FILLER_46_771 ();
 b15zdnd11an1n64x5 FILLER_46_790 ();
 b15zdnd11an1n64x5 FILLER_46_854 ();
 b15zdnd11an1n64x5 FILLER_46_918 ();
 b15zdnd11an1n64x5 FILLER_46_982 ();
 b15zdnd11an1n64x5 FILLER_46_1046 ();
 b15zdnd11an1n64x5 FILLER_46_1110 ();
 b15zdnd11an1n64x5 FILLER_46_1174 ();
 b15zdnd11an1n64x5 FILLER_46_1238 ();
 b15zdnd11an1n64x5 FILLER_46_1302 ();
 b15zdnd11an1n64x5 FILLER_46_1366 ();
 b15zdnd11an1n32x5 FILLER_46_1430 ();
 b15zdnd11an1n16x5 FILLER_46_1462 ();
 b15zdnd11an1n08x5 FILLER_46_2265 ();
 b15zdnd00an1n02x5 FILLER_46_2273 ();
 b15zdnd00an1n01x5 FILLER_46_2275 ();
 b15zdnd11an1n64x5 FILLER_47_0 ();
 b15zdnd11an1n64x5 FILLER_47_64 ();
 b15zdnd11an1n64x5 FILLER_47_128 ();
 b15zdnd11an1n64x5 FILLER_47_192 ();
 b15zdnd11an1n64x5 FILLER_47_256 ();
 b15zdnd11an1n64x5 FILLER_47_320 ();
 b15zdnd11an1n64x5 FILLER_47_384 ();
 b15zdnd11an1n64x5 FILLER_47_448 ();
 b15zdnd11an1n64x5 FILLER_47_512 ();
 b15zdnd11an1n64x5 FILLER_47_576 ();
 b15zdnd11an1n32x5 FILLER_47_640 ();
 b15zdnd11an1n16x5 FILLER_47_672 ();
 b15zdnd11an1n64x5 FILLER_47_730 ();
 b15zdnd11an1n64x5 FILLER_47_794 ();
 b15zdnd11an1n64x5 FILLER_47_858 ();
 b15zdnd11an1n64x5 FILLER_47_922 ();
 b15zdnd11an1n64x5 FILLER_47_986 ();
 b15zdnd11an1n64x5 FILLER_47_1050 ();
 b15zdnd11an1n64x5 FILLER_47_1114 ();
 b15zdnd11an1n64x5 FILLER_47_1178 ();
 b15zdnd11an1n64x5 FILLER_47_1242 ();
 b15zdnd11an1n64x5 FILLER_47_1306 ();
 b15zdnd11an1n64x5 FILLER_47_1370 ();
 b15zdnd11an1n32x5 FILLER_47_1434 ();
 b15zdnd11an1n16x5 FILLER_47_1466 ();
 b15zdnd11an1n04x5 FILLER_47_1482 ();
 b15zdnd11an1n16x5 FILLER_47_2257 ();
 b15zdnd11an1n08x5 FILLER_47_2273 ();
 b15zdnd00an1n02x5 FILLER_47_2281 ();
 b15zdnd00an1n01x5 FILLER_47_2283 ();
 b15zdnd11an1n64x5 FILLER_48_8 ();
 b15zdnd11an1n64x5 FILLER_48_72 ();
 b15zdnd11an1n64x5 FILLER_48_136 ();
 b15zdnd11an1n64x5 FILLER_48_200 ();
 b15zdnd11an1n64x5 FILLER_48_264 ();
 b15zdnd11an1n64x5 FILLER_48_328 ();
 b15zdnd11an1n64x5 FILLER_48_392 ();
 b15zdnd11an1n64x5 FILLER_48_456 ();
 b15zdnd11an1n64x5 FILLER_48_520 ();
 b15zdnd11an1n64x5 FILLER_48_584 ();
 b15zdnd11an1n64x5 FILLER_48_648 ();
 b15zdnd11an1n04x5 FILLER_48_712 ();
 b15zdnd00an1n02x5 FILLER_48_716 ();
 b15zdnd11an1n64x5 FILLER_48_726 ();
 b15zdnd11an1n64x5 FILLER_48_790 ();
 b15zdnd11an1n64x5 FILLER_48_854 ();
 b15zdnd11an1n64x5 FILLER_48_918 ();
 b15zdnd11an1n64x5 FILLER_48_982 ();
 b15zdnd11an1n64x5 FILLER_48_1046 ();
 b15zdnd11an1n64x5 FILLER_48_1110 ();
 b15zdnd11an1n64x5 FILLER_48_1174 ();
 b15zdnd11an1n64x5 FILLER_48_1238 ();
 b15zdnd11an1n64x5 FILLER_48_1302 ();
 b15zdnd11an1n64x5 FILLER_48_1366 ();
 b15zdnd11an1n32x5 FILLER_48_1430 ();
 b15zdnd11an1n16x5 FILLER_48_1462 ();
 b15zdnd11an1n08x5 FILLER_48_2265 ();
 b15zdnd00an1n02x5 FILLER_48_2273 ();
 b15zdnd00an1n01x5 FILLER_48_2275 ();
 b15zdnd11an1n64x5 FILLER_49_0 ();
 b15zdnd11an1n64x5 FILLER_49_64 ();
 b15zdnd11an1n64x5 FILLER_49_128 ();
 b15zdnd11an1n64x5 FILLER_49_192 ();
 b15zdnd11an1n64x5 FILLER_49_256 ();
 b15zdnd11an1n64x5 FILLER_49_320 ();
 b15zdnd11an1n64x5 FILLER_49_384 ();
 b15zdnd11an1n64x5 FILLER_49_448 ();
 b15zdnd11an1n64x5 FILLER_49_512 ();
 b15zdnd11an1n64x5 FILLER_49_576 ();
 b15zdnd11an1n64x5 FILLER_49_640 ();
 b15zdnd11an1n64x5 FILLER_49_704 ();
 b15zdnd11an1n64x5 FILLER_49_768 ();
 b15zdnd11an1n64x5 FILLER_49_832 ();
 b15zdnd11an1n64x5 FILLER_49_896 ();
 b15zdnd11an1n64x5 FILLER_49_960 ();
 b15zdnd11an1n64x5 FILLER_49_1024 ();
 b15zdnd11an1n64x5 FILLER_49_1088 ();
 b15zdnd11an1n64x5 FILLER_49_1152 ();
 b15zdnd11an1n64x5 FILLER_49_1216 ();
 b15zdnd11an1n64x5 FILLER_49_1280 ();
 b15zdnd11an1n64x5 FILLER_49_1344 ();
 b15zdnd11an1n64x5 FILLER_49_1408 ();
 b15zdnd11an1n08x5 FILLER_49_1472 ();
 b15zdnd11an1n04x5 FILLER_49_1480 ();
 b15zdnd00an1n02x5 FILLER_49_1484 ();
 b15zdnd11an1n16x5 FILLER_49_2257 ();
 b15zdnd11an1n08x5 FILLER_49_2273 ();
 b15zdnd00an1n02x5 FILLER_49_2281 ();
 b15zdnd00an1n01x5 FILLER_49_2283 ();
 b15zdnd11an1n64x5 FILLER_50_8 ();
 b15zdnd11an1n64x5 FILLER_50_72 ();
 b15zdnd11an1n64x5 FILLER_50_136 ();
 b15zdnd11an1n64x5 FILLER_50_200 ();
 b15zdnd11an1n64x5 FILLER_50_264 ();
 b15zdnd11an1n64x5 FILLER_50_328 ();
 b15zdnd11an1n08x5 FILLER_50_392 ();
 b15zdnd00an1n02x5 FILLER_50_400 ();
 b15zdnd11an1n64x5 FILLER_50_414 ();
 b15zdnd11an1n64x5 FILLER_50_478 ();
 b15zdnd11an1n16x5 FILLER_50_542 ();
 b15zdnd00an1n01x5 FILLER_50_558 ();
 b15zdnd11an1n64x5 FILLER_50_601 ();
 b15zdnd11an1n32x5 FILLER_50_665 ();
 b15zdnd11an1n16x5 FILLER_50_697 ();
 b15zdnd11an1n04x5 FILLER_50_713 ();
 b15zdnd00an1n01x5 FILLER_50_717 ();
 b15zdnd11an1n64x5 FILLER_50_726 ();
 b15zdnd11an1n64x5 FILLER_50_790 ();
 b15zdnd11an1n64x5 FILLER_50_854 ();
 b15zdnd11an1n64x5 FILLER_50_918 ();
 b15zdnd11an1n64x5 FILLER_50_982 ();
 b15zdnd11an1n64x5 FILLER_50_1046 ();
 b15zdnd11an1n64x5 FILLER_50_1110 ();
 b15zdnd11an1n64x5 FILLER_50_1174 ();
 b15zdnd11an1n64x5 FILLER_50_1238 ();
 b15zdnd11an1n64x5 FILLER_50_1302 ();
 b15zdnd11an1n16x5 FILLER_50_1366 ();
 b15zdnd11an1n04x5 FILLER_50_1382 ();
 b15zdnd00an1n02x5 FILLER_50_1386 ();
 b15zdnd00an1n01x5 FILLER_50_1388 ();
 b15zdnd11an1n64x5 FILLER_50_1400 ();
 b15zdnd11an1n08x5 FILLER_50_1464 ();
 b15zdnd11an1n04x5 FILLER_50_1472 ();
 b15zdnd00an1n02x5 FILLER_50_1476 ();
 b15zdnd11an1n08x5 FILLER_50_2265 ();
 b15zdnd00an1n02x5 FILLER_50_2273 ();
 b15zdnd00an1n01x5 FILLER_50_2275 ();
 b15zdnd11an1n64x5 FILLER_51_0 ();
 b15zdnd11an1n64x5 FILLER_51_64 ();
 b15zdnd11an1n64x5 FILLER_51_128 ();
 b15zdnd11an1n64x5 FILLER_51_192 ();
 b15zdnd11an1n64x5 FILLER_51_256 ();
 b15zdnd11an1n64x5 FILLER_51_320 ();
 b15zdnd11an1n64x5 FILLER_51_384 ();
 b15zdnd11an1n64x5 FILLER_51_448 ();
 b15zdnd11an1n64x5 FILLER_51_512 ();
 b15zdnd11an1n64x5 FILLER_51_576 ();
 b15zdnd00an1n02x5 FILLER_51_640 ();
 b15zdnd11an1n04x5 FILLER_51_645 ();
 b15zdnd11an1n08x5 FILLER_51_652 ();
 b15zdnd11an1n64x5 FILLER_51_663 ();
 b15zdnd11an1n64x5 FILLER_51_727 ();
 b15zdnd11an1n64x5 FILLER_51_791 ();
 b15zdnd11an1n64x5 FILLER_51_855 ();
 b15zdnd11an1n64x5 FILLER_51_919 ();
 b15zdnd11an1n64x5 FILLER_51_983 ();
 b15zdnd11an1n64x5 FILLER_51_1047 ();
 b15zdnd11an1n64x5 FILLER_51_1111 ();
 b15zdnd11an1n64x5 FILLER_51_1175 ();
 b15zdnd11an1n64x5 FILLER_51_1239 ();
 b15zdnd11an1n64x5 FILLER_51_1303 ();
 b15zdnd11an1n64x5 FILLER_51_1367 ();
 b15zdnd11an1n32x5 FILLER_51_1431 ();
 b15zdnd11an1n16x5 FILLER_51_1463 ();
 b15zdnd11an1n04x5 FILLER_51_1479 ();
 b15zdnd00an1n02x5 FILLER_51_1483 ();
 b15zdnd00an1n01x5 FILLER_51_1485 ();
 b15zdnd11an1n16x5 FILLER_51_2257 ();
 b15zdnd11an1n08x5 FILLER_51_2273 ();
 b15zdnd00an1n02x5 FILLER_51_2281 ();
 b15zdnd00an1n01x5 FILLER_51_2283 ();
 b15zdnd11an1n64x5 FILLER_52_8 ();
 b15zdnd11an1n64x5 FILLER_52_72 ();
 b15zdnd11an1n64x5 FILLER_52_136 ();
 b15zdnd11an1n64x5 FILLER_52_200 ();
 b15zdnd11an1n64x5 FILLER_52_264 ();
 b15zdnd11an1n64x5 FILLER_52_328 ();
 b15zdnd11an1n64x5 FILLER_52_392 ();
 b15zdnd11an1n64x5 FILLER_52_456 ();
 b15zdnd11an1n64x5 FILLER_52_520 ();
 b15zdnd11an1n32x5 FILLER_52_584 ();
 b15zdnd00an1n01x5 FILLER_52_616 ();
 b15zdnd11an1n32x5 FILLER_52_661 ();
 b15zdnd11an1n16x5 FILLER_52_693 ();
 b15zdnd11an1n08x5 FILLER_52_709 ();
 b15zdnd00an1n01x5 FILLER_52_717 ();
 b15zdnd11an1n32x5 FILLER_52_726 ();
 b15zdnd11an1n16x5 FILLER_52_758 ();
 b15zdnd11an1n04x5 FILLER_52_774 ();
 b15zdnd00an1n01x5 FILLER_52_778 ();
 b15zdnd11an1n64x5 FILLER_52_821 ();
 b15zdnd11an1n16x5 FILLER_52_885 ();
 b15zdnd00an1n01x5 FILLER_52_901 ();
 b15zdnd11an1n64x5 FILLER_52_905 ();
 b15zdnd11an1n64x5 FILLER_52_969 ();
 b15zdnd11an1n64x5 FILLER_52_1033 ();
 b15zdnd11an1n64x5 FILLER_52_1097 ();
 b15zdnd11an1n64x5 FILLER_52_1161 ();
 b15zdnd11an1n64x5 FILLER_52_1225 ();
 b15zdnd11an1n64x5 FILLER_52_1289 ();
 b15zdnd11an1n64x5 FILLER_52_1353 ();
 b15zdnd11an1n32x5 FILLER_52_1417 ();
 b15zdnd11an1n16x5 FILLER_52_1449 ();
 b15zdnd11an1n08x5 FILLER_52_1465 ();
 b15zdnd11an1n04x5 FILLER_52_1473 ();
 b15zdnd00an1n01x5 FILLER_52_1477 ();
 b15zdnd11an1n08x5 FILLER_52_2265 ();
 b15zdnd00an1n02x5 FILLER_52_2273 ();
 b15zdnd00an1n01x5 FILLER_52_2275 ();
 b15zdnd11an1n64x5 FILLER_53_0 ();
 b15zdnd11an1n64x5 FILLER_53_64 ();
 b15zdnd11an1n64x5 FILLER_53_128 ();
 b15zdnd11an1n64x5 FILLER_53_192 ();
 b15zdnd11an1n64x5 FILLER_53_256 ();
 b15zdnd11an1n64x5 FILLER_53_320 ();
 b15zdnd11an1n16x5 FILLER_53_384 ();
 b15zdnd00an1n02x5 FILLER_53_400 ();
 b15zdnd00an1n01x5 FILLER_53_402 ();
 b15zdnd11an1n32x5 FILLER_53_414 ();
 b15zdnd00an1n02x5 FILLER_53_446 ();
 b15zdnd11an1n32x5 FILLER_53_493 ();
 b15zdnd11an1n16x5 FILLER_53_525 ();
 b15zdnd11an1n04x5 FILLER_53_541 ();
 b15zdnd00an1n02x5 FILLER_53_545 ();
 b15zdnd00an1n01x5 FILLER_53_547 ();
 b15zdnd11an1n64x5 FILLER_53_590 ();
 b15zdnd11an1n32x5 FILLER_53_654 ();
 b15zdnd11an1n16x5 FILLER_53_686 ();
 b15zdnd11an1n08x5 FILLER_53_702 ();
 b15zdnd11an1n32x5 FILLER_53_754 ();
 b15zdnd11an1n16x5 FILLER_53_786 ();
 b15zdnd11an1n04x5 FILLER_53_802 ();
 b15zdnd00an1n01x5 FILLER_53_806 ();
 b15zdnd11an1n32x5 FILLER_53_849 ();
 b15zdnd11an1n16x5 FILLER_53_881 ();
 b15zdnd11an1n04x5 FILLER_53_897 ();
 b15zdnd11an1n64x5 FILLER_53_904 ();
 b15zdnd11an1n64x5 FILLER_53_968 ();
 b15zdnd11an1n64x5 FILLER_53_1032 ();
 b15zdnd11an1n64x5 FILLER_53_1096 ();
 b15zdnd11an1n64x5 FILLER_53_1160 ();
 b15zdnd11an1n32x5 FILLER_53_1224 ();
 b15zdnd11an1n16x5 FILLER_53_1256 ();
 b15zdnd11an1n04x5 FILLER_53_1272 ();
 b15zdnd00an1n02x5 FILLER_53_1276 ();
 b15zdnd00an1n01x5 FILLER_53_1278 ();
 b15zdnd11an1n64x5 FILLER_53_1293 ();
 b15zdnd11an1n64x5 FILLER_53_1357 ();
 b15zdnd11an1n64x5 FILLER_53_1421 ();
 b15zdnd00an1n01x5 FILLER_53_1485 ();
 b15zdnd11an1n16x5 FILLER_53_2257 ();
 b15zdnd11an1n08x5 FILLER_53_2273 ();
 b15zdnd00an1n02x5 FILLER_53_2281 ();
 b15zdnd00an1n01x5 FILLER_53_2283 ();
 b15zdnd11an1n64x5 FILLER_54_8 ();
 b15zdnd11an1n64x5 FILLER_54_72 ();
 b15zdnd11an1n64x5 FILLER_54_136 ();
 b15zdnd11an1n64x5 FILLER_54_200 ();
 b15zdnd11an1n64x5 FILLER_54_264 ();
 b15zdnd11an1n64x5 FILLER_54_328 ();
 b15zdnd11an1n64x5 FILLER_54_392 ();
 b15zdnd11an1n64x5 FILLER_54_456 ();
 b15zdnd11an1n64x5 FILLER_54_520 ();
 b15zdnd11an1n64x5 FILLER_54_584 ();
 b15zdnd11an1n64x5 FILLER_54_648 ();
 b15zdnd11an1n04x5 FILLER_54_712 ();
 b15zdnd00an1n02x5 FILLER_54_716 ();
 b15zdnd11an1n04x5 FILLER_54_726 ();
 b15zdnd00an1n02x5 FILLER_54_730 ();
 b15zdnd11an1n04x5 FILLER_54_735 ();
 b15zdnd11an1n04x5 FILLER_54_742 ();
 b15zdnd11an1n64x5 FILLER_54_749 ();
 b15zdnd11an1n64x5 FILLER_54_813 ();
 b15zdnd00an1n02x5 FILLER_54_877 ();
 b15zdnd00an1n01x5 FILLER_54_879 ();
 b15zdnd11an1n64x5 FILLER_54_924 ();
 b15zdnd11an1n64x5 FILLER_54_988 ();
 b15zdnd11an1n64x5 FILLER_54_1052 ();
 b15zdnd11an1n64x5 FILLER_54_1116 ();
 b15zdnd11an1n64x5 FILLER_54_1180 ();
 b15zdnd11an1n64x5 FILLER_54_1244 ();
 b15zdnd11an1n64x5 FILLER_54_1308 ();
 b15zdnd11an1n64x5 FILLER_54_1372 ();
 b15zdnd11an1n32x5 FILLER_54_1436 ();
 b15zdnd11an1n08x5 FILLER_54_1468 ();
 b15zdnd00an1n02x5 FILLER_54_1476 ();
 b15zdnd11an1n08x5 FILLER_54_2265 ();
 b15zdnd00an1n02x5 FILLER_54_2273 ();
 b15zdnd00an1n01x5 FILLER_54_2275 ();
 b15zdnd11an1n64x5 FILLER_55_0 ();
 b15zdnd11an1n64x5 FILLER_55_64 ();
 b15zdnd11an1n64x5 FILLER_55_128 ();
 b15zdnd11an1n64x5 FILLER_55_192 ();
 b15zdnd11an1n64x5 FILLER_55_256 ();
 b15zdnd11an1n64x5 FILLER_55_320 ();
 b15zdnd11an1n64x5 FILLER_55_384 ();
 b15zdnd11an1n64x5 FILLER_55_448 ();
 b15zdnd11an1n64x5 FILLER_55_512 ();
 b15zdnd11an1n64x5 FILLER_55_576 ();
 b15zdnd11an1n64x5 FILLER_55_640 ();
 b15zdnd00an1n02x5 FILLER_55_704 ();
 b15zdnd11an1n64x5 FILLER_55_748 ();
 b15zdnd11an1n64x5 FILLER_55_812 ();
 b15zdnd11an1n16x5 FILLER_55_876 ();
 b15zdnd11an1n04x5 FILLER_55_892 ();
 b15zdnd00an1n02x5 FILLER_55_896 ();
 b15zdnd00an1n01x5 FILLER_55_898 ();
 b15zdnd11an1n64x5 FILLER_55_902 ();
 b15zdnd11an1n64x5 FILLER_55_966 ();
 b15zdnd11an1n64x5 FILLER_55_1030 ();
 b15zdnd11an1n64x5 FILLER_55_1094 ();
 b15zdnd11an1n64x5 FILLER_55_1158 ();
 b15zdnd11an1n64x5 FILLER_55_1222 ();
 b15zdnd11an1n64x5 FILLER_55_1286 ();
 b15zdnd11an1n64x5 FILLER_55_1350 ();
 b15zdnd11an1n64x5 FILLER_55_1414 ();
 b15zdnd11an1n08x5 FILLER_55_1478 ();
 b15zdnd11an1n16x5 FILLER_55_2257 ();
 b15zdnd11an1n08x5 FILLER_55_2273 ();
 b15zdnd00an1n02x5 FILLER_55_2281 ();
 b15zdnd00an1n01x5 FILLER_55_2283 ();
 b15zdnd11an1n64x5 FILLER_56_8 ();
 b15zdnd11an1n64x5 FILLER_56_72 ();
 b15zdnd11an1n64x5 FILLER_56_136 ();
 b15zdnd11an1n64x5 FILLER_56_200 ();
 b15zdnd11an1n64x5 FILLER_56_264 ();
 b15zdnd11an1n32x5 FILLER_56_328 ();
 b15zdnd11an1n16x5 FILLER_56_360 ();
 b15zdnd11an1n08x5 FILLER_56_376 ();
 b15zdnd11an1n04x5 FILLER_56_384 ();
 b15zdnd11an1n64x5 FILLER_56_402 ();
 b15zdnd11an1n64x5 FILLER_56_466 ();
 b15zdnd11an1n64x5 FILLER_56_530 ();
 b15zdnd11an1n64x5 FILLER_56_594 ();
 b15zdnd11an1n32x5 FILLER_56_658 ();
 b15zdnd11an1n16x5 FILLER_56_690 ();
 b15zdnd11an1n08x5 FILLER_56_706 ();
 b15zdnd11an1n04x5 FILLER_56_714 ();
 b15zdnd11an1n64x5 FILLER_56_726 ();
 b15zdnd11an1n64x5 FILLER_56_790 ();
 b15zdnd11an1n64x5 FILLER_56_854 ();
 b15zdnd11an1n64x5 FILLER_56_918 ();
 b15zdnd11an1n32x5 FILLER_56_982 ();
 b15zdnd11an1n08x5 FILLER_56_1014 ();
 b15zdnd11an1n64x5 FILLER_56_1064 ();
 b15zdnd11an1n64x5 FILLER_56_1128 ();
 b15zdnd11an1n64x5 FILLER_56_1192 ();
 b15zdnd11an1n64x5 FILLER_56_1256 ();
 b15zdnd11an1n64x5 FILLER_56_1320 ();
 b15zdnd11an1n64x5 FILLER_56_1384 ();
 b15zdnd11an1n16x5 FILLER_56_1448 ();
 b15zdnd11an1n08x5 FILLER_56_1464 ();
 b15zdnd11an1n04x5 FILLER_56_1472 ();
 b15zdnd00an1n02x5 FILLER_56_1476 ();
 b15zdnd11an1n08x5 FILLER_56_2265 ();
 b15zdnd00an1n02x5 FILLER_56_2273 ();
 b15zdnd00an1n01x5 FILLER_56_2275 ();
 b15zdnd11an1n64x5 FILLER_57_0 ();
 b15zdnd11an1n64x5 FILLER_57_64 ();
 b15zdnd11an1n64x5 FILLER_57_128 ();
 b15zdnd11an1n64x5 FILLER_57_192 ();
 b15zdnd11an1n64x5 FILLER_57_256 ();
 b15zdnd11an1n64x5 FILLER_57_320 ();
 b15zdnd11an1n64x5 FILLER_57_384 ();
 b15zdnd11an1n64x5 FILLER_57_448 ();
 b15zdnd11an1n08x5 FILLER_57_512 ();
 b15zdnd11an1n04x5 FILLER_57_520 ();
 b15zdnd11an1n64x5 FILLER_57_566 ();
 b15zdnd11an1n08x5 FILLER_57_630 ();
 b15zdnd11an1n64x5 FILLER_57_680 ();
 b15zdnd11an1n64x5 FILLER_57_744 ();
 b15zdnd11an1n64x5 FILLER_57_808 ();
 b15zdnd11an1n64x5 FILLER_57_872 ();
 b15zdnd11an1n64x5 FILLER_57_936 ();
 b15zdnd11an1n64x5 FILLER_57_1000 ();
 b15zdnd11an1n64x5 FILLER_57_1064 ();
 b15zdnd11an1n64x5 FILLER_57_1128 ();
 b15zdnd11an1n64x5 FILLER_57_1192 ();
 b15zdnd11an1n64x5 FILLER_57_1256 ();
 b15zdnd11an1n64x5 FILLER_57_1320 ();
 b15zdnd11an1n64x5 FILLER_57_1384 ();
 b15zdnd11an1n32x5 FILLER_57_1448 ();
 b15zdnd11an1n04x5 FILLER_57_1480 ();
 b15zdnd00an1n02x5 FILLER_57_1484 ();
 b15zdnd11an1n16x5 FILLER_57_2257 ();
 b15zdnd11an1n08x5 FILLER_57_2273 ();
 b15zdnd00an1n02x5 FILLER_57_2281 ();
 b15zdnd00an1n01x5 FILLER_57_2283 ();
 b15zdnd11an1n64x5 FILLER_58_8 ();
 b15zdnd11an1n64x5 FILLER_58_72 ();
 b15zdnd11an1n64x5 FILLER_58_136 ();
 b15zdnd11an1n64x5 FILLER_58_200 ();
 b15zdnd11an1n64x5 FILLER_58_264 ();
 b15zdnd11an1n64x5 FILLER_58_328 ();
 b15zdnd11an1n64x5 FILLER_58_409 ();
 b15zdnd11an1n64x5 FILLER_58_473 ();
 b15zdnd11an1n64x5 FILLER_58_537 ();
 b15zdnd11an1n64x5 FILLER_58_601 ();
 b15zdnd11an1n32x5 FILLER_58_665 ();
 b15zdnd11an1n16x5 FILLER_58_697 ();
 b15zdnd11an1n04x5 FILLER_58_713 ();
 b15zdnd00an1n01x5 FILLER_58_717 ();
 b15zdnd11an1n64x5 FILLER_58_726 ();
 b15zdnd11an1n64x5 FILLER_58_790 ();
 b15zdnd11an1n32x5 FILLER_58_854 ();
 b15zdnd11an1n04x5 FILLER_58_886 ();
 b15zdnd11an1n64x5 FILLER_58_932 ();
 b15zdnd11an1n64x5 FILLER_58_996 ();
 b15zdnd11an1n64x5 FILLER_58_1060 ();
 b15zdnd11an1n64x5 FILLER_58_1124 ();
 b15zdnd11an1n64x5 FILLER_58_1188 ();
 b15zdnd11an1n64x5 FILLER_58_1252 ();
 b15zdnd11an1n64x5 FILLER_58_1316 ();
 b15zdnd11an1n64x5 FILLER_58_1380 ();
 b15zdnd11an1n32x5 FILLER_58_1444 ();
 b15zdnd00an1n02x5 FILLER_58_1476 ();
 b15zdnd11an1n08x5 FILLER_58_2265 ();
 b15zdnd00an1n02x5 FILLER_58_2273 ();
 b15zdnd00an1n01x5 FILLER_58_2275 ();
 b15zdnd11an1n64x5 FILLER_59_0 ();
 b15zdnd11an1n64x5 FILLER_59_64 ();
 b15zdnd11an1n64x5 FILLER_59_128 ();
 b15zdnd11an1n64x5 FILLER_59_192 ();
 b15zdnd11an1n64x5 FILLER_59_256 ();
 b15zdnd11an1n64x5 FILLER_59_320 ();
 b15zdnd11an1n64x5 FILLER_59_384 ();
 b15zdnd11an1n64x5 FILLER_59_448 ();
 b15zdnd11an1n64x5 FILLER_59_512 ();
 b15zdnd11an1n32x5 FILLER_59_576 ();
 b15zdnd11an1n08x5 FILLER_59_608 ();
 b15zdnd00an1n02x5 FILLER_59_616 ();
 b15zdnd11an1n64x5 FILLER_59_660 ();
 b15zdnd11an1n64x5 FILLER_59_724 ();
 b15zdnd11an1n64x5 FILLER_59_788 ();
 b15zdnd11an1n64x5 FILLER_59_852 ();
 b15zdnd11an1n64x5 FILLER_59_916 ();
 b15zdnd11an1n64x5 FILLER_59_980 ();
 b15zdnd11an1n64x5 FILLER_59_1044 ();
 b15zdnd11an1n64x5 FILLER_59_1108 ();
 b15zdnd11an1n64x5 FILLER_59_1172 ();
 b15zdnd11an1n64x5 FILLER_59_1236 ();
 b15zdnd11an1n64x5 FILLER_59_1300 ();
 b15zdnd11an1n64x5 FILLER_59_1364 ();
 b15zdnd11an1n32x5 FILLER_59_1428 ();
 b15zdnd11an1n16x5 FILLER_59_1460 ();
 b15zdnd11an1n08x5 FILLER_59_1476 ();
 b15zdnd00an1n02x5 FILLER_59_1484 ();
 b15zdnd11an1n16x5 FILLER_59_2257 ();
 b15zdnd11an1n08x5 FILLER_59_2273 ();
 b15zdnd00an1n02x5 FILLER_59_2281 ();
 b15zdnd00an1n01x5 FILLER_59_2283 ();
 b15zdnd11an1n64x5 FILLER_60_8 ();
 b15zdnd11an1n64x5 FILLER_60_72 ();
 b15zdnd11an1n64x5 FILLER_60_136 ();
 b15zdnd11an1n64x5 FILLER_60_200 ();
 b15zdnd11an1n64x5 FILLER_60_264 ();
 b15zdnd11an1n64x5 FILLER_60_328 ();
 b15zdnd11an1n08x5 FILLER_60_392 ();
 b15zdnd11an1n04x5 FILLER_60_400 ();
 b15zdnd00an1n01x5 FILLER_60_404 ();
 b15zdnd11an1n32x5 FILLER_60_413 ();
 b15zdnd11an1n04x5 FILLER_60_445 ();
 b15zdnd00an1n02x5 FILLER_60_449 ();
 b15zdnd00an1n01x5 FILLER_60_451 ();
 b15zdnd11an1n64x5 FILLER_60_497 ();
 b15zdnd11an1n64x5 FILLER_60_561 ();
 b15zdnd11an1n64x5 FILLER_60_625 ();
 b15zdnd11an1n16x5 FILLER_60_689 ();
 b15zdnd11an1n08x5 FILLER_60_705 ();
 b15zdnd11an1n04x5 FILLER_60_713 ();
 b15zdnd00an1n01x5 FILLER_60_717 ();
 b15zdnd11an1n64x5 FILLER_60_726 ();
 b15zdnd11an1n64x5 FILLER_60_790 ();
 b15zdnd11an1n64x5 FILLER_60_854 ();
 b15zdnd11an1n64x5 FILLER_60_918 ();
 b15zdnd11an1n64x5 FILLER_60_982 ();
 b15zdnd11an1n64x5 FILLER_60_1046 ();
 b15zdnd11an1n64x5 FILLER_60_1110 ();
 b15zdnd11an1n64x5 FILLER_60_1174 ();
 b15zdnd11an1n64x5 FILLER_60_1238 ();
 b15zdnd11an1n64x5 FILLER_60_1302 ();
 b15zdnd11an1n64x5 FILLER_60_1366 ();
 b15zdnd11an1n32x5 FILLER_60_1430 ();
 b15zdnd11an1n16x5 FILLER_60_1462 ();
 b15zdnd11an1n08x5 FILLER_60_2265 ();
 b15zdnd00an1n02x5 FILLER_60_2273 ();
 b15zdnd00an1n01x5 FILLER_60_2275 ();
 b15zdnd11an1n64x5 FILLER_61_0 ();
 b15zdnd11an1n64x5 FILLER_61_64 ();
 b15zdnd11an1n64x5 FILLER_61_128 ();
 b15zdnd11an1n64x5 FILLER_61_192 ();
 b15zdnd11an1n64x5 FILLER_61_256 ();
 b15zdnd11an1n64x5 FILLER_61_320 ();
 b15zdnd11an1n04x5 FILLER_61_384 ();
 b15zdnd11an1n64x5 FILLER_61_433 ();
 b15zdnd11an1n16x5 FILLER_61_497 ();
 b15zdnd11an1n08x5 FILLER_61_513 ();
 b15zdnd00an1n01x5 FILLER_61_521 ();
 b15zdnd11an1n64x5 FILLER_61_564 ();
 b15zdnd11an1n16x5 FILLER_61_628 ();
 b15zdnd11an1n64x5 FILLER_61_647 ();
 b15zdnd11an1n64x5 FILLER_61_711 ();
 b15zdnd11an1n32x5 FILLER_61_775 ();
 b15zdnd11an1n16x5 FILLER_61_807 ();
 b15zdnd11an1n08x5 FILLER_61_823 ();
 b15zdnd11an1n04x5 FILLER_61_831 ();
 b15zdnd00an1n02x5 FILLER_61_835 ();
 b15zdnd00an1n01x5 FILLER_61_837 ();
 b15zdnd11an1n64x5 FILLER_61_880 ();
 b15zdnd11an1n32x5 FILLER_61_944 ();
 b15zdnd11an1n08x5 FILLER_61_976 ();
 b15zdnd00an1n01x5 FILLER_61_984 ();
 b15zdnd11an1n64x5 FILLER_61_988 ();
 b15zdnd11an1n64x5 FILLER_61_1052 ();
 b15zdnd11an1n64x5 FILLER_61_1116 ();
 b15zdnd11an1n64x5 FILLER_61_1180 ();
 b15zdnd11an1n64x5 FILLER_61_1244 ();
 b15zdnd11an1n64x5 FILLER_61_1308 ();
 b15zdnd11an1n64x5 FILLER_61_1372 ();
 b15zdnd11an1n32x5 FILLER_61_1436 ();
 b15zdnd11an1n16x5 FILLER_61_1468 ();
 b15zdnd00an1n02x5 FILLER_61_1484 ();
 b15zdnd11an1n16x5 FILLER_61_2257 ();
 b15zdnd11an1n08x5 FILLER_61_2273 ();
 b15zdnd00an1n02x5 FILLER_61_2281 ();
 b15zdnd00an1n01x5 FILLER_61_2283 ();
 b15zdnd11an1n64x5 FILLER_62_8 ();
 b15zdnd11an1n64x5 FILLER_62_72 ();
 b15zdnd11an1n64x5 FILLER_62_136 ();
 b15zdnd11an1n64x5 FILLER_62_200 ();
 b15zdnd11an1n64x5 FILLER_62_264 ();
 b15zdnd11an1n64x5 FILLER_62_328 ();
 b15zdnd11an1n64x5 FILLER_62_392 ();
 b15zdnd11an1n64x5 FILLER_62_456 ();
 b15zdnd11an1n64x5 FILLER_62_520 ();
 b15zdnd11an1n32x5 FILLER_62_584 ();
 b15zdnd11an1n16x5 FILLER_62_616 ();
 b15zdnd11an1n04x5 FILLER_62_632 ();
 b15zdnd00an1n02x5 FILLER_62_636 ();
 b15zdnd00an1n01x5 FILLER_62_638 ();
 b15zdnd11an1n04x5 FILLER_62_642 ();
 b15zdnd00an1n01x5 FILLER_62_646 ();
 b15zdnd11an1n64x5 FILLER_62_650 ();
 b15zdnd11an1n04x5 FILLER_62_714 ();
 b15zdnd11an1n64x5 FILLER_62_726 ();
 b15zdnd11an1n64x5 FILLER_62_790 ();
 b15zdnd11an1n64x5 FILLER_62_854 ();
 b15zdnd11an1n32x5 FILLER_62_918 ();
 b15zdnd11an1n08x5 FILLER_62_950 ();
 b15zdnd00an1n02x5 FILLER_62_958 ();
 b15zdnd00an1n01x5 FILLER_62_960 ();
 b15zdnd11an1n64x5 FILLER_62_1005 ();
 b15zdnd11an1n64x5 FILLER_62_1069 ();
 b15zdnd11an1n64x5 FILLER_62_1133 ();
 b15zdnd11an1n64x5 FILLER_62_1197 ();
 b15zdnd11an1n64x5 FILLER_62_1261 ();
 b15zdnd11an1n64x5 FILLER_62_1325 ();
 b15zdnd11an1n64x5 FILLER_62_1389 ();
 b15zdnd11an1n16x5 FILLER_62_1453 ();
 b15zdnd11an1n08x5 FILLER_62_1469 ();
 b15zdnd00an1n01x5 FILLER_62_1477 ();
 b15zdnd11an1n08x5 FILLER_62_2265 ();
 b15zdnd00an1n02x5 FILLER_62_2273 ();
 b15zdnd00an1n01x5 FILLER_62_2275 ();
 b15zdnd11an1n64x5 FILLER_63_0 ();
 b15zdnd11an1n64x5 FILLER_63_64 ();
 b15zdnd11an1n64x5 FILLER_63_128 ();
 b15zdnd11an1n64x5 FILLER_63_192 ();
 b15zdnd11an1n64x5 FILLER_63_256 ();
 b15zdnd11an1n64x5 FILLER_63_320 ();
 b15zdnd11an1n64x5 FILLER_63_384 ();
 b15zdnd11an1n64x5 FILLER_63_448 ();
 b15zdnd11an1n64x5 FILLER_63_512 ();
 b15zdnd11an1n16x5 FILLER_63_576 ();
 b15zdnd11an1n08x5 FILLER_63_592 ();
 b15zdnd11an1n04x5 FILLER_63_600 ();
 b15zdnd00an1n02x5 FILLER_63_604 ();
 b15zdnd11an1n64x5 FILLER_63_650 ();
 b15zdnd11an1n64x5 FILLER_63_714 ();
 b15zdnd11an1n64x5 FILLER_63_778 ();
 b15zdnd11an1n64x5 FILLER_63_842 ();
 b15zdnd11an1n64x5 FILLER_63_906 ();
 b15zdnd11an1n04x5 FILLER_63_970 ();
 b15zdnd00an1n02x5 FILLER_63_974 ();
 b15zdnd00an1n01x5 FILLER_63_976 ();
 b15zdnd11an1n04x5 FILLER_63_980 ();
 b15zdnd11an1n64x5 FILLER_63_987 ();
 b15zdnd11an1n64x5 FILLER_63_1051 ();
 b15zdnd11an1n64x5 FILLER_63_1115 ();
 b15zdnd11an1n64x5 FILLER_63_1179 ();
 b15zdnd11an1n64x5 FILLER_63_1243 ();
 b15zdnd11an1n64x5 FILLER_63_1307 ();
 b15zdnd11an1n64x5 FILLER_63_1371 ();
 b15zdnd11an1n32x5 FILLER_63_1435 ();
 b15zdnd11an1n16x5 FILLER_63_1467 ();
 b15zdnd00an1n02x5 FILLER_63_1483 ();
 b15zdnd00an1n01x5 FILLER_63_1485 ();
 b15zdnd11an1n16x5 FILLER_63_2257 ();
 b15zdnd11an1n08x5 FILLER_63_2273 ();
 b15zdnd00an1n02x5 FILLER_63_2281 ();
 b15zdnd00an1n01x5 FILLER_63_2283 ();
 b15zdnd11an1n64x5 FILLER_64_8 ();
 b15zdnd11an1n64x5 FILLER_64_72 ();
 b15zdnd11an1n64x5 FILLER_64_136 ();
 b15zdnd11an1n64x5 FILLER_64_200 ();
 b15zdnd11an1n64x5 FILLER_64_264 ();
 b15zdnd11an1n64x5 FILLER_64_328 ();
 b15zdnd11an1n32x5 FILLER_64_392 ();
 b15zdnd11an1n16x5 FILLER_64_424 ();
 b15zdnd00an1n02x5 FILLER_64_440 ();
 b15zdnd11an1n64x5 FILLER_64_487 ();
 b15zdnd11an1n08x5 FILLER_64_551 ();
 b15zdnd00an1n02x5 FILLER_64_559 ();
 b15zdnd11an1n64x5 FILLER_64_603 ();
 b15zdnd11an1n32x5 FILLER_64_667 ();
 b15zdnd11an1n16x5 FILLER_64_699 ();
 b15zdnd00an1n02x5 FILLER_64_715 ();
 b15zdnd00an1n01x5 FILLER_64_717 ();
 b15zdnd11an1n64x5 FILLER_64_726 ();
 b15zdnd11an1n64x5 FILLER_64_790 ();
 b15zdnd11an1n64x5 FILLER_64_854 ();
 b15zdnd11an1n64x5 FILLER_64_918 ();
 b15zdnd11an1n64x5 FILLER_64_982 ();
 b15zdnd11an1n64x5 FILLER_64_1046 ();
 b15zdnd11an1n64x5 FILLER_64_1110 ();
 b15zdnd11an1n64x5 FILLER_64_1174 ();
 b15zdnd11an1n64x5 FILLER_64_1238 ();
 b15zdnd11an1n64x5 FILLER_64_1302 ();
 b15zdnd11an1n64x5 FILLER_64_1366 ();
 b15zdnd11an1n32x5 FILLER_64_1430 ();
 b15zdnd11an1n16x5 FILLER_64_1462 ();
 b15zdnd11an1n08x5 FILLER_64_2265 ();
 b15zdnd00an1n02x5 FILLER_64_2273 ();
 b15zdnd00an1n01x5 FILLER_64_2275 ();
 b15zdnd11an1n64x5 FILLER_65_0 ();
 b15zdnd11an1n64x5 FILLER_65_64 ();
 b15zdnd11an1n64x5 FILLER_65_128 ();
 b15zdnd11an1n64x5 FILLER_65_192 ();
 b15zdnd11an1n64x5 FILLER_65_256 ();
 b15zdnd11an1n64x5 FILLER_65_320 ();
 b15zdnd11an1n16x5 FILLER_65_384 ();
 b15zdnd00an1n02x5 FILLER_65_400 ();
 b15zdnd00an1n01x5 FILLER_65_402 ();
 b15zdnd11an1n64x5 FILLER_65_445 ();
 b15zdnd11an1n64x5 FILLER_65_509 ();
 b15zdnd11an1n64x5 FILLER_65_573 ();
 b15zdnd11an1n64x5 FILLER_65_637 ();
 b15zdnd11an1n64x5 FILLER_65_701 ();
 b15zdnd11an1n64x5 FILLER_65_765 ();
 b15zdnd11an1n64x5 FILLER_65_829 ();
 b15zdnd11an1n64x5 FILLER_65_893 ();
 b15zdnd11an1n08x5 FILLER_65_957 ();
 b15zdnd00an1n01x5 FILLER_65_965 ();
 b15zdnd11an1n64x5 FILLER_65_1010 ();
 b15zdnd11an1n64x5 FILLER_65_1074 ();
 b15zdnd11an1n64x5 FILLER_65_1138 ();
 b15zdnd11an1n64x5 FILLER_65_1202 ();
 b15zdnd11an1n64x5 FILLER_65_1266 ();
 b15zdnd11an1n64x5 FILLER_65_1330 ();
 b15zdnd11an1n64x5 FILLER_65_1394 ();
 b15zdnd11an1n16x5 FILLER_65_1458 ();
 b15zdnd11an1n08x5 FILLER_65_1474 ();
 b15zdnd11an1n04x5 FILLER_65_1482 ();
 b15zdnd11an1n16x5 FILLER_65_2257 ();
 b15zdnd11an1n08x5 FILLER_65_2273 ();
 b15zdnd00an1n02x5 FILLER_65_2281 ();
 b15zdnd00an1n01x5 FILLER_65_2283 ();
 b15zdnd11an1n64x5 FILLER_66_8 ();
 b15zdnd11an1n64x5 FILLER_66_72 ();
 b15zdnd11an1n64x5 FILLER_66_136 ();
 b15zdnd11an1n64x5 FILLER_66_200 ();
 b15zdnd11an1n64x5 FILLER_66_264 ();
 b15zdnd11an1n64x5 FILLER_66_328 ();
 b15zdnd11an1n64x5 FILLER_66_392 ();
 b15zdnd11an1n64x5 FILLER_66_456 ();
 b15zdnd11an1n64x5 FILLER_66_520 ();
 b15zdnd11an1n64x5 FILLER_66_584 ();
 b15zdnd11an1n64x5 FILLER_66_648 ();
 b15zdnd11an1n04x5 FILLER_66_712 ();
 b15zdnd00an1n02x5 FILLER_66_716 ();
 b15zdnd11an1n64x5 FILLER_66_726 ();
 b15zdnd11an1n04x5 FILLER_66_790 ();
 b15zdnd11an1n64x5 FILLER_66_802 ();
 b15zdnd11an1n64x5 FILLER_66_866 ();
 b15zdnd11an1n32x5 FILLER_66_930 ();
 b15zdnd11an1n16x5 FILLER_66_962 ();
 b15zdnd11an1n04x5 FILLER_66_978 ();
 b15zdnd00an1n02x5 FILLER_66_982 ();
 b15zdnd11an1n04x5 FILLER_66_987 ();
 b15zdnd11an1n64x5 FILLER_66_994 ();
 b15zdnd11an1n64x5 FILLER_66_1058 ();
 b15zdnd11an1n64x5 FILLER_66_1122 ();
 b15zdnd11an1n64x5 FILLER_66_1186 ();
 b15zdnd11an1n64x5 FILLER_66_1250 ();
 b15zdnd11an1n64x5 FILLER_66_1314 ();
 b15zdnd11an1n64x5 FILLER_66_1378 ();
 b15zdnd11an1n32x5 FILLER_66_1442 ();
 b15zdnd11an1n04x5 FILLER_66_1474 ();
 b15zdnd11an1n08x5 FILLER_66_2265 ();
 b15zdnd00an1n02x5 FILLER_66_2273 ();
 b15zdnd00an1n01x5 FILLER_66_2275 ();
 b15zdnd11an1n64x5 FILLER_67_0 ();
 b15zdnd11an1n64x5 FILLER_67_64 ();
 b15zdnd11an1n04x5 FILLER_67_128 ();
 b15zdnd00an1n02x5 FILLER_67_132 ();
 b15zdnd11an1n64x5 FILLER_67_153 ();
 b15zdnd11an1n64x5 FILLER_67_217 ();
 b15zdnd11an1n64x5 FILLER_67_281 ();
 b15zdnd11an1n64x5 FILLER_67_345 ();
 b15zdnd11an1n64x5 FILLER_67_409 ();
 b15zdnd11an1n64x5 FILLER_67_473 ();
 b15zdnd11an1n64x5 FILLER_67_537 ();
 b15zdnd11an1n64x5 FILLER_67_601 ();
 b15zdnd11an1n64x5 FILLER_67_665 ();
 b15zdnd11an1n64x5 FILLER_67_729 ();
 b15zdnd11an1n64x5 FILLER_67_793 ();
 b15zdnd11an1n64x5 FILLER_67_857 ();
 b15zdnd11an1n64x5 FILLER_67_921 ();
 b15zdnd00an1n02x5 FILLER_67_985 ();
 b15zdnd00an1n01x5 FILLER_67_987 ();
 b15zdnd11an1n64x5 FILLER_67_991 ();
 b15zdnd11an1n64x5 FILLER_67_1055 ();
 b15zdnd11an1n64x5 FILLER_67_1119 ();
 b15zdnd11an1n64x5 FILLER_67_1183 ();
 b15zdnd11an1n64x5 FILLER_67_1247 ();
 b15zdnd11an1n16x5 FILLER_67_1311 ();
 b15zdnd00an1n01x5 FILLER_67_1327 ();
 b15zdnd11an1n04x5 FILLER_67_1331 ();
 b15zdnd11an1n64x5 FILLER_67_1338 ();
 b15zdnd11an1n64x5 FILLER_67_1402 ();
 b15zdnd11an1n16x5 FILLER_67_1466 ();
 b15zdnd11an1n04x5 FILLER_67_1482 ();
 b15zdnd11an1n16x5 FILLER_67_2257 ();
 b15zdnd11an1n08x5 FILLER_67_2273 ();
 b15zdnd00an1n02x5 FILLER_67_2281 ();
 b15zdnd00an1n01x5 FILLER_67_2283 ();
 b15zdnd11an1n64x5 FILLER_68_8 ();
 b15zdnd11an1n64x5 FILLER_68_72 ();
 b15zdnd11an1n64x5 FILLER_68_136 ();
 b15zdnd11an1n64x5 FILLER_68_200 ();
 b15zdnd11an1n64x5 FILLER_68_264 ();
 b15zdnd11an1n64x5 FILLER_68_328 ();
 b15zdnd11an1n64x5 FILLER_68_392 ();
 b15zdnd11an1n64x5 FILLER_68_456 ();
 b15zdnd11an1n64x5 FILLER_68_520 ();
 b15zdnd11an1n64x5 FILLER_68_584 ();
 b15zdnd11an1n64x5 FILLER_68_648 ();
 b15zdnd11an1n04x5 FILLER_68_712 ();
 b15zdnd00an1n02x5 FILLER_68_716 ();
 b15zdnd11an1n64x5 FILLER_68_726 ();
 b15zdnd11an1n64x5 FILLER_68_790 ();
 b15zdnd11an1n16x5 FILLER_68_854 ();
 b15zdnd11an1n04x5 FILLER_68_870 ();
 b15zdnd00an1n02x5 FILLER_68_874 ();
 b15zdnd00an1n01x5 FILLER_68_876 ();
 b15zdnd11an1n32x5 FILLER_68_886 ();
 b15zdnd11an1n16x5 FILLER_68_918 ();
 b15zdnd11an1n08x5 FILLER_68_934 ();
 b15zdnd11an1n04x5 FILLER_68_942 ();
 b15zdnd00an1n01x5 FILLER_68_946 ();
 b15zdnd11an1n64x5 FILLER_68_991 ();
 b15zdnd11an1n64x5 FILLER_68_1055 ();
 b15zdnd11an1n64x5 FILLER_68_1119 ();
 b15zdnd11an1n64x5 FILLER_68_1183 ();
 b15zdnd11an1n32x5 FILLER_68_1247 ();
 b15zdnd11an1n08x5 FILLER_68_1279 ();
 b15zdnd11an1n04x5 FILLER_68_1287 ();
 b15zdnd00an1n02x5 FILLER_68_1291 ();
 b15zdnd00an1n01x5 FILLER_68_1293 ();
 b15zdnd11an1n64x5 FILLER_68_1303 ();
 b15zdnd11an1n64x5 FILLER_68_1367 ();
 b15zdnd11an1n32x5 FILLER_68_1431 ();
 b15zdnd11an1n08x5 FILLER_68_1463 ();
 b15zdnd11an1n04x5 FILLER_68_1471 ();
 b15zdnd00an1n02x5 FILLER_68_1475 ();
 b15zdnd00an1n01x5 FILLER_68_1477 ();
 b15zdnd11an1n08x5 FILLER_68_2265 ();
 b15zdnd00an1n02x5 FILLER_68_2273 ();
 b15zdnd00an1n01x5 FILLER_68_2275 ();
 b15zdnd11an1n64x5 FILLER_69_0 ();
 b15zdnd11an1n64x5 FILLER_69_64 ();
 b15zdnd11an1n64x5 FILLER_69_128 ();
 b15zdnd11an1n64x5 FILLER_69_192 ();
 b15zdnd11an1n64x5 FILLER_69_256 ();
 b15zdnd11an1n32x5 FILLER_69_320 ();
 b15zdnd11an1n16x5 FILLER_69_352 ();
 b15zdnd11an1n08x5 FILLER_69_368 ();
 b15zdnd11an1n04x5 FILLER_69_376 ();
 b15zdnd00an1n01x5 FILLER_69_380 ();
 b15zdnd11an1n64x5 FILLER_69_412 ();
 b15zdnd11an1n64x5 FILLER_69_476 ();
 b15zdnd11an1n64x5 FILLER_69_540 ();
 b15zdnd11an1n64x5 FILLER_69_604 ();
 b15zdnd11an1n64x5 FILLER_69_668 ();
 b15zdnd11an1n64x5 FILLER_69_732 ();
 b15zdnd11an1n64x5 FILLER_69_796 ();
 b15zdnd11an1n64x5 FILLER_69_860 ();
 b15zdnd11an1n32x5 FILLER_69_924 ();
 b15zdnd11an1n08x5 FILLER_69_956 ();
 b15zdnd11an1n04x5 FILLER_69_967 ();
 b15zdnd11an1n04x5 FILLER_69_974 ();
 b15zdnd11an1n64x5 FILLER_69_981 ();
 b15zdnd11an1n64x5 FILLER_69_1045 ();
 b15zdnd11an1n64x5 FILLER_69_1109 ();
 b15zdnd11an1n64x5 FILLER_69_1173 ();
 b15zdnd11an1n32x5 FILLER_69_1237 ();
 b15zdnd11an1n16x5 FILLER_69_1269 ();
 b15zdnd11an1n08x5 FILLER_69_1285 ();
 b15zdnd11an1n04x5 FILLER_69_1293 ();
 b15zdnd11an1n04x5 FILLER_69_1300 ();
 b15zdnd11an1n08x5 FILLER_69_1307 ();
 b15zdnd00an1n02x5 FILLER_69_1315 ();
 b15zdnd00an1n01x5 FILLER_69_1317 ();
 b15zdnd11an1n64x5 FILLER_69_1362 ();
 b15zdnd11an1n32x5 FILLER_69_1426 ();
 b15zdnd11an1n16x5 FILLER_69_1458 ();
 b15zdnd11an1n08x5 FILLER_69_1474 ();
 b15zdnd11an1n04x5 FILLER_69_1482 ();
 b15zdnd11an1n16x5 FILLER_69_2257 ();
 b15zdnd11an1n08x5 FILLER_69_2273 ();
 b15zdnd00an1n02x5 FILLER_69_2281 ();
 b15zdnd00an1n01x5 FILLER_69_2283 ();
 b15zdnd11an1n64x5 FILLER_70_8 ();
 b15zdnd11an1n64x5 FILLER_70_72 ();
 b15zdnd11an1n64x5 FILLER_70_136 ();
 b15zdnd11an1n64x5 FILLER_70_200 ();
 b15zdnd11an1n64x5 FILLER_70_264 ();
 b15zdnd11an1n64x5 FILLER_70_328 ();
 b15zdnd11an1n64x5 FILLER_70_392 ();
 b15zdnd11an1n64x5 FILLER_70_456 ();
 b15zdnd11an1n64x5 FILLER_70_520 ();
 b15zdnd11an1n64x5 FILLER_70_584 ();
 b15zdnd11an1n64x5 FILLER_70_648 ();
 b15zdnd11an1n04x5 FILLER_70_712 ();
 b15zdnd00an1n02x5 FILLER_70_716 ();
 b15zdnd11an1n64x5 FILLER_70_726 ();
 b15zdnd11an1n64x5 FILLER_70_790 ();
 b15zdnd11an1n64x5 FILLER_70_854 ();
 b15zdnd11an1n32x5 FILLER_70_918 ();
 b15zdnd11an1n08x5 FILLER_70_950 ();
 b15zdnd00an1n02x5 FILLER_70_958 ();
 b15zdnd00an1n01x5 FILLER_70_960 ();
 b15zdnd11an1n64x5 FILLER_70_1005 ();
 b15zdnd11an1n64x5 FILLER_70_1069 ();
 b15zdnd11an1n64x5 FILLER_70_1133 ();
 b15zdnd11an1n64x5 FILLER_70_1197 ();
 b15zdnd11an1n16x5 FILLER_70_1261 ();
 b15zdnd11an1n04x5 FILLER_70_1277 ();
 b15zdnd00an1n01x5 FILLER_70_1281 ();
 b15zdnd11an1n08x5 FILLER_70_1326 ();
 b15zdnd00an1n02x5 FILLER_70_1334 ();
 b15zdnd00an1n01x5 FILLER_70_1336 ();
 b15zdnd11an1n04x5 FILLER_70_1340 ();
 b15zdnd11an1n64x5 FILLER_70_1347 ();
 b15zdnd11an1n64x5 FILLER_70_1411 ();
 b15zdnd00an1n02x5 FILLER_70_1475 ();
 b15zdnd00an1n01x5 FILLER_70_1477 ();
 b15zdnd11an1n08x5 FILLER_70_2265 ();
 b15zdnd00an1n02x5 FILLER_70_2273 ();
 b15zdnd00an1n01x5 FILLER_70_2275 ();
 b15zdnd11an1n64x5 FILLER_71_0 ();
 b15zdnd11an1n64x5 FILLER_71_64 ();
 b15zdnd11an1n64x5 FILLER_71_128 ();
 b15zdnd11an1n64x5 FILLER_71_192 ();
 b15zdnd11an1n64x5 FILLER_71_256 ();
 b15zdnd11an1n64x5 FILLER_71_320 ();
 b15zdnd11an1n64x5 FILLER_71_384 ();
 b15zdnd11an1n64x5 FILLER_71_448 ();
 b15zdnd11an1n64x5 FILLER_71_512 ();
 b15zdnd11an1n08x5 FILLER_71_576 ();
 b15zdnd11an1n64x5 FILLER_71_626 ();
 b15zdnd11an1n64x5 FILLER_71_690 ();
 b15zdnd11an1n64x5 FILLER_71_754 ();
 b15zdnd11an1n64x5 FILLER_71_818 ();
 b15zdnd11an1n64x5 FILLER_71_882 ();
 b15zdnd11an1n64x5 FILLER_71_946 ();
 b15zdnd11an1n64x5 FILLER_71_1010 ();
 b15zdnd11an1n64x5 FILLER_71_1074 ();
 b15zdnd11an1n64x5 FILLER_71_1138 ();
 b15zdnd11an1n64x5 FILLER_71_1202 ();
 b15zdnd11an1n16x5 FILLER_71_1266 ();
 b15zdnd00an1n01x5 FILLER_71_1282 ();
 b15zdnd11an1n08x5 FILLER_71_1325 ();
 b15zdnd00an1n01x5 FILLER_71_1333 ();
 b15zdnd11an1n04x5 FILLER_71_1337 ();
 b15zdnd11an1n64x5 FILLER_71_1344 ();
 b15zdnd11an1n64x5 FILLER_71_1408 ();
 b15zdnd00an1n01x5 FILLER_71_1472 ();
 b15zdnd00an1n02x5 FILLER_71_1484 ();
 b15zdnd11an1n16x5 FILLER_71_2257 ();
 b15zdnd11an1n08x5 FILLER_71_2273 ();
 b15zdnd00an1n02x5 FILLER_71_2281 ();
 b15zdnd00an1n01x5 FILLER_71_2283 ();
 b15zdnd11an1n64x5 FILLER_72_8 ();
 b15zdnd11an1n64x5 FILLER_72_72 ();
 b15zdnd11an1n64x5 FILLER_72_136 ();
 b15zdnd00an1n01x5 FILLER_72_200 ();
 b15zdnd11an1n64x5 FILLER_72_234 ();
 b15zdnd11an1n64x5 FILLER_72_298 ();
 b15zdnd11an1n64x5 FILLER_72_362 ();
 b15zdnd11an1n64x5 FILLER_72_426 ();
 b15zdnd11an1n08x5 FILLER_72_490 ();
 b15zdnd11an1n04x5 FILLER_72_498 ();
 b15zdnd00an1n02x5 FILLER_72_502 ();
 b15zdnd11an1n64x5 FILLER_72_546 ();
 b15zdnd11an1n64x5 FILLER_72_610 ();
 b15zdnd11an1n32x5 FILLER_72_674 ();
 b15zdnd11an1n08x5 FILLER_72_706 ();
 b15zdnd11an1n04x5 FILLER_72_714 ();
 b15zdnd11an1n64x5 FILLER_72_726 ();
 b15zdnd11an1n64x5 FILLER_72_790 ();
 b15zdnd11an1n64x5 FILLER_72_854 ();
 b15zdnd11an1n16x5 FILLER_72_918 ();
 b15zdnd11an1n04x5 FILLER_72_978 ();
 b15zdnd11an1n64x5 FILLER_72_985 ();
 b15zdnd11an1n64x5 FILLER_72_1049 ();
 b15zdnd11an1n64x5 FILLER_72_1113 ();
 b15zdnd11an1n64x5 FILLER_72_1177 ();
 b15zdnd11an1n32x5 FILLER_72_1241 ();
 b15zdnd11an1n08x5 FILLER_72_1273 ();
 b15zdnd00an1n01x5 FILLER_72_1281 ();
 b15zdnd11an1n08x5 FILLER_72_1290 ();
 b15zdnd11an1n04x5 FILLER_72_1298 ();
 b15zdnd00an1n01x5 FILLER_72_1302 ();
 b15zdnd11an1n08x5 FILLER_72_1306 ();
 b15zdnd11an1n04x5 FILLER_72_1314 ();
 b15zdnd00an1n01x5 FILLER_72_1318 ();
 b15zdnd11an1n64x5 FILLER_72_1363 ();
 b15zdnd11an1n32x5 FILLER_72_1427 ();
 b15zdnd11an1n16x5 FILLER_72_1459 ();
 b15zdnd00an1n02x5 FILLER_72_1475 ();
 b15zdnd00an1n01x5 FILLER_72_1477 ();
 b15zdnd11an1n08x5 FILLER_72_2265 ();
 b15zdnd00an1n02x5 FILLER_72_2273 ();
 b15zdnd00an1n01x5 FILLER_72_2275 ();
 b15zdnd11an1n64x5 FILLER_73_0 ();
 b15zdnd11an1n64x5 FILLER_73_64 ();
 b15zdnd11an1n64x5 FILLER_73_128 ();
 b15zdnd11an1n64x5 FILLER_73_192 ();
 b15zdnd11an1n64x5 FILLER_73_256 ();
 b15zdnd11an1n64x5 FILLER_73_320 ();
 b15zdnd11an1n64x5 FILLER_73_384 ();
 b15zdnd11an1n64x5 FILLER_73_448 ();
 b15zdnd11an1n64x5 FILLER_73_512 ();
 b15zdnd11an1n64x5 FILLER_73_576 ();
 b15zdnd11an1n16x5 FILLER_73_640 ();
 b15zdnd11an1n08x5 FILLER_73_656 ();
 b15zdnd11an1n04x5 FILLER_73_664 ();
 b15zdnd11an1n08x5 FILLER_73_671 ();
 b15zdnd00an1n02x5 FILLER_73_679 ();
 b15zdnd00an1n01x5 FILLER_73_681 ();
 b15zdnd11an1n64x5 FILLER_73_691 ();
 b15zdnd11an1n64x5 FILLER_73_755 ();
 b15zdnd11an1n64x5 FILLER_73_819 ();
 b15zdnd11an1n64x5 FILLER_73_883 ();
 b15zdnd11an1n04x5 FILLER_73_947 ();
 b15zdnd11an1n04x5 FILLER_73_954 ();
 b15zdnd11an1n08x5 FILLER_73_961 ();
 b15zdnd00an1n02x5 FILLER_73_969 ();
 b15zdnd00an1n01x5 FILLER_73_971 ();
 b15zdnd11an1n04x5 FILLER_73_975 ();
 b15zdnd11an1n64x5 FILLER_73_982 ();
 b15zdnd11an1n64x5 FILLER_73_1046 ();
 b15zdnd11an1n64x5 FILLER_73_1110 ();
 b15zdnd11an1n64x5 FILLER_73_1174 ();
 b15zdnd11an1n64x5 FILLER_73_1238 ();
 b15zdnd11an1n64x5 FILLER_73_1302 ();
 b15zdnd11an1n64x5 FILLER_73_1366 ();
 b15zdnd11an1n32x5 FILLER_73_1430 ();
 b15zdnd11an1n16x5 FILLER_73_1462 ();
 b15zdnd11an1n08x5 FILLER_73_1478 ();
 b15zdnd11an1n16x5 FILLER_73_2257 ();
 b15zdnd11an1n08x5 FILLER_73_2273 ();
 b15zdnd00an1n02x5 FILLER_73_2281 ();
 b15zdnd00an1n01x5 FILLER_73_2283 ();
 b15zdnd11an1n64x5 FILLER_74_8 ();
 b15zdnd11an1n64x5 FILLER_74_72 ();
 b15zdnd11an1n64x5 FILLER_74_136 ();
 b15zdnd11an1n64x5 FILLER_74_200 ();
 b15zdnd11an1n64x5 FILLER_74_264 ();
 b15zdnd11an1n64x5 FILLER_74_328 ();
 b15zdnd11an1n64x5 FILLER_74_392 ();
 b15zdnd11an1n64x5 FILLER_74_456 ();
 b15zdnd11an1n64x5 FILLER_74_520 ();
 b15zdnd11an1n64x5 FILLER_74_584 ();
 b15zdnd11an1n08x5 FILLER_74_648 ();
 b15zdnd00an1n01x5 FILLER_74_656 ();
 b15zdnd11an1n04x5 FILLER_74_660 ();
 b15zdnd11an1n16x5 FILLER_74_689 ();
 b15zdnd11an1n08x5 FILLER_74_705 ();
 b15zdnd11an1n04x5 FILLER_74_713 ();
 b15zdnd00an1n01x5 FILLER_74_717 ();
 b15zdnd11an1n64x5 FILLER_74_726 ();
 b15zdnd11an1n32x5 FILLER_74_790 ();
 b15zdnd11an1n16x5 FILLER_74_822 ();
 b15zdnd11an1n08x5 FILLER_74_838 ();
 b15zdnd00an1n02x5 FILLER_74_846 ();
 b15zdnd11an1n32x5 FILLER_74_890 ();
 b15zdnd11an1n16x5 FILLER_74_922 ();
 b15zdnd11an1n08x5 FILLER_74_938 ();
 b15zdnd11an1n04x5 FILLER_74_946 ();
 b15zdnd11an1n64x5 FILLER_74_953 ();
 b15zdnd11an1n64x5 FILLER_74_1017 ();
 b15zdnd11an1n64x5 FILLER_74_1081 ();
 b15zdnd11an1n64x5 FILLER_74_1145 ();
 b15zdnd11an1n64x5 FILLER_74_1209 ();
 b15zdnd11an1n64x5 FILLER_74_1273 ();
 b15zdnd11an1n64x5 FILLER_74_1337 ();
 b15zdnd11an1n64x5 FILLER_74_1401 ();
 b15zdnd11an1n08x5 FILLER_74_1465 ();
 b15zdnd11an1n04x5 FILLER_74_1473 ();
 b15zdnd00an1n01x5 FILLER_74_1477 ();
 b15zdnd11an1n08x5 FILLER_74_2265 ();
 b15zdnd00an1n02x5 FILLER_74_2273 ();
 b15zdnd00an1n01x5 FILLER_74_2275 ();
 b15zdnd11an1n64x5 FILLER_75_0 ();
 b15zdnd11an1n64x5 FILLER_75_64 ();
 b15zdnd11an1n64x5 FILLER_75_128 ();
 b15zdnd11an1n64x5 FILLER_75_192 ();
 b15zdnd11an1n64x5 FILLER_75_256 ();
 b15zdnd11an1n64x5 FILLER_75_320 ();
 b15zdnd11an1n64x5 FILLER_75_384 ();
 b15zdnd11an1n64x5 FILLER_75_448 ();
 b15zdnd11an1n64x5 FILLER_75_512 ();
 b15zdnd11an1n64x5 FILLER_75_576 ();
 b15zdnd00an1n02x5 FILLER_75_640 ();
 b15zdnd00an1n01x5 FILLER_75_642 ();
 b15zdnd11an1n64x5 FILLER_75_646 ();
 b15zdnd11an1n64x5 FILLER_75_710 ();
 b15zdnd11an1n16x5 FILLER_75_774 ();
 b15zdnd11an1n08x5 FILLER_75_790 ();
 b15zdnd11an1n32x5 FILLER_75_807 ();
 b15zdnd11an1n08x5 FILLER_75_839 ();
 b15zdnd00an1n02x5 FILLER_75_847 ();
 b15zdnd11an1n64x5 FILLER_75_891 ();
 b15zdnd11an1n64x5 FILLER_75_955 ();
 b15zdnd11an1n64x5 FILLER_75_1019 ();
 b15zdnd11an1n64x5 FILLER_75_1083 ();
 b15zdnd11an1n64x5 FILLER_75_1147 ();
 b15zdnd11an1n64x5 FILLER_75_1211 ();
 b15zdnd11an1n64x5 FILLER_75_1275 ();
 b15zdnd11an1n64x5 FILLER_75_1339 ();
 b15zdnd11an1n64x5 FILLER_75_1403 ();
 b15zdnd11an1n16x5 FILLER_75_1467 ();
 b15zdnd00an1n02x5 FILLER_75_1483 ();
 b15zdnd00an1n01x5 FILLER_75_1485 ();
 b15zdnd11an1n16x5 FILLER_75_2257 ();
 b15zdnd11an1n08x5 FILLER_75_2273 ();
 b15zdnd00an1n02x5 FILLER_75_2281 ();
 b15zdnd00an1n01x5 FILLER_75_2283 ();
 b15zdnd11an1n64x5 FILLER_76_8 ();
 b15zdnd11an1n64x5 FILLER_76_72 ();
 b15zdnd11an1n64x5 FILLER_76_136 ();
 b15zdnd11an1n64x5 FILLER_76_200 ();
 b15zdnd11an1n64x5 FILLER_76_264 ();
 b15zdnd11an1n32x5 FILLER_76_328 ();
 b15zdnd11an1n16x5 FILLER_76_360 ();
 b15zdnd11an1n08x5 FILLER_76_376 ();
 b15zdnd11an1n04x5 FILLER_76_384 ();
 b15zdnd00an1n02x5 FILLER_76_388 ();
 b15zdnd00an1n01x5 FILLER_76_390 ();
 b15zdnd11an1n64x5 FILLER_76_436 ();
 b15zdnd11an1n32x5 FILLER_76_500 ();
 b15zdnd11an1n16x5 FILLER_76_532 ();
 b15zdnd11an1n08x5 FILLER_76_548 ();
 b15zdnd11an1n04x5 FILLER_76_556 ();
 b15zdnd11an1n16x5 FILLER_76_602 ();
 b15zdnd11an1n08x5 FILLER_76_618 ();
 b15zdnd00an1n02x5 FILLER_76_626 ();
 b15zdnd00an1n01x5 FILLER_76_628 ();
 b15zdnd11an1n04x5 FILLER_76_632 ();
 b15zdnd11an1n32x5 FILLER_76_661 ();
 b15zdnd11an1n16x5 FILLER_76_693 ();
 b15zdnd11an1n08x5 FILLER_76_709 ();
 b15zdnd00an1n01x5 FILLER_76_717 ();
 b15zdnd11an1n64x5 FILLER_76_726 ();
 b15zdnd11an1n64x5 FILLER_76_790 ();
 b15zdnd11an1n04x5 FILLER_76_854 ();
 b15zdnd00an1n02x5 FILLER_76_858 ();
 b15zdnd11an1n64x5 FILLER_76_902 ();
 b15zdnd11an1n64x5 FILLER_76_966 ();
 b15zdnd11an1n64x5 FILLER_76_1030 ();
 b15zdnd11an1n64x5 FILLER_76_1094 ();
 b15zdnd11an1n64x5 FILLER_76_1158 ();
 b15zdnd11an1n64x5 FILLER_76_1222 ();
 b15zdnd11an1n64x5 FILLER_76_1286 ();
 b15zdnd11an1n64x5 FILLER_76_1350 ();
 b15zdnd11an1n64x5 FILLER_76_1414 ();
 b15zdnd11an1n08x5 FILLER_76_2265 ();
 b15zdnd00an1n02x5 FILLER_76_2273 ();
 b15zdnd00an1n01x5 FILLER_76_2275 ();
 b15zdnd11an1n64x5 FILLER_77_0 ();
 b15zdnd11an1n64x5 FILLER_77_64 ();
 b15zdnd11an1n64x5 FILLER_77_128 ();
 b15zdnd11an1n64x5 FILLER_77_192 ();
 b15zdnd11an1n64x5 FILLER_77_256 ();
 b15zdnd11an1n64x5 FILLER_77_320 ();
 b15zdnd11an1n64x5 FILLER_77_384 ();
 b15zdnd11an1n64x5 FILLER_77_448 ();
 b15zdnd11an1n64x5 FILLER_77_512 ();
 b15zdnd11an1n64x5 FILLER_77_576 ();
 b15zdnd11an1n64x5 FILLER_77_640 ();
 b15zdnd11an1n64x5 FILLER_77_704 ();
 b15zdnd11an1n64x5 FILLER_77_768 ();
 b15zdnd11an1n16x5 FILLER_77_832 ();
 b15zdnd11an1n08x5 FILLER_77_848 ();
 b15zdnd11an1n04x5 FILLER_77_856 ();
 b15zdnd11an1n64x5 FILLER_77_902 ();
 b15zdnd11an1n32x5 FILLER_77_966 ();
 b15zdnd11an1n16x5 FILLER_77_998 ();
 b15zdnd11an1n08x5 FILLER_77_1014 ();
 b15zdnd11an1n04x5 FILLER_77_1022 ();
 b15zdnd00an1n01x5 FILLER_77_1026 ();
 b15zdnd11an1n64x5 FILLER_77_1069 ();
 b15zdnd11an1n64x5 FILLER_77_1133 ();
 b15zdnd11an1n64x5 FILLER_77_1197 ();
 b15zdnd11an1n32x5 FILLER_77_1261 ();
 b15zdnd11an1n08x5 FILLER_77_1293 ();
 b15zdnd00an1n02x5 FILLER_77_1301 ();
 b15zdnd00an1n01x5 FILLER_77_1303 ();
 b15zdnd11an1n64x5 FILLER_77_1313 ();
 b15zdnd11an1n64x5 FILLER_77_1377 ();
 b15zdnd11an1n32x5 FILLER_77_1441 ();
 b15zdnd11an1n08x5 FILLER_77_1473 ();
 b15zdnd11an1n04x5 FILLER_77_1481 ();
 b15zdnd00an1n01x5 FILLER_77_1485 ();
 b15zdnd11an1n16x5 FILLER_77_2257 ();
 b15zdnd11an1n08x5 FILLER_77_2273 ();
 b15zdnd00an1n02x5 FILLER_77_2281 ();
 b15zdnd00an1n01x5 FILLER_77_2283 ();
 b15zdnd11an1n64x5 FILLER_78_8 ();
 b15zdnd11an1n64x5 FILLER_78_72 ();
 b15zdnd11an1n64x5 FILLER_78_136 ();
 b15zdnd11an1n64x5 FILLER_78_200 ();
 b15zdnd11an1n64x5 FILLER_78_264 ();
 b15zdnd11an1n64x5 FILLER_78_328 ();
 b15zdnd11an1n64x5 FILLER_78_392 ();
 b15zdnd11an1n64x5 FILLER_78_456 ();
 b15zdnd11an1n64x5 FILLER_78_520 ();
 b15zdnd11an1n64x5 FILLER_78_584 ();
 b15zdnd11an1n64x5 FILLER_78_648 ();
 b15zdnd11an1n04x5 FILLER_78_712 ();
 b15zdnd00an1n02x5 FILLER_78_716 ();
 b15zdnd11an1n64x5 FILLER_78_726 ();
 b15zdnd11an1n32x5 FILLER_78_790 ();
 b15zdnd11an1n16x5 FILLER_78_822 ();
 b15zdnd11an1n08x5 FILLER_78_838 ();
 b15zdnd11an1n64x5 FILLER_78_888 ();
 b15zdnd11an1n64x5 FILLER_78_952 ();
 b15zdnd11an1n64x5 FILLER_78_1016 ();
 b15zdnd11an1n64x5 FILLER_78_1080 ();
 b15zdnd11an1n64x5 FILLER_78_1144 ();
 b15zdnd11an1n64x5 FILLER_78_1208 ();
 b15zdnd11an1n16x5 FILLER_78_1272 ();
 b15zdnd11an1n04x5 FILLER_78_1288 ();
 b15zdnd00an1n02x5 FILLER_78_1292 ();
 b15zdnd11an1n32x5 FILLER_78_1303 ();
 b15zdnd11an1n16x5 FILLER_78_1335 ();
 b15zdnd11an1n08x5 FILLER_78_1351 ();
 b15zdnd11an1n04x5 FILLER_78_1359 ();
 b15zdnd11an1n64x5 FILLER_78_1405 ();
 b15zdnd11an1n08x5 FILLER_78_1469 ();
 b15zdnd00an1n01x5 FILLER_78_1477 ();
 b15zdnd11an1n08x5 FILLER_78_2265 ();
 b15zdnd00an1n02x5 FILLER_78_2273 ();
 b15zdnd00an1n01x5 FILLER_78_2275 ();
 b15zdnd11an1n64x5 FILLER_79_0 ();
 b15zdnd11an1n64x5 FILLER_79_64 ();
 b15zdnd11an1n64x5 FILLER_79_128 ();
 b15zdnd11an1n64x5 FILLER_79_192 ();
 b15zdnd11an1n64x5 FILLER_79_256 ();
 b15zdnd11an1n64x5 FILLER_79_320 ();
 b15zdnd11an1n64x5 FILLER_79_384 ();
 b15zdnd11an1n64x5 FILLER_79_448 ();
 b15zdnd11an1n32x5 FILLER_79_512 ();
 b15zdnd11an1n16x5 FILLER_79_544 ();
 b15zdnd11an1n08x5 FILLER_79_560 ();
 b15zdnd11an1n04x5 FILLER_79_568 ();
 b15zdnd00an1n02x5 FILLER_79_572 ();
 b15zdnd00an1n01x5 FILLER_79_574 ();
 b15zdnd11an1n64x5 FILLER_79_617 ();
 b15zdnd11an1n64x5 FILLER_79_681 ();
 b15zdnd11an1n64x5 FILLER_79_745 ();
 b15zdnd11an1n64x5 FILLER_79_809 ();
 b15zdnd11an1n64x5 FILLER_79_873 ();
 b15zdnd11an1n64x5 FILLER_79_937 ();
 b15zdnd11an1n64x5 FILLER_79_1001 ();
 b15zdnd11an1n64x5 FILLER_79_1065 ();
 b15zdnd11an1n64x5 FILLER_79_1129 ();
 b15zdnd11an1n64x5 FILLER_79_1193 ();
 b15zdnd11an1n64x5 FILLER_79_1257 ();
 b15zdnd11an1n32x5 FILLER_79_1321 ();
 b15zdnd11an1n08x5 FILLER_79_1353 ();
 b15zdnd11an1n04x5 FILLER_79_1361 ();
 b15zdnd00an1n01x5 FILLER_79_1365 ();
 b15zdnd11an1n64x5 FILLER_79_1408 ();
 b15zdnd11an1n08x5 FILLER_79_1472 ();
 b15zdnd11an1n04x5 FILLER_79_1480 ();
 b15zdnd00an1n02x5 FILLER_79_1484 ();
 b15zdnd11an1n16x5 FILLER_79_2257 ();
 b15zdnd11an1n08x5 FILLER_79_2273 ();
 b15zdnd00an1n02x5 FILLER_79_2281 ();
 b15zdnd00an1n01x5 FILLER_79_2283 ();
 b15zdnd11an1n64x5 FILLER_80_8 ();
 b15zdnd11an1n64x5 FILLER_80_72 ();
 b15zdnd11an1n64x5 FILLER_80_136 ();
 b15zdnd11an1n64x5 FILLER_80_200 ();
 b15zdnd11an1n64x5 FILLER_80_264 ();
 b15zdnd11an1n64x5 FILLER_80_328 ();
 b15zdnd00an1n02x5 FILLER_80_392 ();
 b15zdnd00an1n01x5 FILLER_80_394 ();
 b15zdnd11an1n32x5 FILLER_80_415 ();
 b15zdnd00an1n02x5 FILLER_80_447 ();
 b15zdnd11an1n32x5 FILLER_80_494 ();
 b15zdnd11an1n08x5 FILLER_80_526 ();
 b15zdnd11an1n04x5 FILLER_80_534 ();
 b15zdnd11an1n64x5 FILLER_80_580 ();
 b15zdnd11an1n08x5 FILLER_80_644 ();
 b15zdnd00an1n01x5 FILLER_80_652 ();
 b15zdnd11an1n32x5 FILLER_80_656 ();
 b15zdnd11an1n16x5 FILLER_80_688 ();
 b15zdnd11an1n08x5 FILLER_80_704 ();
 b15zdnd11an1n04x5 FILLER_80_712 ();
 b15zdnd00an1n02x5 FILLER_80_716 ();
 b15zdnd11an1n64x5 FILLER_80_726 ();
 b15zdnd11an1n64x5 FILLER_80_790 ();
 b15zdnd11an1n64x5 FILLER_80_854 ();
 b15zdnd11an1n64x5 FILLER_80_918 ();
 b15zdnd11an1n64x5 FILLER_80_982 ();
 b15zdnd11an1n64x5 FILLER_80_1046 ();
 b15zdnd11an1n64x5 FILLER_80_1110 ();
 b15zdnd11an1n64x5 FILLER_80_1174 ();
 b15zdnd11an1n64x5 FILLER_80_1238 ();
 b15zdnd11an1n04x5 FILLER_80_1302 ();
 b15zdnd00an1n01x5 FILLER_80_1306 ();
 b15zdnd11an1n64x5 FILLER_80_1310 ();
 b15zdnd11an1n64x5 FILLER_80_1374 ();
 b15zdnd11an1n32x5 FILLER_80_1438 ();
 b15zdnd11an1n08x5 FILLER_80_1470 ();
 b15zdnd11an1n08x5 FILLER_80_2265 ();
 b15zdnd00an1n02x5 FILLER_80_2273 ();
 b15zdnd00an1n01x5 FILLER_80_2275 ();
 b15zdnd11an1n64x5 FILLER_81_0 ();
 b15zdnd11an1n64x5 FILLER_81_64 ();
 b15zdnd11an1n64x5 FILLER_81_128 ();
 b15zdnd11an1n64x5 FILLER_81_192 ();
 b15zdnd11an1n64x5 FILLER_81_256 ();
 b15zdnd11an1n64x5 FILLER_81_320 ();
 b15zdnd11an1n64x5 FILLER_81_384 ();
 b15zdnd11an1n64x5 FILLER_81_448 ();
 b15zdnd11an1n64x5 FILLER_81_512 ();
 b15zdnd11an1n32x5 FILLER_81_576 ();
 b15zdnd11an1n16x5 FILLER_81_608 ();
 b15zdnd11an1n08x5 FILLER_81_624 ();
 b15zdnd11an1n64x5 FILLER_81_676 ();
 b15zdnd11an1n64x5 FILLER_81_740 ();
 b15zdnd11an1n64x5 FILLER_81_804 ();
 b15zdnd11an1n64x5 FILLER_81_868 ();
 b15zdnd11an1n64x5 FILLER_81_932 ();
 b15zdnd11an1n64x5 FILLER_81_996 ();
 b15zdnd11an1n64x5 FILLER_81_1060 ();
 b15zdnd11an1n64x5 FILLER_81_1124 ();
 b15zdnd11an1n64x5 FILLER_81_1188 ();
 b15zdnd11an1n16x5 FILLER_81_1252 ();
 b15zdnd11an1n08x5 FILLER_81_1268 ();
 b15zdnd11an1n04x5 FILLER_81_1276 ();
 b15zdnd11an1n64x5 FILLER_81_1324 ();
 b15zdnd11an1n64x5 FILLER_81_1388 ();
 b15zdnd11an1n16x5 FILLER_81_1452 ();
 b15zdnd11an1n04x5 FILLER_81_1468 ();
 b15zdnd00an1n01x5 FILLER_81_1472 ();
 b15zdnd00an1n02x5 FILLER_81_1484 ();
 b15zdnd11an1n16x5 FILLER_81_2257 ();
 b15zdnd11an1n08x5 FILLER_81_2273 ();
 b15zdnd00an1n02x5 FILLER_81_2281 ();
 b15zdnd00an1n01x5 FILLER_81_2283 ();
 b15zdnd11an1n64x5 FILLER_82_8 ();
 b15zdnd11an1n64x5 FILLER_82_72 ();
 b15zdnd11an1n64x5 FILLER_82_136 ();
 b15zdnd11an1n64x5 FILLER_82_200 ();
 b15zdnd11an1n64x5 FILLER_82_264 ();
 b15zdnd11an1n64x5 FILLER_82_328 ();
 b15zdnd11an1n32x5 FILLER_82_392 ();
 b15zdnd11an1n08x5 FILLER_82_424 ();
 b15zdnd11an1n04x5 FILLER_82_432 ();
 b15zdnd00an1n01x5 FILLER_82_436 ();
 b15zdnd11an1n64x5 FILLER_82_482 ();
 b15zdnd11an1n64x5 FILLER_82_546 ();
 b15zdnd11an1n32x5 FILLER_82_610 ();
 b15zdnd00an1n02x5 FILLER_82_642 ();
 b15zdnd00an1n01x5 FILLER_82_644 ();
 b15zdnd11an1n16x5 FILLER_82_687 ();
 b15zdnd11an1n08x5 FILLER_82_703 ();
 b15zdnd11an1n04x5 FILLER_82_711 ();
 b15zdnd00an1n02x5 FILLER_82_715 ();
 b15zdnd00an1n01x5 FILLER_82_717 ();
 b15zdnd11an1n64x5 FILLER_82_726 ();
 b15zdnd11an1n64x5 FILLER_82_790 ();
 b15zdnd11an1n64x5 FILLER_82_854 ();
 b15zdnd11an1n64x5 FILLER_82_918 ();
 b15zdnd11an1n64x5 FILLER_82_982 ();
 b15zdnd11an1n64x5 FILLER_82_1046 ();
 b15zdnd11an1n64x5 FILLER_82_1110 ();
 b15zdnd11an1n64x5 FILLER_82_1174 ();
 b15zdnd11an1n32x5 FILLER_82_1238 ();
 b15zdnd11an1n16x5 FILLER_82_1270 ();
 b15zdnd11an1n08x5 FILLER_82_1286 ();
 b15zdnd11an1n04x5 FILLER_82_1294 ();
 b15zdnd00an1n01x5 FILLER_82_1298 ();
 b15zdnd11an1n64x5 FILLER_82_1343 ();
 b15zdnd11an1n64x5 FILLER_82_1407 ();
 b15zdnd11an1n04x5 FILLER_82_1471 ();
 b15zdnd00an1n02x5 FILLER_82_1475 ();
 b15zdnd00an1n01x5 FILLER_82_1477 ();
 b15zdnd11an1n08x5 FILLER_82_2265 ();
 b15zdnd00an1n02x5 FILLER_82_2273 ();
 b15zdnd00an1n01x5 FILLER_82_2275 ();
 b15zdnd11an1n64x5 FILLER_83_0 ();
 b15zdnd11an1n64x5 FILLER_83_64 ();
 b15zdnd11an1n64x5 FILLER_83_128 ();
 b15zdnd11an1n64x5 FILLER_83_192 ();
 b15zdnd11an1n64x5 FILLER_83_256 ();
 b15zdnd11an1n64x5 FILLER_83_320 ();
 b15zdnd11an1n64x5 FILLER_83_384 ();
 b15zdnd11an1n64x5 FILLER_83_448 ();
 b15zdnd11an1n64x5 FILLER_83_512 ();
 b15zdnd11an1n64x5 FILLER_83_576 ();
 b15zdnd11an1n08x5 FILLER_83_640 ();
 b15zdnd11an1n04x5 FILLER_83_648 ();
 b15zdnd11an1n04x5 FILLER_83_655 ();
 b15zdnd00an1n02x5 FILLER_83_659 ();
 b15zdnd11an1n64x5 FILLER_83_664 ();
 b15zdnd11an1n64x5 FILLER_83_728 ();
 b15zdnd11an1n64x5 FILLER_83_792 ();
 b15zdnd11an1n64x5 FILLER_83_856 ();
 b15zdnd11an1n64x5 FILLER_83_920 ();
 b15zdnd11an1n64x5 FILLER_83_984 ();
 b15zdnd11an1n64x5 FILLER_83_1048 ();
 b15zdnd11an1n64x5 FILLER_83_1112 ();
 b15zdnd11an1n64x5 FILLER_83_1176 ();
 b15zdnd11an1n32x5 FILLER_83_1240 ();
 b15zdnd11an1n08x5 FILLER_83_1272 ();
 b15zdnd11an1n04x5 FILLER_83_1324 ();
 b15zdnd11an1n04x5 FILLER_83_1331 ();
 b15zdnd11an1n64x5 FILLER_83_1338 ();
 b15zdnd11an1n64x5 FILLER_83_1402 ();
 b15zdnd11an1n16x5 FILLER_83_1466 ();
 b15zdnd11an1n04x5 FILLER_83_1482 ();
 b15zdnd11an1n16x5 FILLER_83_2257 ();
 b15zdnd11an1n08x5 FILLER_83_2273 ();
 b15zdnd00an1n02x5 FILLER_83_2281 ();
 b15zdnd00an1n01x5 FILLER_83_2283 ();
 b15zdnd11an1n64x5 FILLER_84_8 ();
 b15zdnd11an1n64x5 FILLER_84_72 ();
 b15zdnd11an1n64x5 FILLER_84_136 ();
 b15zdnd11an1n64x5 FILLER_84_200 ();
 b15zdnd11an1n64x5 FILLER_84_264 ();
 b15zdnd11an1n64x5 FILLER_84_328 ();
 b15zdnd00an1n02x5 FILLER_84_392 ();
 b15zdnd11an1n64x5 FILLER_84_402 ();
 b15zdnd11an1n64x5 FILLER_84_466 ();
 b15zdnd11an1n64x5 FILLER_84_530 ();
 b15zdnd11an1n64x5 FILLER_84_594 ();
 b15zdnd11an1n32x5 FILLER_84_658 ();
 b15zdnd11an1n16x5 FILLER_84_690 ();
 b15zdnd11an1n08x5 FILLER_84_706 ();
 b15zdnd11an1n04x5 FILLER_84_714 ();
 b15zdnd11an1n64x5 FILLER_84_726 ();
 b15zdnd11an1n64x5 FILLER_84_790 ();
 b15zdnd11an1n64x5 FILLER_84_854 ();
 b15zdnd11an1n64x5 FILLER_84_918 ();
 b15zdnd11an1n64x5 FILLER_84_982 ();
 b15zdnd11an1n64x5 FILLER_84_1046 ();
 b15zdnd11an1n64x5 FILLER_84_1110 ();
 b15zdnd11an1n64x5 FILLER_84_1174 ();
 b15zdnd11an1n16x5 FILLER_84_1238 ();
 b15zdnd11an1n08x5 FILLER_84_1254 ();
 b15zdnd00an1n02x5 FILLER_84_1262 ();
 b15zdnd00an1n01x5 FILLER_84_1264 ();
 b15zdnd11an1n04x5 FILLER_84_1272 ();
 b15zdnd11an1n04x5 FILLER_84_1320 ();
 b15zdnd11an1n04x5 FILLER_84_1327 ();
 b15zdnd11an1n04x5 FILLER_84_1334 ();
 b15zdnd11an1n04x5 FILLER_84_1341 ();
 b15zdnd11an1n16x5 FILLER_84_1348 ();
 b15zdnd11an1n04x5 FILLER_84_1364 ();
 b15zdnd11an1n64x5 FILLER_84_1376 ();
 b15zdnd11an1n32x5 FILLER_84_1440 ();
 b15zdnd11an1n04x5 FILLER_84_1472 ();
 b15zdnd00an1n02x5 FILLER_84_1476 ();
 b15zdnd11an1n08x5 FILLER_84_2265 ();
 b15zdnd00an1n02x5 FILLER_84_2273 ();
 b15zdnd00an1n01x5 FILLER_84_2275 ();
 b15zdnd11an1n64x5 FILLER_85_0 ();
 b15zdnd11an1n64x5 FILLER_85_64 ();
 b15zdnd11an1n64x5 FILLER_85_128 ();
 b15zdnd11an1n64x5 FILLER_85_192 ();
 b15zdnd11an1n64x5 FILLER_85_256 ();
 b15zdnd11an1n64x5 FILLER_85_320 ();
 b15zdnd11an1n64x5 FILLER_85_384 ();
 b15zdnd11an1n64x5 FILLER_85_448 ();
 b15zdnd11an1n64x5 FILLER_85_512 ();
 b15zdnd11an1n64x5 FILLER_85_576 ();
 b15zdnd11an1n64x5 FILLER_85_640 ();
 b15zdnd11an1n64x5 FILLER_85_704 ();
 b15zdnd11an1n64x5 FILLER_85_768 ();
 b15zdnd11an1n64x5 FILLER_85_832 ();
 b15zdnd11an1n64x5 FILLER_85_896 ();
 b15zdnd11an1n64x5 FILLER_85_960 ();
 b15zdnd11an1n64x5 FILLER_85_1024 ();
 b15zdnd11an1n64x5 FILLER_85_1088 ();
 b15zdnd11an1n64x5 FILLER_85_1152 ();
 b15zdnd11an1n32x5 FILLER_85_1216 ();
 b15zdnd11an1n16x5 FILLER_85_1248 ();
 b15zdnd11an1n08x5 FILLER_85_1264 ();
 b15zdnd00an1n02x5 FILLER_85_1272 ();
 b15zdnd11an1n04x5 FILLER_85_1316 ();
 b15zdnd11an1n04x5 FILLER_85_1323 ();
 b15zdnd11an1n04x5 FILLER_85_1330 ();
 b15zdnd11an1n64x5 FILLER_85_1337 ();
 b15zdnd11an1n64x5 FILLER_85_1401 ();
 b15zdnd11an1n16x5 FILLER_85_1465 ();
 b15zdnd11an1n04x5 FILLER_85_1481 ();
 b15zdnd00an1n01x5 FILLER_85_1485 ();
 b15zdnd11an1n16x5 FILLER_85_2257 ();
 b15zdnd11an1n08x5 FILLER_85_2273 ();
 b15zdnd00an1n02x5 FILLER_85_2281 ();
 b15zdnd00an1n01x5 FILLER_85_2283 ();
 b15zdnd11an1n64x5 FILLER_86_8 ();
 b15zdnd11an1n64x5 FILLER_86_72 ();
 b15zdnd11an1n64x5 FILLER_86_136 ();
 b15zdnd11an1n64x5 FILLER_86_200 ();
 b15zdnd11an1n64x5 FILLER_86_264 ();
 b15zdnd11an1n64x5 FILLER_86_328 ();
 b15zdnd11an1n64x5 FILLER_86_392 ();
 b15zdnd11an1n64x5 FILLER_86_456 ();
 b15zdnd11an1n64x5 FILLER_86_520 ();
 b15zdnd11an1n64x5 FILLER_86_584 ();
 b15zdnd11an1n64x5 FILLER_86_648 ();
 b15zdnd11an1n04x5 FILLER_86_712 ();
 b15zdnd00an1n02x5 FILLER_86_716 ();
 b15zdnd11an1n64x5 FILLER_86_726 ();
 b15zdnd11an1n64x5 FILLER_86_790 ();
 b15zdnd11an1n64x5 FILLER_86_854 ();
 b15zdnd11an1n64x5 FILLER_86_918 ();
 b15zdnd11an1n64x5 FILLER_86_982 ();
 b15zdnd11an1n64x5 FILLER_86_1046 ();
 b15zdnd11an1n64x5 FILLER_86_1110 ();
 b15zdnd11an1n64x5 FILLER_86_1174 ();
 b15zdnd11an1n32x5 FILLER_86_1238 ();
 b15zdnd11an1n16x5 FILLER_86_1270 ();
 b15zdnd11an1n04x5 FILLER_86_1286 ();
 b15zdnd00an1n02x5 FILLER_86_1290 ();
 b15zdnd11an1n04x5 FILLER_86_1295 ();
 b15zdnd11an1n04x5 FILLER_86_1302 ();
 b15zdnd11an1n04x5 FILLER_86_1309 ();
 b15zdnd11an1n04x5 FILLER_86_1316 ();
 b15zdnd11an1n04x5 FILLER_86_1323 ();
 b15zdnd11an1n64x5 FILLER_86_1330 ();
 b15zdnd11an1n64x5 FILLER_86_1394 ();
 b15zdnd11an1n16x5 FILLER_86_1458 ();
 b15zdnd11an1n04x5 FILLER_86_1474 ();
 b15zdnd11an1n08x5 FILLER_86_2265 ();
 b15zdnd00an1n02x5 FILLER_86_2273 ();
 b15zdnd00an1n01x5 FILLER_86_2275 ();
 b15zdnd11an1n64x5 FILLER_87_0 ();
 b15zdnd11an1n64x5 FILLER_87_64 ();
 b15zdnd11an1n64x5 FILLER_87_128 ();
 b15zdnd11an1n64x5 FILLER_87_192 ();
 b15zdnd11an1n64x5 FILLER_87_256 ();
 b15zdnd11an1n64x5 FILLER_87_320 ();
 b15zdnd11an1n16x5 FILLER_87_384 ();
 b15zdnd11an1n08x5 FILLER_87_400 ();
 b15zdnd00an1n01x5 FILLER_87_408 ();
 b15zdnd11an1n64x5 FILLER_87_419 ();
 b15zdnd11an1n64x5 FILLER_87_483 ();
 b15zdnd11an1n64x5 FILLER_87_547 ();
 b15zdnd11an1n64x5 FILLER_87_611 ();
 b15zdnd11an1n64x5 FILLER_87_675 ();
 b15zdnd11an1n64x5 FILLER_87_739 ();
 b15zdnd11an1n64x5 FILLER_87_803 ();
 b15zdnd11an1n64x5 FILLER_87_867 ();
 b15zdnd11an1n64x5 FILLER_87_931 ();
 b15zdnd11an1n64x5 FILLER_87_995 ();
 b15zdnd11an1n64x5 FILLER_87_1059 ();
 b15zdnd11an1n64x5 FILLER_87_1123 ();
 b15zdnd11an1n64x5 FILLER_87_1187 ();
 b15zdnd11an1n32x5 FILLER_87_1251 ();
 b15zdnd11an1n08x5 FILLER_87_1283 ();
 b15zdnd11an1n04x5 FILLER_87_1291 ();
 b15zdnd11an1n04x5 FILLER_87_1298 ();
 b15zdnd11an1n04x5 FILLER_87_1305 ();
 b15zdnd11an1n04x5 FILLER_87_1312 ();
 b15zdnd11an1n32x5 FILLER_87_1319 ();
 b15zdnd11an1n08x5 FILLER_87_1351 ();
 b15zdnd11an1n04x5 FILLER_87_1359 ();
 b15zdnd11an1n64x5 FILLER_87_1371 ();
 b15zdnd11an1n32x5 FILLER_87_1435 ();
 b15zdnd11an1n16x5 FILLER_87_1467 ();
 b15zdnd00an1n02x5 FILLER_87_1483 ();
 b15zdnd00an1n01x5 FILLER_87_1485 ();
 b15zdnd11an1n16x5 FILLER_87_2257 ();
 b15zdnd11an1n08x5 FILLER_87_2273 ();
 b15zdnd00an1n02x5 FILLER_87_2281 ();
 b15zdnd00an1n01x5 FILLER_87_2283 ();
 b15zdnd11an1n64x5 FILLER_88_8 ();
 b15zdnd11an1n64x5 FILLER_88_72 ();
 b15zdnd11an1n64x5 FILLER_88_136 ();
 b15zdnd11an1n64x5 FILLER_88_200 ();
 b15zdnd11an1n64x5 FILLER_88_264 ();
 b15zdnd11an1n64x5 FILLER_88_328 ();
 b15zdnd11an1n64x5 FILLER_88_392 ();
 b15zdnd11an1n64x5 FILLER_88_456 ();
 b15zdnd11an1n64x5 FILLER_88_520 ();
 b15zdnd11an1n32x5 FILLER_88_584 ();
 b15zdnd00an1n02x5 FILLER_88_616 ();
 b15zdnd11an1n64x5 FILLER_88_626 ();
 b15zdnd11an1n16x5 FILLER_88_690 ();
 b15zdnd11an1n08x5 FILLER_88_706 ();
 b15zdnd11an1n04x5 FILLER_88_714 ();
 b15zdnd11an1n64x5 FILLER_88_726 ();
 b15zdnd11an1n64x5 FILLER_88_790 ();
 b15zdnd11an1n64x5 FILLER_88_854 ();
 b15zdnd11an1n64x5 FILLER_88_918 ();
 b15zdnd11an1n32x5 FILLER_88_982 ();
 b15zdnd11an1n16x5 FILLER_88_1014 ();
 b15zdnd11an1n08x5 FILLER_88_1030 ();
 b15zdnd00an1n02x5 FILLER_88_1038 ();
 b15zdnd00an1n01x5 FILLER_88_1040 ();
 b15zdnd11an1n64x5 FILLER_88_1083 ();
 b15zdnd11an1n64x5 FILLER_88_1147 ();
 b15zdnd11an1n64x5 FILLER_88_1211 ();
 b15zdnd11an1n64x5 FILLER_88_1275 ();
 b15zdnd11an1n64x5 FILLER_88_1339 ();
 b15zdnd11an1n64x5 FILLER_88_1403 ();
 b15zdnd11an1n08x5 FILLER_88_1467 ();
 b15zdnd00an1n02x5 FILLER_88_1475 ();
 b15zdnd00an1n01x5 FILLER_88_1477 ();
 b15zdnd11an1n08x5 FILLER_88_2265 ();
 b15zdnd00an1n02x5 FILLER_88_2273 ();
 b15zdnd00an1n01x5 FILLER_88_2275 ();
 b15zdnd11an1n64x5 FILLER_89_0 ();
 b15zdnd11an1n64x5 FILLER_89_64 ();
 b15zdnd11an1n64x5 FILLER_89_128 ();
 b15zdnd11an1n64x5 FILLER_89_192 ();
 b15zdnd11an1n64x5 FILLER_89_256 ();
 b15zdnd11an1n64x5 FILLER_89_320 ();
 b15zdnd11an1n64x5 FILLER_89_384 ();
 b15zdnd11an1n64x5 FILLER_89_448 ();
 b15zdnd11an1n64x5 FILLER_89_512 ();
 b15zdnd11an1n64x5 FILLER_89_576 ();
 b15zdnd11an1n64x5 FILLER_89_640 ();
 b15zdnd11an1n64x5 FILLER_89_704 ();
 b15zdnd11an1n64x5 FILLER_89_768 ();
 b15zdnd11an1n64x5 FILLER_89_832 ();
 b15zdnd11an1n64x5 FILLER_89_896 ();
 b15zdnd11an1n64x5 FILLER_89_960 ();
 b15zdnd11an1n16x5 FILLER_89_1024 ();
 b15zdnd11an1n04x5 FILLER_89_1040 ();
 b15zdnd11an1n64x5 FILLER_89_1052 ();
 b15zdnd11an1n64x5 FILLER_89_1116 ();
 b15zdnd11an1n64x5 FILLER_89_1180 ();
 b15zdnd11an1n64x5 FILLER_89_1244 ();
 b15zdnd11an1n64x5 FILLER_89_1308 ();
 b15zdnd11an1n64x5 FILLER_89_1372 ();
 b15zdnd11an1n32x5 FILLER_89_1436 ();
 b15zdnd11an1n16x5 FILLER_89_1468 ();
 b15zdnd00an1n02x5 FILLER_89_1484 ();
 b15zdnd11an1n16x5 FILLER_89_2257 ();
 b15zdnd11an1n08x5 FILLER_89_2273 ();
 b15zdnd00an1n02x5 FILLER_89_2281 ();
 b15zdnd00an1n01x5 FILLER_89_2283 ();
 b15zdnd11an1n64x5 FILLER_90_8 ();
 b15zdnd11an1n64x5 FILLER_90_72 ();
 b15zdnd11an1n64x5 FILLER_90_136 ();
 b15zdnd11an1n64x5 FILLER_90_200 ();
 b15zdnd11an1n64x5 FILLER_90_264 ();
 b15zdnd11an1n64x5 FILLER_90_328 ();
 b15zdnd11an1n16x5 FILLER_90_392 ();
 b15zdnd11an1n04x5 FILLER_90_408 ();
 b15zdnd00an1n01x5 FILLER_90_412 ();
 b15zdnd11an1n64x5 FILLER_90_425 ();
 b15zdnd11an1n64x5 FILLER_90_489 ();
 b15zdnd11an1n64x5 FILLER_90_553 ();
 b15zdnd11an1n64x5 FILLER_90_617 ();
 b15zdnd11an1n32x5 FILLER_90_681 ();
 b15zdnd11an1n04x5 FILLER_90_713 ();
 b15zdnd00an1n01x5 FILLER_90_717 ();
 b15zdnd11an1n64x5 FILLER_90_726 ();
 b15zdnd11an1n64x5 FILLER_90_790 ();
 b15zdnd11an1n64x5 FILLER_90_854 ();
 b15zdnd11an1n64x5 FILLER_90_918 ();
 b15zdnd11an1n64x5 FILLER_90_982 ();
 b15zdnd11an1n64x5 FILLER_90_1046 ();
 b15zdnd11an1n64x5 FILLER_90_1110 ();
 b15zdnd11an1n64x5 FILLER_90_1174 ();
 b15zdnd11an1n64x5 FILLER_90_1238 ();
 b15zdnd11an1n16x5 FILLER_90_1302 ();
 b15zdnd11an1n04x5 FILLER_90_1318 ();
 b15zdnd00an1n02x5 FILLER_90_1322 ();
 b15zdnd11an1n64x5 FILLER_90_1366 ();
 b15zdnd11an1n32x5 FILLER_90_1430 ();
 b15zdnd11an1n16x5 FILLER_90_1462 ();
 b15zdnd11an1n08x5 FILLER_90_2265 ();
 b15zdnd00an1n02x5 FILLER_90_2273 ();
 b15zdnd00an1n01x5 FILLER_90_2275 ();
 b15zdnd11an1n08x5 FILLER_91_0 ();
 b15zdnd11an1n16x5 FILLER_91_15 ();
 b15zdnd00an1n02x5 FILLER_91_31 ();
 b15zdnd00an1n01x5 FILLER_91_33 ();
 b15zdnd11an1n64x5 FILLER_91_38 ();
 b15zdnd11an1n64x5 FILLER_91_102 ();
 b15zdnd11an1n64x5 FILLER_91_166 ();
 b15zdnd11an1n64x5 FILLER_91_230 ();
 b15zdnd11an1n64x5 FILLER_91_294 ();
 b15zdnd11an1n64x5 FILLER_91_358 ();
 b15zdnd11an1n64x5 FILLER_91_422 ();
 b15zdnd11an1n64x5 FILLER_91_486 ();
 b15zdnd11an1n64x5 FILLER_91_550 ();
 b15zdnd11an1n64x5 FILLER_91_614 ();
 b15zdnd11an1n64x5 FILLER_91_678 ();
 b15zdnd11an1n64x5 FILLER_91_742 ();
 b15zdnd11an1n64x5 FILLER_91_806 ();
 b15zdnd11an1n64x5 FILLER_91_870 ();
 b15zdnd11an1n64x5 FILLER_91_934 ();
 b15zdnd11an1n64x5 FILLER_91_998 ();
 b15zdnd11an1n64x5 FILLER_91_1062 ();
 b15zdnd11an1n64x5 FILLER_91_1126 ();
 b15zdnd11an1n64x5 FILLER_91_1190 ();
 b15zdnd11an1n64x5 FILLER_91_1254 ();
 b15zdnd00an1n01x5 FILLER_91_1318 ();
 b15zdnd11an1n64x5 FILLER_91_1361 ();
 b15zdnd11an1n32x5 FILLER_91_1425 ();
 b15zdnd11an1n16x5 FILLER_91_1457 ();
 b15zdnd11an1n08x5 FILLER_91_1473 ();
 b15zdnd11an1n04x5 FILLER_91_1481 ();
 b15zdnd00an1n01x5 FILLER_91_1485 ();
 b15zdnd11an1n16x5 FILLER_91_2257 ();
 b15zdnd11an1n08x5 FILLER_91_2273 ();
 b15zdnd00an1n02x5 FILLER_91_2281 ();
 b15zdnd00an1n01x5 FILLER_91_2283 ();
 b15zdnd11an1n04x5 FILLER_92_8 ();
 b15zdnd00an1n01x5 FILLER_92_12 ();
 b15zdnd11an1n64x5 FILLER_92_55 ();
 b15zdnd11an1n64x5 FILLER_92_119 ();
 b15zdnd11an1n64x5 FILLER_92_183 ();
 b15zdnd11an1n64x5 FILLER_92_247 ();
 b15zdnd11an1n64x5 FILLER_92_311 ();
 b15zdnd11an1n64x5 FILLER_92_375 ();
 b15zdnd11an1n64x5 FILLER_92_439 ();
 b15zdnd11an1n64x5 FILLER_92_503 ();
 b15zdnd11an1n64x5 FILLER_92_567 ();
 b15zdnd11an1n08x5 FILLER_92_631 ();
 b15zdnd00an1n01x5 FILLER_92_639 ();
 b15zdnd11an1n64x5 FILLER_92_643 ();
 b15zdnd00an1n01x5 FILLER_92_707 ();
 b15zdnd00an1n02x5 FILLER_92_716 ();
 b15zdnd11an1n64x5 FILLER_92_726 ();
 b15zdnd11an1n64x5 FILLER_92_790 ();
 b15zdnd11an1n64x5 FILLER_92_854 ();
 b15zdnd11an1n64x5 FILLER_92_918 ();
 b15zdnd11an1n64x5 FILLER_92_982 ();
 b15zdnd11an1n64x5 FILLER_92_1046 ();
 b15zdnd11an1n64x5 FILLER_92_1110 ();
 b15zdnd11an1n64x5 FILLER_92_1174 ();
 b15zdnd11an1n64x5 FILLER_92_1238 ();
 b15zdnd11an1n64x5 FILLER_92_1302 ();
 b15zdnd11an1n64x5 FILLER_92_1366 ();
 b15zdnd11an1n32x5 FILLER_92_1430 ();
 b15zdnd11an1n16x5 FILLER_92_1462 ();
 b15zdnd11an1n08x5 FILLER_92_2265 ();
 b15zdnd00an1n02x5 FILLER_92_2273 ();
 b15zdnd00an1n01x5 FILLER_92_2275 ();
 b15zdnd11an1n04x5 FILLER_93_0 ();
 b15zdnd00an1n02x5 FILLER_93_4 ();
 b15zdnd00an1n01x5 FILLER_93_6 ();
 b15zdnd11an1n64x5 FILLER_93_49 ();
 b15zdnd11an1n64x5 FILLER_93_113 ();
 b15zdnd11an1n64x5 FILLER_93_177 ();
 b15zdnd11an1n64x5 FILLER_93_241 ();
 b15zdnd11an1n64x5 FILLER_93_305 ();
 b15zdnd11an1n32x5 FILLER_93_369 ();
 b15zdnd00an1n02x5 FILLER_93_401 ();
 b15zdnd11an1n64x5 FILLER_93_419 ();
 b15zdnd11an1n64x5 FILLER_93_483 ();
 b15zdnd11an1n64x5 FILLER_93_547 ();
 b15zdnd11an1n16x5 FILLER_93_611 ();
 b15zdnd11an1n04x5 FILLER_93_627 ();
 b15zdnd11an1n04x5 FILLER_93_634 ();
 b15zdnd11an1n64x5 FILLER_93_680 ();
 b15zdnd11an1n64x5 FILLER_93_744 ();
 b15zdnd11an1n64x5 FILLER_93_808 ();
 b15zdnd11an1n64x5 FILLER_93_872 ();
 b15zdnd11an1n64x5 FILLER_93_936 ();
 b15zdnd11an1n64x5 FILLER_93_1000 ();
 b15zdnd11an1n64x5 FILLER_93_1064 ();
 b15zdnd11an1n64x5 FILLER_93_1128 ();
 b15zdnd11an1n64x5 FILLER_93_1192 ();
 b15zdnd11an1n64x5 FILLER_93_1256 ();
 b15zdnd11an1n64x5 FILLER_93_1320 ();
 b15zdnd11an1n64x5 FILLER_93_1384 ();
 b15zdnd11an1n32x5 FILLER_93_1448 ();
 b15zdnd11an1n04x5 FILLER_93_1480 ();
 b15zdnd00an1n02x5 FILLER_93_1484 ();
 b15zdnd11an1n16x5 FILLER_93_2257 ();
 b15zdnd11an1n08x5 FILLER_93_2273 ();
 b15zdnd00an1n02x5 FILLER_93_2281 ();
 b15zdnd00an1n01x5 FILLER_93_2283 ();
 b15zdnd11an1n08x5 FILLER_94_8 ();
 b15zdnd11an1n04x5 FILLER_94_16 ();
 b15zdnd00an1n02x5 FILLER_94_20 ();
 b15zdnd00an1n01x5 FILLER_94_22 ();
 b15zdnd11an1n08x5 FILLER_94_27 ();
 b15zdnd11an1n04x5 FILLER_94_35 ();
 b15zdnd11an1n64x5 FILLER_94_46 ();
 b15zdnd11an1n64x5 FILLER_94_110 ();
 b15zdnd11an1n64x5 FILLER_94_174 ();
 b15zdnd11an1n64x5 FILLER_94_238 ();
 b15zdnd11an1n64x5 FILLER_94_302 ();
 b15zdnd11an1n64x5 FILLER_94_366 ();
 b15zdnd11an1n64x5 FILLER_94_430 ();
 b15zdnd11an1n64x5 FILLER_94_494 ();
 b15zdnd11an1n32x5 FILLER_94_558 ();
 b15zdnd11an1n16x5 FILLER_94_590 ();
 b15zdnd11an1n08x5 FILLER_94_606 ();
 b15zdnd11an1n04x5 FILLER_94_614 ();
 b15zdnd11an1n04x5 FILLER_94_662 ();
 b15zdnd11an1n32x5 FILLER_94_669 ();
 b15zdnd11an1n16x5 FILLER_94_701 ();
 b15zdnd00an1n01x5 FILLER_94_717 ();
 b15zdnd11an1n64x5 FILLER_94_726 ();
 b15zdnd11an1n64x5 FILLER_94_790 ();
 b15zdnd11an1n64x5 FILLER_94_854 ();
 b15zdnd11an1n64x5 FILLER_94_918 ();
 b15zdnd11an1n64x5 FILLER_94_982 ();
 b15zdnd11an1n64x5 FILLER_94_1046 ();
 b15zdnd11an1n64x5 FILLER_94_1110 ();
 b15zdnd11an1n64x5 FILLER_94_1174 ();
 b15zdnd11an1n64x5 FILLER_94_1238 ();
 b15zdnd11an1n64x5 FILLER_94_1302 ();
 b15zdnd11an1n64x5 FILLER_94_1366 ();
 b15zdnd11an1n32x5 FILLER_94_1430 ();
 b15zdnd11an1n16x5 FILLER_94_1462 ();
 b15zdnd11an1n08x5 FILLER_94_2265 ();
 b15zdnd00an1n02x5 FILLER_94_2273 ();
 b15zdnd00an1n01x5 FILLER_94_2275 ();
 b15zdnd11an1n64x5 FILLER_95_0 ();
 b15zdnd11an1n64x5 FILLER_95_64 ();
 b15zdnd11an1n64x5 FILLER_95_128 ();
 b15zdnd11an1n64x5 FILLER_95_192 ();
 b15zdnd11an1n64x5 FILLER_95_256 ();
 b15zdnd11an1n64x5 FILLER_95_320 ();
 b15zdnd11an1n64x5 FILLER_95_384 ();
 b15zdnd00an1n02x5 FILLER_95_448 ();
 b15zdnd11an1n64x5 FILLER_95_492 ();
 b15zdnd11an1n64x5 FILLER_95_556 ();
 b15zdnd11an1n64x5 FILLER_95_620 ();
 b15zdnd11an1n16x5 FILLER_95_684 ();
 b15zdnd11an1n04x5 FILLER_95_700 ();
 b15zdnd11an1n64x5 FILLER_95_746 ();
 b15zdnd11an1n64x5 FILLER_95_810 ();
 b15zdnd11an1n64x5 FILLER_95_874 ();
 b15zdnd11an1n64x5 FILLER_95_938 ();
 b15zdnd11an1n64x5 FILLER_95_1002 ();
 b15zdnd11an1n64x5 FILLER_95_1066 ();
 b15zdnd11an1n64x5 FILLER_95_1130 ();
 b15zdnd11an1n64x5 FILLER_95_1194 ();
 b15zdnd11an1n64x5 FILLER_95_1258 ();
 b15zdnd11an1n64x5 FILLER_95_1322 ();
 b15zdnd11an1n64x5 FILLER_95_1386 ();
 b15zdnd11an1n32x5 FILLER_95_1450 ();
 b15zdnd11an1n04x5 FILLER_95_1482 ();
 b15zdnd00an1n02x5 FILLER_95_2257 ();
 b15zdnd11an1n16x5 FILLER_95_2262 ();
 b15zdnd11an1n04x5 FILLER_95_2278 ();
 b15zdnd00an1n02x5 FILLER_95_2282 ();
 b15zdnd11an1n64x5 FILLER_96_8 ();
 b15zdnd11an1n64x5 FILLER_96_72 ();
 b15zdnd11an1n64x5 FILLER_96_136 ();
 b15zdnd11an1n64x5 FILLER_96_200 ();
 b15zdnd11an1n64x5 FILLER_96_264 ();
 b15zdnd11an1n32x5 FILLER_96_328 ();
 b15zdnd11an1n16x5 FILLER_96_360 ();
 b15zdnd11an1n08x5 FILLER_96_376 ();
 b15zdnd00an1n01x5 FILLER_96_384 ();
 b15zdnd11an1n64x5 FILLER_96_430 ();
 b15zdnd11an1n64x5 FILLER_96_494 ();
 b15zdnd11an1n64x5 FILLER_96_558 ();
 b15zdnd11an1n32x5 FILLER_96_622 ();
 b15zdnd00an1n02x5 FILLER_96_654 ();
 b15zdnd11an1n16x5 FILLER_96_700 ();
 b15zdnd00an1n02x5 FILLER_96_716 ();
 b15zdnd11an1n64x5 FILLER_96_726 ();
 b15zdnd11an1n64x5 FILLER_96_790 ();
 b15zdnd11an1n64x5 FILLER_96_854 ();
 b15zdnd11an1n64x5 FILLER_96_918 ();
 b15zdnd11an1n64x5 FILLER_96_982 ();
 b15zdnd11an1n64x5 FILLER_96_1046 ();
 b15zdnd11an1n64x5 FILLER_96_1110 ();
 b15zdnd11an1n64x5 FILLER_96_1174 ();
 b15zdnd11an1n64x5 FILLER_96_1238 ();
 b15zdnd11an1n64x5 FILLER_96_1302 ();
 b15zdnd11an1n64x5 FILLER_96_1366 ();
 b15zdnd11an1n32x5 FILLER_96_1430 ();
 b15zdnd11an1n16x5 FILLER_96_1462 ();
 b15zdnd00an1n02x5 FILLER_96_2265 ();
 b15zdnd11an1n04x5 FILLER_96_2270 ();
 b15zdnd00an1n02x5 FILLER_96_2274 ();
 b15zdnd11an1n64x5 FILLER_97_0 ();
 b15zdnd11an1n64x5 FILLER_97_64 ();
 b15zdnd11an1n64x5 FILLER_97_128 ();
 b15zdnd11an1n64x5 FILLER_97_192 ();
 b15zdnd11an1n64x5 FILLER_97_256 ();
 b15zdnd11an1n64x5 FILLER_97_320 ();
 b15zdnd11an1n08x5 FILLER_97_384 ();
 b15zdnd11an1n04x5 FILLER_97_392 ();
 b15zdnd00an1n01x5 FILLER_97_396 ();
 b15zdnd11an1n04x5 FILLER_97_413 ();
 b15zdnd11an1n16x5 FILLER_97_431 ();
 b15zdnd00an1n02x5 FILLER_97_447 ();
 b15zdnd11an1n64x5 FILLER_97_494 ();
 b15zdnd11an1n64x5 FILLER_97_558 ();
 b15zdnd11an1n32x5 FILLER_97_622 ();
 b15zdnd11an1n16x5 FILLER_97_654 ();
 b15zdnd00an1n02x5 FILLER_97_670 ();
 b15zdnd00an1n01x5 FILLER_97_672 ();
 b15zdnd11an1n04x5 FILLER_97_676 ();
 b15zdnd11an1n64x5 FILLER_97_683 ();
 b15zdnd11an1n64x5 FILLER_97_747 ();
 b15zdnd11an1n64x5 FILLER_97_811 ();
 b15zdnd11an1n64x5 FILLER_97_875 ();
 b15zdnd11an1n64x5 FILLER_97_939 ();
 b15zdnd11an1n64x5 FILLER_97_1003 ();
 b15zdnd11an1n64x5 FILLER_97_1067 ();
 b15zdnd11an1n64x5 FILLER_97_1131 ();
 b15zdnd11an1n64x5 FILLER_97_1195 ();
 b15zdnd11an1n64x5 FILLER_97_1259 ();
 b15zdnd11an1n64x5 FILLER_97_1323 ();
 b15zdnd11an1n64x5 FILLER_97_1387 ();
 b15zdnd11an1n32x5 FILLER_97_1451 ();
 b15zdnd00an1n02x5 FILLER_97_1483 ();
 b15zdnd00an1n01x5 FILLER_97_1485 ();
 b15zdnd00an1n02x5 FILLER_97_2257 ();
 b15zdnd11an1n16x5 FILLER_97_2262 ();
 b15zdnd11an1n04x5 FILLER_97_2278 ();
 b15zdnd00an1n02x5 FILLER_97_2282 ();
 b15zdnd11an1n64x5 FILLER_98_8 ();
 b15zdnd11an1n64x5 FILLER_98_72 ();
 b15zdnd11an1n64x5 FILLER_98_136 ();
 b15zdnd11an1n64x5 FILLER_98_200 ();
 b15zdnd11an1n64x5 FILLER_98_264 ();
 b15zdnd11an1n64x5 FILLER_98_328 ();
 b15zdnd11an1n64x5 FILLER_98_392 ();
 b15zdnd11an1n64x5 FILLER_98_456 ();
 b15zdnd11an1n64x5 FILLER_98_520 ();
 b15zdnd11an1n64x5 FILLER_98_584 ();
 b15zdnd11an1n16x5 FILLER_98_648 ();
 b15zdnd11an1n08x5 FILLER_98_664 ();
 b15zdnd11an1n04x5 FILLER_98_672 ();
 b15zdnd00an1n02x5 FILLER_98_676 ();
 b15zdnd00an1n01x5 FILLER_98_678 ();
 b15zdnd11an1n32x5 FILLER_98_682 ();
 b15zdnd11an1n04x5 FILLER_98_714 ();
 b15zdnd11an1n64x5 FILLER_98_726 ();
 b15zdnd11an1n64x5 FILLER_98_790 ();
 b15zdnd11an1n04x5 FILLER_98_854 ();
 b15zdnd11an1n64x5 FILLER_98_885 ();
 b15zdnd11an1n64x5 FILLER_98_949 ();
 b15zdnd11an1n08x5 FILLER_98_1013 ();
 b15zdnd11an1n04x5 FILLER_98_1021 ();
 b15zdnd00an1n01x5 FILLER_98_1025 ();
 b15zdnd11an1n64x5 FILLER_98_1068 ();
 b15zdnd11an1n64x5 FILLER_98_1132 ();
 b15zdnd11an1n32x5 FILLER_98_1196 ();
 b15zdnd11an1n16x5 FILLER_98_1228 ();
 b15zdnd11an1n08x5 FILLER_98_1244 ();
 b15zdnd11an1n04x5 FILLER_98_1252 ();
 b15zdnd00an1n01x5 FILLER_98_1256 ();
 b15zdnd11an1n64x5 FILLER_98_1284 ();
 b15zdnd11an1n64x5 FILLER_98_1348 ();
 b15zdnd11an1n64x5 FILLER_98_1412 ();
 b15zdnd00an1n02x5 FILLER_98_1476 ();
 b15zdnd11an1n08x5 FILLER_98_2265 ();
 b15zdnd00an1n02x5 FILLER_98_2273 ();
 b15zdnd00an1n01x5 FILLER_98_2275 ();
 b15zdnd11an1n64x5 FILLER_99_0 ();
 b15zdnd11an1n64x5 FILLER_99_64 ();
 b15zdnd11an1n64x5 FILLER_99_128 ();
 b15zdnd11an1n64x5 FILLER_99_192 ();
 b15zdnd11an1n64x5 FILLER_99_256 ();
 b15zdnd11an1n32x5 FILLER_99_320 ();
 b15zdnd11an1n16x5 FILLER_99_352 ();
 b15zdnd11an1n04x5 FILLER_99_368 ();
 b15zdnd11an1n64x5 FILLER_99_395 ();
 b15zdnd11an1n16x5 FILLER_99_459 ();
 b15zdnd00an1n01x5 FILLER_99_475 ();
 b15zdnd11an1n64x5 FILLER_99_508 ();
 b15zdnd11an1n16x5 FILLER_99_572 ();
 b15zdnd11an1n08x5 FILLER_99_588 ();
 b15zdnd11an1n64x5 FILLER_99_604 ();
 b15zdnd11an1n64x5 FILLER_99_668 ();
 b15zdnd11an1n64x5 FILLER_99_732 ();
 b15zdnd11an1n32x5 FILLER_99_796 ();
 b15zdnd11an1n16x5 FILLER_99_828 ();
 b15zdnd11an1n08x5 FILLER_99_844 ();
 b15zdnd11an1n04x5 FILLER_99_852 ();
 b15zdnd00an1n02x5 FILLER_99_856 ();
 b15zdnd11an1n64x5 FILLER_99_861 ();
 b15zdnd11an1n64x5 FILLER_99_925 ();
 b15zdnd11an1n64x5 FILLER_99_989 ();
 b15zdnd11an1n64x5 FILLER_99_1053 ();
 b15zdnd11an1n64x5 FILLER_99_1117 ();
 b15zdnd11an1n64x5 FILLER_99_1181 ();
 b15zdnd11an1n08x5 FILLER_99_1245 ();
 b15zdnd11an1n04x5 FILLER_99_1253 ();
 b15zdnd00an1n01x5 FILLER_99_1257 ();
 b15zdnd11an1n64x5 FILLER_99_1261 ();
 b15zdnd11an1n64x5 FILLER_99_1325 ();
 b15zdnd11an1n64x5 FILLER_99_1389 ();
 b15zdnd11an1n32x5 FILLER_99_1453 ();
 b15zdnd00an1n01x5 FILLER_99_1485 ();
 b15zdnd00an1n02x5 FILLER_99_2257 ();
 b15zdnd11an1n16x5 FILLER_99_2262 ();
 b15zdnd11an1n04x5 FILLER_99_2278 ();
 b15zdnd00an1n02x5 FILLER_99_2282 ();
 b15zdnd00an1n02x5 FILLER_100_8 ();
 b15zdnd00an1n01x5 FILLER_100_10 ();
 b15zdnd11an1n08x5 FILLER_100_18 ();
 b15zdnd11an1n04x5 FILLER_100_26 ();
 b15zdnd00an1n01x5 FILLER_100_30 ();
 b15zdnd11an1n64x5 FILLER_100_35 ();
 b15zdnd11an1n32x5 FILLER_100_99 ();
 b15zdnd11an1n04x5 FILLER_100_131 ();
 b15zdnd11an1n64x5 FILLER_100_144 ();
 b15zdnd11an1n64x5 FILLER_100_208 ();
 b15zdnd11an1n64x5 FILLER_100_272 ();
 b15zdnd11an1n32x5 FILLER_100_336 ();
 b15zdnd11an1n08x5 FILLER_100_368 ();
 b15zdnd11an1n04x5 FILLER_100_376 ();
 b15zdnd00an1n01x5 FILLER_100_380 ();
 b15zdnd11an1n64x5 FILLER_100_387 ();
 b15zdnd11an1n08x5 FILLER_100_451 ();
 b15zdnd11an1n04x5 FILLER_100_459 ();
 b15zdnd11an1n64x5 FILLER_100_495 ();
 b15zdnd11an1n64x5 FILLER_100_559 ();
 b15zdnd11an1n64x5 FILLER_100_623 ();
 b15zdnd11an1n16x5 FILLER_100_687 ();
 b15zdnd11an1n08x5 FILLER_100_703 ();
 b15zdnd11an1n04x5 FILLER_100_711 ();
 b15zdnd00an1n02x5 FILLER_100_715 ();
 b15zdnd00an1n01x5 FILLER_100_717 ();
 b15zdnd11an1n64x5 FILLER_100_726 ();
 b15zdnd11an1n64x5 FILLER_100_790 ();
 b15zdnd11an1n64x5 FILLER_100_854 ();
 b15zdnd11an1n64x5 FILLER_100_918 ();
 b15zdnd11an1n64x5 FILLER_100_982 ();
 b15zdnd11an1n64x5 FILLER_100_1046 ();
 b15zdnd11an1n64x5 FILLER_100_1110 ();
 b15zdnd11an1n64x5 FILLER_100_1174 ();
 b15zdnd11an1n64x5 FILLER_100_1238 ();
 b15zdnd11an1n64x5 FILLER_100_1302 ();
 b15zdnd11an1n64x5 FILLER_100_1366 ();
 b15zdnd11an1n32x5 FILLER_100_1430 ();
 b15zdnd11an1n16x5 FILLER_100_1462 ();
 b15zdnd11an1n08x5 FILLER_100_2265 ();
 b15zdnd00an1n02x5 FILLER_100_2273 ();
 b15zdnd00an1n01x5 FILLER_100_2275 ();
 b15zdnd11an1n08x5 FILLER_101_0 ();
 b15zdnd00an1n02x5 FILLER_101_8 ();
 b15zdnd00an1n01x5 FILLER_101_10 ();
 b15zdnd11an1n64x5 FILLER_101_53 ();
 b15zdnd11an1n64x5 FILLER_101_117 ();
 b15zdnd11an1n64x5 FILLER_101_181 ();
 b15zdnd11an1n64x5 FILLER_101_245 ();
 b15zdnd11an1n64x5 FILLER_101_309 ();
 b15zdnd11an1n64x5 FILLER_101_373 ();
 b15zdnd11an1n64x5 FILLER_101_437 ();
 b15zdnd11an1n64x5 FILLER_101_501 ();
 b15zdnd11an1n64x5 FILLER_101_565 ();
 b15zdnd11an1n64x5 FILLER_101_629 ();
 b15zdnd11an1n64x5 FILLER_101_693 ();
 b15zdnd11an1n64x5 FILLER_101_757 ();
 b15zdnd11an1n64x5 FILLER_101_821 ();
 b15zdnd11an1n64x5 FILLER_101_885 ();
 b15zdnd11an1n64x5 FILLER_101_949 ();
 b15zdnd11an1n64x5 FILLER_101_1013 ();
 b15zdnd11an1n64x5 FILLER_101_1077 ();
 b15zdnd11an1n64x5 FILLER_101_1141 ();
 b15zdnd11an1n64x5 FILLER_101_1205 ();
 b15zdnd11an1n64x5 FILLER_101_1269 ();
 b15zdnd11an1n64x5 FILLER_101_1333 ();
 b15zdnd11an1n64x5 FILLER_101_1397 ();
 b15zdnd11an1n16x5 FILLER_101_1461 ();
 b15zdnd11an1n08x5 FILLER_101_1477 ();
 b15zdnd00an1n01x5 FILLER_101_1485 ();
 b15zdnd00an1n02x5 FILLER_101_2257 ();
 b15zdnd11an1n16x5 FILLER_101_2262 ();
 b15zdnd11an1n04x5 FILLER_101_2278 ();
 b15zdnd00an1n02x5 FILLER_101_2282 ();
 b15zdnd00an1n02x5 FILLER_102_8 ();
 b15zdnd11an1n64x5 FILLER_102_52 ();
 b15zdnd11an1n64x5 FILLER_102_116 ();
 b15zdnd11an1n64x5 FILLER_102_180 ();
 b15zdnd11an1n64x5 FILLER_102_244 ();
 b15zdnd11an1n64x5 FILLER_102_308 ();
 b15zdnd11an1n64x5 FILLER_102_372 ();
 b15zdnd11an1n64x5 FILLER_102_436 ();
 b15zdnd11an1n64x5 FILLER_102_500 ();
 b15zdnd11an1n64x5 FILLER_102_564 ();
 b15zdnd11an1n64x5 FILLER_102_628 ();
 b15zdnd11an1n16x5 FILLER_102_692 ();
 b15zdnd11an1n08x5 FILLER_102_708 ();
 b15zdnd00an1n02x5 FILLER_102_716 ();
 b15zdnd11an1n64x5 FILLER_102_726 ();
 b15zdnd11an1n64x5 FILLER_102_790 ();
 b15zdnd11an1n64x5 FILLER_102_854 ();
 b15zdnd11an1n64x5 FILLER_102_918 ();
 b15zdnd11an1n64x5 FILLER_102_982 ();
 b15zdnd11an1n64x5 FILLER_102_1046 ();
 b15zdnd11an1n64x5 FILLER_102_1110 ();
 b15zdnd11an1n64x5 FILLER_102_1174 ();
 b15zdnd11an1n64x5 FILLER_102_1238 ();
 b15zdnd11an1n64x5 FILLER_102_1302 ();
 b15zdnd11an1n64x5 FILLER_102_1366 ();
 b15zdnd11an1n32x5 FILLER_102_1430 ();
 b15zdnd11an1n16x5 FILLER_102_1462 ();
 b15zdnd00an1n02x5 FILLER_102_2265 ();
 b15zdnd00an1n01x5 FILLER_102_2267 ();
 b15zdnd11an1n04x5 FILLER_102_2271 ();
 b15zdnd00an1n01x5 FILLER_102_2275 ();
 b15zdnd11an1n16x5 FILLER_103_0 ();
 b15zdnd00an1n02x5 FILLER_103_16 ();
 b15zdnd00an1n01x5 FILLER_103_18 ();
 b15zdnd11an1n04x5 FILLER_103_23 ();
 b15zdnd00an1n02x5 FILLER_103_27 ();
 b15zdnd11an1n64x5 FILLER_103_36 ();
 b15zdnd11an1n64x5 FILLER_103_100 ();
 b15zdnd11an1n64x5 FILLER_103_164 ();
 b15zdnd11an1n64x5 FILLER_103_228 ();
 b15zdnd11an1n64x5 FILLER_103_292 ();
 b15zdnd11an1n64x5 FILLER_103_356 ();
 b15zdnd11an1n64x5 FILLER_103_420 ();
 b15zdnd11an1n64x5 FILLER_103_484 ();
 b15zdnd11an1n64x5 FILLER_103_548 ();
 b15zdnd11an1n64x5 FILLER_103_612 ();
 b15zdnd11an1n64x5 FILLER_103_676 ();
 b15zdnd11an1n64x5 FILLER_103_740 ();
 b15zdnd11an1n64x5 FILLER_103_804 ();
 b15zdnd11an1n64x5 FILLER_103_868 ();
 b15zdnd11an1n64x5 FILLER_103_932 ();
 b15zdnd11an1n64x5 FILLER_103_996 ();
 b15zdnd11an1n64x5 FILLER_103_1060 ();
 b15zdnd11an1n64x5 FILLER_103_1124 ();
 b15zdnd11an1n64x5 FILLER_103_1188 ();
 b15zdnd11an1n64x5 FILLER_103_1252 ();
 b15zdnd11an1n64x5 FILLER_103_1316 ();
 b15zdnd11an1n64x5 FILLER_103_1380 ();
 b15zdnd11an1n32x5 FILLER_103_1444 ();
 b15zdnd11an1n04x5 FILLER_103_1476 ();
 b15zdnd00an1n01x5 FILLER_103_1480 ();
 b15zdnd00an1n02x5 FILLER_103_1484 ();
 b15zdnd00an1n02x5 FILLER_103_2257 ();
 b15zdnd11an1n16x5 FILLER_103_2262 ();
 b15zdnd11an1n04x5 FILLER_103_2278 ();
 b15zdnd00an1n02x5 FILLER_103_2282 ();
 b15zdnd11an1n64x5 FILLER_104_8 ();
 b15zdnd11an1n64x5 FILLER_104_72 ();
 b15zdnd11an1n64x5 FILLER_104_136 ();
 b15zdnd11an1n64x5 FILLER_104_200 ();
 b15zdnd11an1n64x5 FILLER_104_264 ();
 b15zdnd11an1n64x5 FILLER_104_328 ();
 b15zdnd11an1n64x5 FILLER_104_392 ();
 b15zdnd11an1n64x5 FILLER_104_456 ();
 b15zdnd11an1n64x5 FILLER_104_520 ();
 b15zdnd11an1n64x5 FILLER_104_584 ();
 b15zdnd11an1n64x5 FILLER_104_648 ();
 b15zdnd11an1n04x5 FILLER_104_712 ();
 b15zdnd00an1n02x5 FILLER_104_716 ();
 b15zdnd11an1n64x5 FILLER_104_726 ();
 b15zdnd11an1n64x5 FILLER_104_790 ();
 b15zdnd11an1n64x5 FILLER_104_854 ();
 b15zdnd11an1n64x5 FILLER_104_918 ();
 b15zdnd11an1n64x5 FILLER_104_982 ();
 b15zdnd11an1n64x5 FILLER_104_1046 ();
 b15zdnd11an1n64x5 FILLER_104_1110 ();
 b15zdnd11an1n64x5 FILLER_104_1174 ();
 b15zdnd11an1n64x5 FILLER_104_1238 ();
 b15zdnd11an1n64x5 FILLER_104_1302 ();
 b15zdnd11an1n64x5 FILLER_104_1366 ();
 b15zdnd11an1n32x5 FILLER_104_1430 ();
 b15zdnd11an1n16x5 FILLER_104_1462 ();
 b15zdnd11an1n08x5 FILLER_104_2265 ();
 b15zdnd00an1n02x5 FILLER_104_2273 ();
 b15zdnd00an1n01x5 FILLER_104_2275 ();
 b15zdnd11an1n64x5 FILLER_105_0 ();
 b15zdnd11an1n64x5 FILLER_105_64 ();
 b15zdnd11an1n64x5 FILLER_105_128 ();
 b15zdnd11an1n64x5 FILLER_105_192 ();
 b15zdnd11an1n64x5 FILLER_105_256 ();
 b15zdnd11an1n64x5 FILLER_105_320 ();
 b15zdnd11an1n64x5 FILLER_105_384 ();
 b15zdnd11an1n64x5 FILLER_105_448 ();
 b15zdnd11an1n64x5 FILLER_105_512 ();
 b15zdnd11an1n64x5 FILLER_105_576 ();
 b15zdnd11an1n64x5 FILLER_105_640 ();
 b15zdnd11an1n64x5 FILLER_105_704 ();
 b15zdnd11an1n64x5 FILLER_105_768 ();
 b15zdnd11an1n64x5 FILLER_105_832 ();
 b15zdnd11an1n64x5 FILLER_105_896 ();
 b15zdnd11an1n64x5 FILLER_105_960 ();
 b15zdnd11an1n32x5 FILLER_105_1024 ();
 b15zdnd11an1n16x5 FILLER_105_1056 ();
 b15zdnd11an1n04x5 FILLER_105_1072 ();
 b15zdnd00an1n01x5 FILLER_105_1076 ();
 b15zdnd11an1n64x5 FILLER_105_1085 ();
 b15zdnd11an1n64x5 FILLER_105_1149 ();
 b15zdnd11an1n64x5 FILLER_105_1213 ();
 b15zdnd11an1n64x5 FILLER_105_1277 ();
 b15zdnd11an1n64x5 FILLER_105_1341 ();
 b15zdnd11an1n64x5 FILLER_105_1405 ();
 b15zdnd00an1n01x5 FILLER_105_1469 ();
 b15zdnd11an1n08x5 FILLER_105_1473 ();
 b15zdnd00an1n02x5 FILLER_105_1484 ();
 b15zdnd11an1n08x5 FILLER_105_2257 ();
 b15zdnd11an1n04x5 FILLER_105_2265 ();
 b15zdnd00an1n02x5 FILLER_105_2269 ();
 b15zdnd00an1n01x5 FILLER_105_2271 ();
 b15zdnd11an1n04x5 FILLER_105_2280 ();
 b15zdnd11an1n64x5 FILLER_106_8 ();
 b15zdnd11an1n64x5 FILLER_106_72 ();
 b15zdnd11an1n64x5 FILLER_106_136 ();
 b15zdnd11an1n64x5 FILLER_106_200 ();
 b15zdnd11an1n64x5 FILLER_106_264 ();
 b15zdnd11an1n64x5 FILLER_106_328 ();
 b15zdnd11an1n64x5 FILLER_106_392 ();
 b15zdnd11an1n64x5 FILLER_106_456 ();
 b15zdnd11an1n64x5 FILLER_106_520 ();
 b15zdnd11an1n64x5 FILLER_106_584 ();
 b15zdnd11an1n64x5 FILLER_106_648 ();
 b15zdnd11an1n04x5 FILLER_106_712 ();
 b15zdnd00an1n02x5 FILLER_106_716 ();
 b15zdnd11an1n64x5 FILLER_106_726 ();
 b15zdnd11an1n64x5 FILLER_106_790 ();
 b15zdnd11an1n64x5 FILLER_106_854 ();
 b15zdnd11an1n64x5 FILLER_106_918 ();
 b15zdnd11an1n64x5 FILLER_106_982 ();
 b15zdnd11an1n64x5 FILLER_106_1046 ();
 b15zdnd11an1n64x5 FILLER_106_1110 ();
 b15zdnd11an1n64x5 FILLER_106_1174 ();
 b15zdnd11an1n64x5 FILLER_106_1238 ();
 b15zdnd11an1n64x5 FILLER_106_1302 ();
 b15zdnd11an1n64x5 FILLER_106_1366 ();
 b15zdnd11an1n32x5 FILLER_106_1430 ();
 b15zdnd11an1n16x5 FILLER_106_1462 ();
 b15zdnd11an1n08x5 FILLER_106_2265 ();
 b15zdnd00an1n02x5 FILLER_106_2273 ();
 b15zdnd00an1n01x5 FILLER_106_2275 ();
 b15zdnd11an1n64x5 FILLER_107_0 ();
 b15zdnd11an1n64x5 FILLER_107_64 ();
 b15zdnd11an1n08x5 FILLER_107_128 ();
 b15zdnd00an1n02x5 FILLER_107_136 ();
 b15zdnd11an1n64x5 FILLER_107_143 ();
 b15zdnd11an1n32x5 FILLER_107_207 ();
 b15zdnd11an1n64x5 FILLER_107_281 ();
 b15zdnd11an1n64x5 FILLER_107_345 ();
 b15zdnd11an1n32x5 FILLER_107_409 ();
 b15zdnd11an1n04x5 FILLER_107_441 ();
 b15zdnd00an1n02x5 FILLER_107_445 ();
 b15zdnd00an1n01x5 FILLER_107_447 ();
 b15zdnd11an1n64x5 FILLER_107_464 ();
 b15zdnd11an1n64x5 FILLER_107_528 ();
 b15zdnd11an1n64x5 FILLER_107_592 ();
 b15zdnd11an1n64x5 FILLER_107_656 ();
 b15zdnd11an1n64x5 FILLER_107_720 ();
 b15zdnd11an1n64x5 FILLER_107_784 ();
 b15zdnd11an1n64x5 FILLER_107_848 ();
 b15zdnd11an1n64x5 FILLER_107_912 ();
 b15zdnd11an1n64x5 FILLER_107_976 ();
 b15zdnd11an1n64x5 FILLER_107_1040 ();
 b15zdnd11an1n64x5 FILLER_107_1104 ();
 b15zdnd11an1n64x5 FILLER_107_1168 ();
 b15zdnd11an1n64x5 FILLER_107_1232 ();
 b15zdnd11an1n64x5 FILLER_107_1296 ();
 b15zdnd11an1n64x5 FILLER_107_1360 ();
 b15zdnd11an1n32x5 FILLER_107_1424 ();
 b15zdnd11an1n16x5 FILLER_107_1456 ();
 b15zdnd11an1n08x5 FILLER_107_1472 ();
 b15zdnd00an1n01x5 FILLER_107_1480 ();
 b15zdnd00an1n02x5 FILLER_107_1484 ();
 b15zdnd11an1n16x5 FILLER_107_2257 ();
 b15zdnd00an1n01x5 FILLER_107_2273 ();
 b15zdnd00an1n02x5 FILLER_107_2282 ();
 b15zdnd11an1n64x5 FILLER_108_8 ();
 b15zdnd11an1n64x5 FILLER_108_72 ();
 b15zdnd11an1n64x5 FILLER_108_136 ();
 b15zdnd11an1n32x5 FILLER_108_200 ();
 b15zdnd11an1n08x5 FILLER_108_232 ();
 b15zdnd00an1n02x5 FILLER_108_240 ();
 b15zdnd00an1n01x5 FILLER_108_242 ();
 b15zdnd11an1n64x5 FILLER_108_285 ();
 b15zdnd11an1n64x5 FILLER_108_349 ();
 b15zdnd11an1n64x5 FILLER_108_413 ();
 b15zdnd11an1n64x5 FILLER_108_477 ();
 b15zdnd11an1n64x5 FILLER_108_541 ();
 b15zdnd11an1n64x5 FILLER_108_605 ();
 b15zdnd11an1n32x5 FILLER_108_669 ();
 b15zdnd11an1n16x5 FILLER_108_701 ();
 b15zdnd00an1n01x5 FILLER_108_717 ();
 b15zdnd11an1n64x5 FILLER_108_726 ();
 b15zdnd11an1n64x5 FILLER_108_790 ();
 b15zdnd11an1n64x5 FILLER_108_854 ();
 b15zdnd11an1n64x5 FILLER_108_918 ();
 b15zdnd11an1n64x5 FILLER_108_982 ();
 b15zdnd11an1n64x5 FILLER_108_1046 ();
 b15zdnd11an1n64x5 FILLER_108_1110 ();
 b15zdnd11an1n64x5 FILLER_108_1174 ();
 b15zdnd11an1n64x5 FILLER_108_1238 ();
 b15zdnd11an1n16x5 FILLER_108_1302 ();
 b15zdnd11an1n08x5 FILLER_108_1318 ();
 b15zdnd11an1n64x5 FILLER_108_1334 ();
 b15zdnd11an1n64x5 FILLER_108_1398 ();
 b15zdnd11an1n16x5 FILLER_108_1462 ();
 b15zdnd11an1n08x5 FILLER_108_2265 ();
 b15zdnd00an1n02x5 FILLER_108_2273 ();
 b15zdnd00an1n01x5 FILLER_108_2275 ();
 b15zdnd11an1n64x5 FILLER_109_0 ();
 b15zdnd11an1n64x5 FILLER_109_64 ();
 b15zdnd11an1n64x5 FILLER_109_128 ();
 b15zdnd11an1n64x5 FILLER_109_192 ();
 b15zdnd11an1n64x5 FILLER_109_256 ();
 b15zdnd11an1n64x5 FILLER_109_320 ();
 b15zdnd11an1n64x5 FILLER_109_384 ();
 b15zdnd11an1n64x5 FILLER_109_448 ();
 b15zdnd11an1n64x5 FILLER_109_512 ();
 b15zdnd11an1n64x5 FILLER_109_576 ();
 b15zdnd11an1n64x5 FILLER_109_640 ();
 b15zdnd11an1n64x5 FILLER_109_704 ();
 b15zdnd11an1n64x5 FILLER_109_768 ();
 b15zdnd11an1n64x5 FILLER_109_832 ();
 b15zdnd11an1n64x5 FILLER_109_896 ();
 b15zdnd11an1n64x5 FILLER_109_960 ();
 b15zdnd11an1n64x5 FILLER_109_1024 ();
 b15zdnd11an1n64x5 FILLER_109_1088 ();
 b15zdnd11an1n64x5 FILLER_109_1152 ();
 b15zdnd11an1n64x5 FILLER_109_1216 ();
 b15zdnd11an1n64x5 FILLER_109_1280 ();
 b15zdnd11an1n64x5 FILLER_109_1344 ();
 b15zdnd11an1n64x5 FILLER_109_1408 ();
 b15zdnd11an1n08x5 FILLER_109_1472 ();
 b15zdnd11an1n04x5 FILLER_109_1480 ();
 b15zdnd00an1n02x5 FILLER_109_1484 ();
 b15zdnd11an1n16x5 FILLER_109_2257 ();
 b15zdnd11an1n08x5 FILLER_109_2273 ();
 b15zdnd00an1n02x5 FILLER_109_2281 ();
 b15zdnd00an1n01x5 FILLER_109_2283 ();
 b15zdnd11an1n64x5 FILLER_110_8 ();
 b15zdnd11an1n64x5 FILLER_110_72 ();
 b15zdnd11an1n64x5 FILLER_110_136 ();
 b15zdnd11an1n64x5 FILLER_110_200 ();
 b15zdnd11an1n64x5 FILLER_110_264 ();
 b15zdnd11an1n64x5 FILLER_110_328 ();
 b15zdnd11an1n64x5 FILLER_110_392 ();
 b15zdnd11an1n64x5 FILLER_110_456 ();
 b15zdnd11an1n64x5 FILLER_110_520 ();
 b15zdnd11an1n64x5 FILLER_110_584 ();
 b15zdnd11an1n64x5 FILLER_110_648 ();
 b15zdnd11an1n04x5 FILLER_110_712 ();
 b15zdnd00an1n02x5 FILLER_110_716 ();
 b15zdnd11an1n64x5 FILLER_110_726 ();
 b15zdnd11an1n64x5 FILLER_110_790 ();
 b15zdnd11an1n64x5 FILLER_110_854 ();
 b15zdnd11an1n64x5 FILLER_110_918 ();
 b15zdnd11an1n64x5 FILLER_110_982 ();
 b15zdnd11an1n64x5 FILLER_110_1046 ();
 b15zdnd11an1n64x5 FILLER_110_1110 ();
 b15zdnd11an1n64x5 FILLER_110_1174 ();
 b15zdnd11an1n64x5 FILLER_110_1238 ();
 b15zdnd11an1n64x5 FILLER_110_1302 ();
 b15zdnd11an1n64x5 FILLER_110_1366 ();
 b15zdnd11an1n32x5 FILLER_110_1430 ();
 b15zdnd11an1n16x5 FILLER_110_1462 ();
 b15zdnd00an1n02x5 FILLER_110_2265 ();
 b15zdnd00an1n02x5 FILLER_110_2274 ();
 b15zdnd11an1n64x5 FILLER_111_0 ();
 b15zdnd11an1n64x5 FILLER_111_64 ();
 b15zdnd11an1n64x5 FILLER_111_128 ();
 b15zdnd11an1n32x5 FILLER_111_192 ();
 b15zdnd11an1n08x5 FILLER_111_224 ();
 b15zdnd11an1n04x5 FILLER_111_232 ();
 b15zdnd11an1n64x5 FILLER_111_278 ();
 b15zdnd11an1n64x5 FILLER_111_342 ();
 b15zdnd11an1n64x5 FILLER_111_406 ();
 b15zdnd11an1n64x5 FILLER_111_470 ();
 b15zdnd11an1n64x5 FILLER_111_534 ();
 b15zdnd11an1n64x5 FILLER_111_598 ();
 b15zdnd11an1n64x5 FILLER_111_662 ();
 b15zdnd11an1n64x5 FILLER_111_726 ();
 b15zdnd11an1n64x5 FILLER_111_790 ();
 b15zdnd11an1n64x5 FILLER_111_854 ();
 b15zdnd11an1n64x5 FILLER_111_918 ();
 b15zdnd11an1n04x5 FILLER_111_982 ();
 b15zdnd00an1n02x5 FILLER_111_986 ();
 b15zdnd11an1n64x5 FILLER_111_997 ();
 b15zdnd11an1n64x5 FILLER_111_1061 ();
 b15zdnd11an1n64x5 FILLER_111_1125 ();
 b15zdnd11an1n64x5 FILLER_111_1189 ();
 b15zdnd11an1n64x5 FILLER_111_1253 ();
 b15zdnd11an1n64x5 FILLER_111_1317 ();
 b15zdnd11an1n64x5 FILLER_111_1381 ();
 b15zdnd11an1n32x5 FILLER_111_1445 ();
 b15zdnd11an1n08x5 FILLER_111_1477 ();
 b15zdnd00an1n01x5 FILLER_111_1485 ();
 b15zdnd11an1n08x5 FILLER_111_2257 ();
 b15zdnd11an1n04x5 FILLER_111_2265 ();
 b15zdnd00an1n02x5 FILLER_111_2269 ();
 b15zdnd00an1n01x5 FILLER_111_2271 ();
 b15zdnd11an1n04x5 FILLER_111_2279 ();
 b15zdnd00an1n01x5 FILLER_111_2283 ();
 b15zdnd11an1n64x5 FILLER_112_8 ();
 b15zdnd11an1n64x5 FILLER_112_72 ();
 b15zdnd11an1n64x5 FILLER_112_136 ();
 b15zdnd11an1n64x5 FILLER_112_200 ();
 b15zdnd11an1n64x5 FILLER_112_264 ();
 b15zdnd11an1n64x5 FILLER_112_328 ();
 b15zdnd11an1n64x5 FILLER_112_392 ();
 b15zdnd11an1n64x5 FILLER_112_456 ();
 b15zdnd11an1n64x5 FILLER_112_520 ();
 b15zdnd11an1n64x5 FILLER_112_584 ();
 b15zdnd11an1n64x5 FILLER_112_648 ();
 b15zdnd11an1n04x5 FILLER_112_712 ();
 b15zdnd00an1n02x5 FILLER_112_716 ();
 b15zdnd11an1n64x5 FILLER_112_726 ();
 b15zdnd11an1n64x5 FILLER_112_790 ();
 b15zdnd11an1n64x5 FILLER_112_854 ();
 b15zdnd11an1n64x5 FILLER_112_918 ();
 b15zdnd11an1n64x5 FILLER_112_982 ();
 b15zdnd11an1n64x5 FILLER_112_1046 ();
 b15zdnd11an1n64x5 FILLER_112_1110 ();
 b15zdnd11an1n64x5 FILLER_112_1174 ();
 b15zdnd11an1n64x5 FILLER_112_1238 ();
 b15zdnd11an1n16x5 FILLER_112_1302 ();
 b15zdnd11an1n64x5 FILLER_112_1326 ();
 b15zdnd11an1n64x5 FILLER_112_1390 ();
 b15zdnd11an1n16x5 FILLER_112_1454 ();
 b15zdnd11an1n08x5 FILLER_112_1470 ();
 b15zdnd11an1n08x5 FILLER_112_2265 ();
 b15zdnd00an1n02x5 FILLER_112_2273 ();
 b15zdnd00an1n01x5 FILLER_112_2275 ();
 b15zdnd11an1n64x5 FILLER_113_0 ();
 b15zdnd11an1n64x5 FILLER_113_64 ();
 b15zdnd11an1n64x5 FILLER_113_128 ();
 b15zdnd11an1n64x5 FILLER_113_192 ();
 b15zdnd11an1n64x5 FILLER_113_256 ();
 b15zdnd11an1n64x5 FILLER_113_320 ();
 b15zdnd11an1n08x5 FILLER_113_384 ();
 b15zdnd11an1n04x5 FILLER_113_392 ();
 b15zdnd00an1n02x5 FILLER_113_396 ();
 b15zdnd00an1n01x5 FILLER_113_398 ();
 b15zdnd11an1n64x5 FILLER_113_427 ();
 b15zdnd11an1n64x5 FILLER_113_491 ();
 b15zdnd11an1n64x5 FILLER_113_555 ();
 b15zdnd11an1n64x5 FILLER_113_619 ();
 b15zdnd11an1n64x5 FILLER_113_683 ();
 b15zdnd11an1n64x5 FILLER_113_747 ();
 b15zdnd11an1n64x5 FILLER_113_811 ();
 b15zdnd11an1n64x5 FILLER_113_875 ();
 b15zdnd11an1n64x5 FILLER_113_939 ();
 b15zdnd11an1n64x5 FILLER_113_1003 ();
 b15zdnd11an1n64x5 FILLER_113_1067 ();
 b15zdnd11an1n64x5 FILLER_113_1131 ();
 b15zdnd11an1n64x5 FILLER_113_1195 ();
 b15zdnd11an1n64x5 FILLER_113_1259 ();
 b15zdnd11an1n64x5 FILLER_113_1323 ();
 b15zdnd11an1n64x5 FILLER_113_1387 ();
 b15zdnd11an1n32x5 FILLER_113_1451 ();
 b15zdnd00an1n02x5 FILLER_113_1483 ();
 b15zdnd00an1n01x5 FILLER_113_1485 ();
 b15zdnd11an1n16x5 FILLER_113_2257 ();
 b15zdnd11an1n08x5 FILLER_113_2273 ();
 b15zdnd00an1n02x5 FILLER_113_2281 ();
 b15zdnd00an1n01x5 FILLER_113_2283 ();
 b15zdnd11an1n64x5 FILLER_114_8 ();
 b15zdnd11an1n64x5 FILLER_114_72 ();
 b15zdnd11an1n64x5 FILLER_114_136 ();
 b15zdnd11an1n32x5 FILLER_114_200 ();
 b15zdnd00an1n02x5 FILLER_114_232 ();
 b15zdnd11an1n64x5 FILLER_114_276 ();
 b15zdnd11an1n64x5 FILLER_114_340 ();
 b15zdnd11an1n64x5 FILLER_114_404 ();
 b15zdnd11an1n64x5 FILLER_114_468 ();
 b15zdnd11an1n64x5 FILLER_114_532 ();
 b15zdnd11an1n64x5 FILLER_114_596 ();
 b15zdnd11an1n32x5 FILLER_114_660 ();
 b15zdnd11an1n16x5 FILLER_114_692 ();
 b15zdnd11an1n08x5 FILLER_114_708 ();
 b15zdnd00an1n02x5 FILLER_114_716 ();
 b15zdnd11an1n64x5 FILLER_114_726 ();
 b15zdnd11an1n64x5 FILLER_114_790 ();
 b15zdnd11an1n64x5 FILLER_114_854 ();
 b15zdnd11an1n64x5 FILLER_114_918 ();
 b15zdnd11an1n64x5 FILLER_114_982 ();
 b15zdnd11an1n64x5 FILLER_114_1046 ();
 b15zdnd11an1n64x5 FILLER_114_1110 ();
 b15zdnd11an1n64x5 FILLER_114_1174 ();
 b15zdnd11an1n64x5 FILLER_114_1238 ();
 b15zdnd11an1n64x5 FILLER_114_1302 ();
 b15zdnd11an1n64x5 FILLER_114_1366 ();
 b15zdnd11an1n32x5 FILLER_114_1430 ();
 b15zdnd11an1n16x5 FILLER_114_1462 ();
 b15zdnd11an1n08x5 FILLER_114_2265 ();
 b15zdnd00an1n02x5 FILLER_114_2273 ();
 b15zdnd00an1n01x5 FILLER_114_2275 ();
 b15zdnd11an1n64x5 FILLER_115_0 ();
 b15zdnd11an1n64x5 FILLER_115_64 ();
 b15zdnd11an1n64x5 FILLER_115_128 ();
 b15zdnd11an1n64x5 FILLER_115_192 ();
 b15zdnd11an1n64x5 FILLER_115_256 ();
 b15zdnd11an1n64x5 FILLER_115_320 ();
 b15zdnd11an1n64x5 FILLER_115_384 ();
 b15zdnd11an1n64x5 FILLER_115_448 ();
 b15zdnd11an1n64x5 FILLER_115_512 ();
 b15zdnd11an1n64x5 FILLER_115_576 ();
 b15zdnd11an1n64x5 FILLER_115_640 ();
 b15zdnd11an1n64x5 FILLER_115_704 ();
 b15zdnd11an1n64x5 FILLER_115_768 ();
 b15zdnd11an1n64x5 FILLER_115_832 ();
 b15zdnd11an1n64x5 FILLER_115_896 ();
 b15zdnd11an1n64x5 FILLER_115_960 ();
 b15zdnd11an1n64x5 FILLER_115_1024 ();
 b15zdnd11an1n64x5 FILLER_115_1088 ();
 b15zdnd11an1n64x5 FILLER_115_1152 ();
 b15zdnd11an1n64x5 FILLER_115_1216 ();
 b15zdnd11an1n64x5 FILLER_115_1280 ();
 b15zdnd11an1n64x5 FILLER_115_1344 ();
 b15zdnd11an1n64x5 FILLER_115_1408 ();
 b15zdnd11an1n08x5 FILLER_115_1472 ();
 b15zdnd11an1n04x5 FILLER_115_1480 ();
 b15zdnd00an1n02x5 FILLER_115_1484 ();
 b15zdnd11an1n16x5 FILLER_115_2257 ();
 b15zdnd11an1n08x5 FILLER_115_2273 ();
 b15zdnd00an1n02x5 FILLER_115_2281 ();
 b15zdnd00an1n01x5 FILLER_115_2283 ();
 b15zdnd11an1n64x5 FILLER_116_8 ();
 b15zdnd11an1n64x5 FILLER_116_72 ();
 b15zdnd11an1n64x5 FILLER_116_136 ();
 b15zdnd11an1n64x5 FILLER_116_200 ();
 b15zdnd11an1n64x5 FILLER_116_264 ();
 b15zdnd11an1n64x5 FILLER_116_328 ();
 b15zdnd11an1n64x5 FILLER_116_392 ();
 b15zdnd11an1n64x5 FILLER_116_456 ();
 b15zdnd11an1n64x5 FILLER_116_520 ();
 b15zdnd11an1n64x5 FILLER_116_584 ();
 b15zdnd11an1n64x5 FILLER_116_648 ();
 b15zdnd11an1n04x5 FILLER_116_712 ();
 b15zdnd00an1n02x5 FILLER_116_716 ();
 b15zdnd11an1n64x5 FILLER_116_726 ();
 b15zdnd11an1n64x5 FILLER_116_790 ();
 b15zdnd11an1n64x5 FILLER_116_854 ();
 b15zdnd11an1n64x5 FILLER_116_918 ();
 b15zdnd11an1n64x5 FILLER_116_982 ();
 b15zdnd11an1n64x5 FILLER_116_1046 ();
 b15zdnd11an1n64x5 FILLER_116_1110 ();
 b15zdnd11an1n64x5 FILLER_116_1174 ();
 b15zdnd11an1n64x5 FILLER_116_1238 ();
 b15zdnd11an1n64x5 FILLER_116_1302 ();
 b15zdnd11an1n64x5 FILLER_116_1366 ();
 b15zdnd11an1n32x5 FILLER_116_1430 ();
 b15zdnd11an1n16x5 FILLER_116_1462 ();
 b15zdnd11an1n08x5 FILLER_116_2265 ();
 b15zdnd00an1n02x5 FILLER_116_2273 ();
 b15zdnd00an1n01x5 FILLER_116_2275 ();
 b15zdnd11an1n64x5 FILLER_117_0 ();
 b15zdnd11an1n64x5 FILLER_117_64 ();
 b15zdnd11an1n64x5 FILLER_117_128 ();
 b15zdnd11an1n64x5 FILLER_117_192 ();
 b15zdnd11an1n64x5 FILLER_117_256 ();
 b15zdnd11an1n64x5 FILLER_117_320 ();
 b15zdnd11an1n64x5 FILLER_117_384 ();
 b15zdnd11an1n64x5 FILLER_117_448 ();
 b15zdnd11an1n64x5 FILLER_117_512 ();
 b15zdnd11an1n64x5 FILLER_117_576 ();
 b15zdnd11an1n64x5 FILLER_117_640 ();
 b15zdnd11an1n64x5 FILLER_117_704 ();
 b15zdnd11an1n64x5 FILLER_117_768 ();
 b15zdnd11an1n64x5 FILLER_117_832 ();
 b15zdnd11an1n64x5 FILLER_117_896 ();
 b15zdnd11an1n64x5 FILLER_117_960 ();
 b15zdnd11an1n64x5 FILLER_117_1024 ();
 b15zdnd11an1n32x5 FILLER_117_1088 ();
 b15zdnd11an1n08x5 FILLER_117_1120 ();
 b15zdnd00an1n02x5 FILLER_117_1128 ();
 b15zdnd11an1n64x5 FILLER_117_1141 ();
 b15zdnd11an1n64x5 FILLER_117_1205 ();
 b15zdnd11an1n64x5 FILLER_117_1269 ();
 b15zdnd11an1n64x5 FILLER_117_1333 ();
 b15zdnd11an1n64x5 FILLER_117_1397 ();
 b15zdnd11an1n08x5 FILLER_117_1461 ();
 b15zdnd11an1n04x5 FILLER_117_1469 ();
 b15zdnd00an1n02x5 FILLER_117_1473 ();
 b15zdnd00an1n01x5 FILLER_117_1475 ();
 b15zdnd00an1n02x5 FILLER_117_1484 ();
 b15zdnd11an1n16x5 FILLER_117_2257 ();
 b15zdnd11an1n08x5 FILLER_117_2273 ();
 b15zdnd00an1n02x5 FILLER_117_2281 ();
 b15zdnd00an1n01x5 FILLER_117_2283 ();
 b15zdnd11an1n64x5 FILLER_118_8 ();
 b15zdnd11an1n64x5 FILLER_118_72 ();
 b15zdnd11an1n64x5 FILLER_118_136 ();
 b15zdnd11an1n64x5 FILLER_118_200 ();
 b15zdnd11an1n64x5 FILLER_118_264 ();
 b15zdnd11an1n64x5 FILLER_118_328 ();
 b15zdnd11an1n64x5 FILLER_118_392 ();
 b15zdnd11an1n64x5 FILLER_118_456 ();
 b15zdnd11an1n64x5 FILLER_118_520 ();
 b15zdnd11an1n64x5 FILLER_118_584 ();
 b15zdnd11an1n64x5 FILLER_118_648 ();
 b15zdnd11an1n04x5 FILLER_118_712 ();
 b15zdnd00an1n02x5 FILLER_118_716 ();
 b15zdnd11an1n64x5 FILLER_118_726 ();
 b15zdnd11an1n64x5 FILLER_118_790 ();
 b15zdnd11an1n64x5 FILLER_118_854 ();
 b15zdnd11an1n64x5 FILLER_118_918 ();
 b15zdnd11an1n16x5 FILLER_118_982 ();
 b15zdnd00an1n02x5 FILLER_118_998 ();
 b15zdnd11an1n64x5 FILLER_118_1044 ();
 b15zdnd11an1n08x5 FILLER_118_1108 ();
 b15zdnd11an1n04x5 FILLER_118_1116 ();
 b15zdnd11an1n16x5 FILLER_118_1131 ();
 b15zdnd11an1n04x5 FILLER_118_1147 ();
 b15zdnd00an1n02x5 FILLER_118_1151 ();
 b15zdnd11an1n64x5 FILLER_118_1195 ();
 b15zdnd11an1n64x5 FILLER_118_1259 ();
 b15zdnd11an1n64x5 FILLER_118_1323 ();
 b15zdnd11an1n64x5 FILLER_118_1387 ();
 b15zdnd11an1n16x5 FILLER_118_1451 ();
 b15zdnd11an1n08x5 FILLER_118_1467 ();
 b15zdnd00an1n02x5 FILLER_118_1475 ();
 b15zdnd00an1n01x5 FILLER_118_1477 ();
 b15zdnd11an1n08x5 FILLER_118_2265 ();
 b15zdnd00an1n02x5 FILLER_118_2273 ();
 b15zdnd00an1n01x5 FILLER_118_2275 ();
 b15zdnd11an1n64x5 FILLER_119_0 ();
 b15zdnd11an1n64x5 FILLER_119_64 ();
 b15zdnd11an1n64x5 FILLER_119_128 ();
 b15zdnd11an1n64x5 FILLER_119_192 ();
 b15zdnd11an1n64x5 FILLER_119_256 ();
 b15zdnd11an1n64x5 FILLER_119_320 ();
 b15zdnd11an1n64x5 FILLER_119_384 ();
 b15zdnd11an1n64x5 FILLER_119_448 ();
 b15zdnd11an1n64x5 FILLER_119_512 ();
 b15zdnd11an1n64x5 FILLER_119_576 ();
 b15zdnd11an1n64x5 FILLER_119_640 ();
 b15zdnd11an1n64x5 FILLER_119_704 ();
 b15zdnd11an1n64x5 FILLER_119_768 ();
 b15zdnd11an1n64x5 FILLER_119_832 ();
 b15zdnd11an1n64x5 FILLER_119_896 ();
 b15zdnd11an1n32x5 FILLER_119_960 ();
 b15zdnd00an1n01x5 FILLER_119_992 ();
 b15zdnd11an1n64x5 FILLER_119_1037 ();
 b15zdnd11an1n64x5 FILLER_119_1101 ();
 b15zdnd11an1n64x5 FILLER_119_1165 ();
 b15zdnd11an1n64x5 FILLER_119_1229 ();
 b15zdnd11an1n64x5 FILLER_119_1293 ();
 b15zdnd11an1n64x5 FILLER_119_1357 ();
 b15zdnd11an1n64x5 FILLER_119_1421 ();
 b15zdnd00an1n01x5 FILLER_119_1485 ();
 b15zdnd11an1n16x5 FILLER_119_2257 ();
 b15zdnd11an1n08x5 FILLER_119_2273 ();
 b15zdnd00an1n02x5 FILLER_119_2281 ();
 b15zdnd00an1n01x5 FILLER_119_2283 ();
 b15zdnd11an1n64x5 FILLER_120_8 ();
 b15zdnd11an1n64x5 FILLER_120_72 ();
 b15zdnd11an1n64x5 FILLER_120_136 ();
 b15zdnd11an1n64x5 FILLER_120_200 ();
 b15zdnd11an1n64x5 FILLER_120_264 ();
 b15zdnd11an1n32x5 FILLER_120_328 ();
 b15zdnd11an1n16x5 FILLER_120_360 ();
 b15zdnd11an1n04x5 FILLER_120_376 ();
 b15zdnd00an1n01x5 FILLER_120_380 ();
 b15zdnd11an1n64x5 FILLER_120_401 ();
 b15zdnd11an1n64x5 FILLER_120_465 ();
 b15zdnd11an1n64x5 FILLER_120_529 ();
 b15zdnd11an1n64x5 FILLER_120_593 ();
 b15zdnd11an1n32x5 FILLER_120_657 ();
 b15zdnd11an1n16x5 FILLER_120_689 ();
 b15zdnd11an1n08x5 FILLER_120_705 ();
 b15zdnd11an1n04x5 FILLER_120_713 ();
 b15zdnd00an1n01x5 FILLER_120_717 ();
 b15zdnd11an1n64x5 FILLER_120_726 ();
 b15zdnd11an1n64x5 FILLER_120_790 ();
 b15zdnd11an1n64x5 FILLER_120_854 ();
 b15zdnd11an1n32x5 FILLER_120_918 ();
 b15zdnd11an1n08x5 FILLER_120_950 ();
 b15zdnd11an1n04x5 FILLER_120_958 ();
 b15zdnd11an1n32x5 FILLER_120_965 ();
 b15zdnd00an1n02x5 FILLER_120_997 ();
 b15zdnd00an1n01x5 FILLER_120_999 ();
 b15zdnd11an1n64x5 FILLER_120_1044 ();
 b15zdnd11an1n64x5 FILLER_120_1108 ();
 b15zdnd11an1n64x5 FILLER_120_1172 ();
 b15zdnd11an1n64x5 FILLER_120_1236 ();
 b15zdnd11an1n64x5 FILLER_120_1300 ();
 b15zdnd11an1n64x5 FILLER_120_1364 ();
 b15zdnd11an1n32x5 FILLER_120_1428 ();
 b15zdnd11an1n16x5 FILLER_120_1460 ();
 b15zdnd00an1n02x5 FILLER_120_1476 ();
 b15zdnd11an1n08x5 FILLER_120_2265 ();
 b15zdnd00an1n02x5 FILLER_120_2273 ();
 b15zdnd00an1n01x5 FILLER_120_2275 ();
 b15zdnd11an1n64x5 FILLER_121_0 ();
 b15zdnd11an1n64x5 FILLER_121_64 ();
 b15zdnd11an1n64x5 FILLER_121_128 ();
 b15zdnd11an1n64x5 FILLER_121_192 ();
 b15zdnd11an1n64x5 FILLER_121_256 ();
 b15zdnd11an1n64x5 FILLER_121_320 ();
 b15zdnd11an1n32x5 FILLER_121_384 ();
 b15zdnd11an1n16x5 FILLER_121_416 ();
 b15zdnd00an1n01x5 FILLER_121_432 ();
 b15zdnd11an1n64x5 FILLER_121_443 ();
 b15zdnd11an1n64x5 FILLER_121_507 ();
 b15zdnd11an1n64x5 FILLER_121_571 ();
 b15zdnd11an1n64x5 FILLER_121_635 ();
 b15zdnd11an1n64x5 FILLER_121_699 ();
 b15zdnd11an1n64x5 FILLER_121_763 ();
 b15zdnd11an1n64x5 FILLER_121_827 ();
 b15zdnd11an1n64x5 FILLER_121_891 ();
 b15zdnd11an1n04x5 FILLER_121_955 ();
 b15zdnd00an1n02x5 FILLER_121_959 ();
 b15zdnd00an1n01x5 FILLER_121_961 ();
 b15zdnd11an1n04x5 FILLER_121_989 ();
 b15zdnd11an1n04x5 FILLER_121_1037 ();
 b15zdnd11an1n04x5 FILLER_121_1044 ();
 b15zdnd11an1n64x5 FILLER_121_1051 ();
 b15zdnd11an1n64x5 FILLER_121_1115 ();
 b15zdnd11an1n64x5 FILLER_121_1179 ();
 b15zdnd11an1n64x5 FILLER_121_1243 ();
 b15zdnd11an1n64x5 FILLER_121_1307 ();
 b15zdnd11an1n64x5 FILLER_121_1371 ();
 b15zdnd11an1n16x5 FILLER_121_1435 ();
 b15zdnd11an1n08x5 FILLER_121_1451 ();
 b15zdnd11an1n04x5 FILLER_121_1459 ();
 b15zdnd00an1n01x5 FILLER_121_1463 ();
 b15zdnd11an1n08x5 FILLER_121_1475 ();
 b15zdnd00an1n02x5 FILLER_121_1483 ();
 b15zdnd00an1n01x5 FILLER_121_1485 ();
 b15zdnd11an1n16x5 FILLER_121_2257 ();
 b15zdnd11an1n08x5 FILLER_121_2273 ();
 b15zdnd00an1n02x5 FILLER_121_2281 ();
 b15zdnd00an1n01x5 FILLER_121_2283 ();
 b15zdnd11an1n64x5 FILLER_122_8 ();
 b15zdnd11an1n64x5 FILLER_122_72 ();
 b15zdnd11an1n64x5 FILLER_122_136 ();
 b15zdnd11an1n64x5 FILLER_122_200 ();
 b15zdnd11an1n64x5 FILLER_122_264 ();
 b15zdnd11an1n64x5 FILLER_122_328 ();
 b15zdnd11an1n04x5 FILLER_122_392 ();
 b15zdnd11an1n32x5 FILLER_122_402 ();
 b15zdnd11an1n08x5 FILLER_122_434 ();
 b15zdnd00an1n01x5 FILLER_122_442 ();
 b15zdnd11an1n64x5 FILLER_122_459 ();
 b15zdnd11an1n64x5 FILLER_122_523 ();
 b15zdnd11an1n64x5 FILLER_122_587 ();
 b15zdnd11an1n64x5 FILLER_122_651 ();
 b15zdnd00an1n02x5 FILLER_122_715 ();
 b15zdnd00an1n01x5 FILLER_122_717 ();
 b15zdnd11an1n64x5 FILLER_122_726 ();
 b15zdnd11an1n64x5 FILLER_122_790 ();
 b15zdnd11an1n64x5 FILLER_122_854 ();
 b15zdnd11an1n64x5 FILLER_122_918 ();
 b15zdnd11an1n04x5 FILLER_122_982 ();
 b15zdnd00an1n02x5 FILLER_122_986 ();
 b15zdnd11an1n04x5 FILLER_122_997 ();
 b15zdnd00an1n02x5 FILLER_122_1001 ();
 b15zdnd11an1n08x5 FILLER_122_1012 ();
 b15zdnd11an1n04x5 FILLER_122_1023 ();
 b15zdnd11an1n04x5 FILLER_122_1030 ();
 b15zdnd11an1n04x5 FILLER_122_1037 ();
 b15zdnd11an1n64x5 FILLER_122_1044 ();
 b15zdnd11an1n64x5 FILLER_122_1119 ();
 b15zdnd11an1n64x5 FILLER_122_1183 ();
 b15zdnd11an1n64x5 FILLER_122_1247 ();
 b15zdnd11an1n64x5 FILLER_122_1311 ();
 b15zdnd11an1n64x5 FILLER_122_1375 ();
 b15zdnd11an1n32x5 FILLER_122_1439 ();
 b15zdnd11an1n04x5 FILLER_122_1471 ();
 b15zdnd00an1n02x5 FILLER_122_1475 ();
 b15zdnd00an1n01x5 FILLER_122_1477 ();
 b15zdnd11an1n08x5 FILLER_122_2265 ();
 b15zdnd00an1n02x5 FILLER_122_2273 ();
 b15zdnd00an1n01x5 FILLER_122_2275 ();
 b15zdnd11an1n64x5 FILLER_123_0 ();
 b15zdnd11an1n64x5 FILLER_123_64 ();
 b15zdnd11an1n64x5 FILLER_123_128 ();
 b15zdnd11an1n64x5 FILLER_123_192 ();
 b15zdnd11an1n64x5 FILLER_123_256 ();
 b15zdnd11an1n64x5 FILLER_123_320 ();
 b15zdnd11an1n16x5 FILLER_123_384 ();
 b15zdnd00an1n02x5 FILLER_123_400 ();
 b15zdnd00an1n01x5 FILLER_123_402 ();
 b15zdnd11an1n64x5 FILLER_123_419 ();
 b15zdnd11an1n64x5 FILLER_123_483 ();
 b15zdnd11an1n64x5 FILLER_123_547 ();
 b15zdnd11an1n64x5 FILLER_123_611 ();
 b15zdnd11an1n64x5 FILLER_123_675 ();
 b15zdnd11an1n64x5 FILLER_123_739 ();
 b15zdnd11an1n64x5 FILLER_123_803 ();
 b15zdnd11an1n64x5 FILLER_123_867 ();
 b15zdnd11an1n64x5 FILLER_123_931 ();
 b15zdnd11an1n08x5 FILLER_123_995 ();
 b15zdnd11an1n04x5 FILLER_123_1006 ();
 b15zdnd11an1n04x5 FILLER_123_1013 ();
 b15zdnd11an1n04x5 FILLER_123_1020 ();
 b15zdnd11an1n04x5 FILLER_123_1027 ();
 b15zdnd11an1n64x5 FILLER_123_1034 ();
 b15zdnd11an1n64x5 FILLER_123_1098 ();
 b15zdnd11an1n64x5 FILLER_123_1162 ();
 b15zdnd11an1n64x5 FILLER_123_1226 ();
 b15zdnd11an1n64x5 FILLER_123_1290 ();
 b15zdnd11an1n64x5 FILLER_123_1354 ();
 b15zdnd11an1n32x5 FILLER_123_1418 ();
 b15zdnd11an1n16x5 FILLER_123_1450 ();
 b15zdnd11an1n04x5 FILLER_123_1466 ();
 b15zdnd00an1n02x5 FILLER_123_1470 ();
 b15zdnd00an1n01x5 FILLER_123_1472 ();
 b15zdnd00an1n02x5 FILLER_123_1484 ();
 b15zdnd11an1n16x5 FILLER_123_2257 ();
 b15zdnd11an1n08x5 FILLER_123_2273 ();
 b15zdnd00an1n02x5 FILLER_123_2281 ();
 b15zdnd00an1n01x5 FILLER_123_2283 ();
 b15zdnd11an1n64x5 FILLER_124_8 ();
 b15zdnd11an1n64x5 FILLER_124_72 ();
 b15zdnd11an1n64x5 FILLER_124_136 ();
 b15zdnd11an1n64x5 FILLER_124_200 ();
 b15zdnd11an1n64x5 FILLER_124_264 ();
 b15zdnd11an1n64x5 FILLER_124_328 ();
 b15zdnd11an1n32x5 FILLER_124_392 ();
 b15zdnd11an1n16x5 FILLER_124_424 ();
 b15zdnd00an1n02x5 FILLER_124_440 ();
 b15zdnd00an1n01x5 FILLER_124_442 ();
 b15zdnd11an1n64x5 FILLER_124_455 ();
 b15zdnd11an1n64x5 FILLER_124_519 ();
 b15zdnd11an1n64x5 FILLER_124_583 ();
 b15zdnd11an1n64x5 FILLER_124_647 ();
 b15zdnd11an1n04x5 FILLER_124_711 ();
 b15zdnd00an1n02x5 FILLER_124_715 ();
 b15zdnd00an1n01x5 FILLER_124_717 ();
 b15zdnd11an1n64x5 FILLER_124_726 ();
 b15zdnd11an1n64x5 FILLER_124_790 ();
 b15zdnd11an1n64x5 FILLER_124_854 ();
 b15zdnd11an1n64x5 FILLER_124_918 ();
 b15zdnd11an1n16x5 FILLER_124_982 ();
 b15zdnd11an1n08x5 FILLER_124_998 ();
 b15zdnd11an1n04x5 FILLER_124_1006 ();
 b15zdnd00an1n02x5 FILLER_124_1010 ();
 b15zdnd00an1n01x5 FILLER_124_1012 ();
 b15zdnd11an1n04x5 FILLER_124_1016 ();
 b15zdnd00an1n02x5 FILLER_124_1020 ();
 b15zdnd00an1n01x5 FILLER_124_1022 ();
 b15zdnd11an1n64x5 FILLER_124_1026 ();
 b15zdnd11an1n64x5 FILLER_124_1090 ();
 b15zdnd11an1n64x5 FILLER_124_1154 ();
 b15zdnd11an1n64x5 FILLER_124_1218 ();
 b15zdnd11an1n64x5 FILLER_124_1282 ();
 b15zdnd11an1n64x5 FILLER_124_1346 ();
 b15zdnd11an1n64x5 FILLER_124_1410 ();
 b15zdnd11an1n04x5 FILLER_124_1474 ();
 b15zdnd11an1n08x5 FILLER_124_2265 ();
 b15zdnd00an1n02x5 FILLER_124_2273 ();
 b15zdnd00an1n01x5 FILLER_124_2275 ();
 b15zdnd11an1n64x5 FILLER_125_0 ();
 b15zdnd11an1n64x5 FILLER_125_64 ();
 b15zdnd11an1n64x5 FILLER_125_128 ();
 b15zdnd11an1n64x5 FILLER_125_192 ();
 b15zdnd11an1n64x5 FILLER_125_256 ();
 b15zdnd11an1n64x5 FILLER_125_320 ();
 b15zdnd11an1n32x5 FILLER_125_384 ();
 b15zdnd11an1n16x5 FILLER_125_416 ();
 b15zdnd11an1n08x5 FILLER_125_432 ();
 b15zdnd00an1n01x5 FILLER_125_440 ();
 b15zdnd11an1n64x5 FILLER_125_451 ();
 b15zdnd11an1n32x5 FILLER_125_515 ();
 b15zdnd11an1n16x5 FILLER_125_547 ();
 b15zdnd11an1n08x5 FILLER_125_563 ();
 b15zdnd11an1n04x5 FILLER_125_571 ();
 b15zdnd11an1n64x5 FILLER_125_617 ();
 b15zdnd11an1n64x5 FILLER_125_681 ();
 b15zdnd11an1n64x5 FILLER_125_745 ();
 b15zdnd11an1n64x5 FILLER_125_809 ();
 b15zdnd11an1n64x5 FILLER_125_873 ();
 b15zdnd11an1n64x5 FILLER_125_937 ();
 b15zdnd11an1n64x5 FILLER_125_1001 ();
 b15zdnd11an1n64x5 FILLER_125_1065 ();
 b15zdnd11an1n64x5 FILLER_125_1129 ();
 b15zdnd11an1n64x5 FILLER_125_1193 ();
 b15zdnd00an1n02x5 FILLER_125_1257 ();
 b15zdnd00an1n01x5 FILLER_125_1259 ();
 b15zdnd11an1n04x5 FILLER_125_1263 ();
 b15zdnd11an1n64x5 FILLER_125_1270 ();
 b15zdnd11an1n32x5 FILLER_125_1334 ();
 b15zdnd11an1n16x5 FILLER_125_1366 ();
 b15zdnd11an1n08x5 FILLER_125_1382 ();
 b15zdnd00an1n02x5 FILLER_125_1390 ();
 b15zdnd00an1n01x5 FILLER_125_1392 ();
 b15zdnd11an1n32x5 FILLER_125_1435 ();
 b15zdnd11an1n16x5 FILLER_125_1467 ();
 b15zdnd00an1n02x5 FILLER_125_1483 ();
 b15zdnd00an1n01x5 FILLER_125_1485 ();
 b15zdnd11an1n04x5 FILLER_125_2257 ();
 b15zdnd00an1n02x5 FILLER_125_2261 ();
 b15zdnd00an1n01x5 FILLER_125_2263 ();
 b15zdnd11an1n08x5 FILLER_125_2271 ();
 b15zdnd11an1n04x5 FILLER_125_2279 ();
 b15zdnd00an1n01x5 FILLER_125_2283 ();
 b15zdnd11an1n64x5 FILLER_126_8 ();
 b15zdnd11an1n64x5 FILLER_126_72 ();
 b15zdnd11an1n64x5 FILLER_126_136 ();
 b15zdnd11an1n64x5 FILLER_126_200 ();
 b15zdnd11an1n64x5 FILLER_126_264 ();
 b15zdnd11an1n64x5 FILLER_126_328 ();
 b15zdnd11an1n64x5 FILLER_126_392 ();
 b15zdnd11an1n64x5 FILLER_126_456 ();
 b15zdnd11an1n32x5 FILLER_126_520 ();
 b15zdnd11an1n04x5 FILLER_126_552 ();
 b15zdnd00an1n02x5 FILLER_126_556 ();
 b15zdnd11an1n32x5 FILLER_126_600 ();
 b15zdnd11an1n16x5 FILLER_126_632 ();
 b15zdnd11an1n04x5 FILLER_126_648 ();
 b15zdnd00an1n02x5 FILLER_126_652 ();
 b15zdnd00an1n01x5 FILLER_126_654 ();
 b15zdnd11an1n32x5 FILLER_126_664 ();
 b15zdnd11an1n16x5 FILLER_126_696 ();
 b15zdnd11an1n04x5 FILLER_126_712 ();
 b15zdnd00an1n02x5 FILLER_126_716 ();
 b15zdnd11an1n64x5 FILLER_126_726 ();
 b15zdnd11an1n64x5 FILLER_126_790 ();
 b15zdnd11an1n64x5 FILLER_126_854 ();
 b15zdnd11an1n64x5 FILLER_126_918 ();
 b15zdnd11an1n32x5 FILLER_126_982 ();
 b15zdnd11an1n16x5 FILLER_126_1014 ();
 b15zdnd11an1n04x5 FILLER_126_1030 ();
 b15zdnd00an1n02x5 FILLER_126_1034 ();
 b15zdnd00an1n01x5 FILLER_126_1036 ();
 b15zdnd11an1n64x5 FILLER_126_1079 ();
 b15zdnd11an1n64x5 FILLER_126_1143 ();
 b15zdnd11an1n32x5 FILLER_126_1207 ();
 b15zdnd00an1n02x5 FILLER_126_1239 ();
 b15zdnd11an1n64x5 FILLER_126_1273 ();
 b15zdnd11an1n16x5 FILLER_126_1337 ();
 b15zdnd11an1n32x5 FILLER_126_1405 ();
 b15zdnd11an1n16x5 FILLER_126_1437 ();
 b15zdnd11an1n08x5 FILLER_126_1453 ();
 b15zdnd11an1n04x5 FILLER_126_1461 ();
 b15zdnd00an1n02x5 FILLER_126_1476 ();
 b15zdnd11an1n08x5 FILLER_126_2265 ();
 b15zdnd00an1n02x5 FILLER_126_2273 ();
 b15zdnd00an1n01x5 FILLER_126_2275 ();
 b15zdnd11an1n64x5 FILLER_127_0 ();
 b15zdnd11an1n64x5 FILLER_127_64 ();
 b15zdnd11an1n64x5 FILLER_127_128 ();
 b15zdnd11an1n64x5 FILLER_127_192 ();
 b15zdnd11an1n64x5 FILLER_127_256 ();
 b15zdnd11an1n64x5 FILLER_127_320 ();
 b15zdnd11an1n64x5 FILLER_127_384 ();
 b15zdnd11an1n64x5 FILLER_127_448 ();
 b15zdnd11an1n64x5 FILLER_127_512 ();
 b15zdnd11an1n04x5 FILLER_127_576 ();
 b15zdnd11an1n16x5 FILLER_127_622 ();
 b15zdnd11an1n08x5 FILLER_127_638 ();
 b15zdnd11an1n04x5 FILLER_127_688 ();
 b15zdnd11an1n64x5 FILLER_127_695 ();
 b15zdnd11an1n64x5 FILLER_127_759 ();
 b15zdnd11an1n64x5 FILLER_127_823 ();
 b15zdnd11an1n64x5 FILLER_127_887 ();
 b15zdnd11an1n64x5 FILLER_127_951 ();
 b15zdnd11an1n64x5 FILLER_127_1015 ();
 b15zdnd11an1n64x5 FILLER_127_1079 ();
 b15zdnd11an1n64x5 FILLER_127_1143 ();
 b15zdnd11an1n64x5 FILLER_127_1207 ();
 b15zdnd11an1n64x5 FILLER_127_1274 ();
 b15zdnd11an1n32x5 FILLER_127_1338 ();
 b15zdnd00an1n02x5 FILLER_127_1370 ();
 b15zdnd11an1n04x5 FILLER_127_1375 ();
 b15zdnd11an1n64x5 FILLER_127_1382 ();
 b15zdnd11an1n32x5 FILLER_127_1446 ();
 b15zdnd11an1n08x5 FILLER_127_1478 ();
 b15zdnd11an1n08x5 FILLER_127_2257 ();
 b15zdnd00an1n02x5 FILLER_127_2265 ();
 b15zdnd11an1n08x5 FILLER_127_2274 ();
 b15zdnd00an1n02x5 FILLER_127_2282 ();
 b15zdnd11an1n64x5 FILLER_128_8 ();
 b15zdnd11an1n64x5 FILLER_128_72 ();
 b15zdnd11an1n64x5 FILLER_128_136 ();
 b15zdnd11an1n64x5 FILLER_128_200 ();
 b15zdnd11an1n64x5 FILLER_128_264 ();
 b15zdnd11an1n64x5 FILLER_128_328 ();
 b15zdnd11an1n64x5 FILLER_128_392 ();
 b15zdnd11an1n64x5 FILLER_128_456 ();
 b15zdnd11an1n64x5 FILLER_128_520 ();
 b15zdnd11an1n32x5 FILLER_128_584 ();
 b15zdnd11an1n08x5 FILLER_128_658 ();
 b15zdnd11an1n04x5 FILLER_128_666 ();
 b15zdnd00an1n02x5 FILLER_128_670 ();
 b15zdnd00an1n02x5 FILLER_128_716 ();
 b15zdnd11an1n64x5 FILLER_128_726 ();
 b15zdnd11an1n64x5 FILLER_128_790 ();
 b15zdnd11an1n64x5 FILLER_128_854 ();
 b15zdnd11an1n64x5 FILLER_128_918 ();
 b15zdnd11an1n64x5 FILLER_128_982 ();
 b15zdnd11an1n64x5 FILLER_128_1046 ();
 b15zdnd11an1n64x5 FILLER_128_1110 ();
 b15zdnd11an1n64x5 FILLER_128_1174 ();
 b15zdnd11an1n08x5 FILLER_128_1238 ();
 b15zdnd11an1n04x5 FILLER_128_1246 ();
 b15zdnd00an1n02x5 FILLER_128_1250 ();
 b15zdnd11an1n04x5 FILLER_128_1255 ();
 b15zdnd11an1n64x5 FILLER_128_1262 ();
 b15zdnd11an1n32x5 FILLER_128_1326 ();
 b15zdnd11an1n16x5 FILLER_128_1358 ();
 b15zdnd11an1n04x5 FILLER_128_1374 ();
 b15zdnd11an1n64x5 FILLER_128_1381 ();
 b15zdnd11an1n32x5 FILLER_128_1445 ();
 b15zdnd00an1n01x5 FILLER_128_1477 ();
 b15zdnd11an1n08x5 FILLER_128_2265 ();
 b15zdnd00an1n02x5 FILLER_128_2273 ();
 b15zdnd00an1n01x5 FILLER_128_2275 ();
 b15zdnd11an1n64x5 FILLER_129_0 ();
 b15zdnd11an1n64x5 FILLER_129_64 ();
 b15zdnd11an1n64x5 FILLER_129_128 ();
 b15zdnd11an1n64x5 FILLER_129_192 ();
 b15zdnd11an1n64x5 FILLER_129_256 ();
 b15zdnd11an1n64x5 FILLER_129_320 ();
 b15zdnd11an1n64x5 FILLER_129_384 ();
 b15zdnd11an1n64x5 FILLER_129_448 ();
 b15zdnd11an1n32x5 FILLER_129_512 ();
 b15zdnd11an1n08x5 FILLER_129_544 ();
 b15zdnd11an1n04x5 FILLER_129_552 ();
 b15zdnd00an1n02x5 FILLER_129_556 ();
 b15zdnd00an1n01x5 FILLER_129_558 ();
 b15zdnd11an1n32x5 FILLER_129_601 ();
 b15zdnd11an1n16x5 FILLER_129_633 ();
 b15zdnd11an1n04x5 FILLER_129_676 ();
 b15zdnd11an1n04x5 FILLER_129_705 ();
 b15zdnd11an1n64x5 FILLER_129_712 ();
 b15zdnd11an1n64x5 FILLER_129_776 ();
 b15zdnd11an1n64x5 FILLER_129_840 ();
 b15zdnd11an1n64x5 FILLER_129_904 ();
 b15zdnd11an1n64x5 FILLER_129_968 ();
 b15zdnd11an1n64x5 FILLER_129_1032 ();
 b15zdnd11an1n64x5 FILLER_129_1096 ();
 b15zdnd11an1n64x5 FILLER_129_1160 ();
 b15zdnd11an1n04x5 FILLER_129_1224 ();
 b15zdnd00an1n01x5 FILLER_129_1228 ();
 b15zdnd11an1n64x5 FILLER_129_1261 ();
 b15zdnd11an1n64x5 FILLER_129_1325 ();
 b15zdnd11an1n64x5 FILLER_129_1389 ();
 b15zdnd11an1n32x5 FILLER_129_1453 ();
 b15zdnd00an1n01x5 FILLER_129_1485 ();
 b15zdnd00an1n02x5 FILLER_129_2257 ();
 b15zdnd00an1n01x5 FILLER_129_2259 ();
 b15zdnd11an1n16x5 FILLER_129_2267 ();
 b15zdnd00an1n01x5 FILLER_129_2283 ();
 b15zdnd11an1n16x5 FILLER_130_8 ();
 b15zdnd11an1n04x5 FILLER_130_24 ();
 b15zdnd00an1n02x5 FILLER_130_28 ();
 b15zdnd00an1n01x5 FILLER_130_30 ();
 b15zdnd11an1n64x5 FILLER_130_35 ();
 b15zdnd11an1n32x5 FILLER_130_99 ();
 b15zdnd00an1n02x5 FILLER_130_131 ();
 b15zdnd11an1n64x5 FILLER_130_151 ();
 b15zdnd11an1n64x5 FILLER_130_215 ();
 b15zdnd11an1n64x5 FILLER_130_279 ();
 b15zdnd11an1n64x5 FILLER_130_343 ();
 b15zdnd11an1n64x5 FILLER_130_407 ();
 b15zdnd11an1n64x5 FILLER_130_471 ();
 b15zdnd11an1n64x5 FILLER_130_535 ();
 b15zdnd11an1n32x5 FILLER_130_599 ();
 b15zdnd11an1n16x5 FILLER_130_631 ();
 b15zdnd00an1n01x5 FILLER_130_647 ();
 b15zdnd11an1n04x5 FILLER_130_690 ();
 b15zdnd11an1n04x5 FILLER_130_703 ();
 b15zdnd11an1n08x5 FILLER_130_710 ();
 b15zdnd11an1n64x5 FILLER_130_726 ();
 b15zdnd11an1n64x5 FILLER_130_790 ();
 b15zdnd11an1n64x5 FILLER_130_854 ();
 b15zdnd11an1n64x5 FILLER_130_918 ();
 b15zdnd11an1n32x5 FILLER_130_982 ();
 b15zdnd11an1n08x5 FILLER_130_1014 ();
 b15zdnd11an1n04x5 FILLER_130_1022 ();
 b15zdnd00an1n02x5 FILLER_130_1026 ();
 b15zdnd00an1n01x5 FILLER_130_1028 ();
 b15zdnd11an1n64x5 FILLER_130_1037 ();
 b15zdnd11an1n64x5 FILLER_130_1101 ();
 b15zdnd11an1n64x5 FILLER_130_1165 ();
 b15zdnd11an1n16x5 FILLER_130_1229 ();
 b15zdnd11an1n08x5 FILLER_130_1245 ();
 b15zdnd00an1n02x5 FILLER_130_1253 ();
 b15zdnd11an1n64x5 FILLER_130_1258 ();
 b15zdnd11an1n64x5 FILLER_130_1322 ();
 b15zdnd11an1n64x5 FILLER_130_1386 ();
 b15zdnd11an1n16x5 FILLER_130_1450 ();
 b15zdnd11an1n08x5 FILLER_130_1466 ();
 b15zdnd11an1n04x5 FILLER_130_1474 ();
 b15zdnd11an1n08x5 FILLER_130_2265 ();
 b15zdnd00an1n02x5 FILLER_130_2273 ();
 b15zdnd00an1n01x5 FILLER_130_2275 ();
 b15zdnd11an1n08x5 FILLER_131_0 ();
 b15zdnd00an1n02x5 FILLER_131_8 ();
 b15zdnd00an1n01x5 FILLER_131_10 ();
 b15zdnd11an1n64x5 FILLER_131_53 ();
 b15zdnd11an1n64x5 FILLER_131_117 ();
 b15zdnd11an1n64x5 FILLER_131_181 ();
 b15zdnd11an1n64x5 FILLER_131_245 ();
 b15zdnd11an1n64x5 FILLER_131_309 ();
 b15zdnd11an1n32x5 FILLER_131_373 ();
 b15zdnd11an1n16x5 FILLER_131_405 ();
 b15zdnd00an1n02x5 FILLER_131_421 ();
 b15zdnd11an1n64x5 FILLER_131_445 ();
 b15zdnd11an1n64x5 FILLER_131_509 ();
 b15zdnd11an1n32x5 FILLER_131_573 ();
 b15zdnd11an1n08x5 FILLER_131_605 ();
 b15zdnd11an1n04x5 FILLER_131_613 ();
 b15zdnd11an1n16x5 FILLER_131_659 ();
 b15zdnd11an1n04x5 FILLER_131_675 ();
 b15zdnd00an1n01x5 FILLER_131_679 ();
 b15zdnd11an1n04x5 FILLER_131_724 ();
 b15zdnd11an1n64x5 FILLER_131_731 ();
 b15zdnd11an1n64x5 FILLER_131_795 ();
 b15zdnd11an1n64x5 FILLER_131_859 ();
 b15zdnd11an1n64x5 FILLER_131_923 ();
 b15zdnd11an1n64x5 FILLER_131_987 ();
 b15zdnd11an1n64x5 FILLER_131_1051 ();
 b15zdnd11an1n64x5 FILLER_131_1115 ();
 b15zdnd11an1n64x5 FILLER_131_1179 ();
 b15zdnd11an1n64x5 FILLER_131_1243 ();
 b15zdnd11an1n64x5 FILLER_131_1307 ();
 b15zdnd11an1n64x5 FILLER_131_1371 ();
 b15zdnd11an1n32x5 FILLER_131_1435 ();
 b15zdnd11an1n16x5 FILLER_131_1467 ();
 b15zdnd00an1n02x5 FILLER_131_1483 ();
 b15zdnd00an1n01x5 FILLER_131_1485 ();
 b15zdnd11an1n16x5 FILLER_131_2257 ();
 b15zdnd11an1n08x5 FILLER_131_2273 ();
 b15zdnd00an1n02x5 FILLER_131_2281 ();
 b15zdnd00an1n01x5 FILLER_131_2283 ();
 b15zdnd11an1n16x5 FILLER_132_8 ();
 b15zdnd00an1n02x5 FILLER_132_24 ();
 b15zdnd11an1n64x5 FILLER_132_38 ();
 b15zdnd11an1n64x5 FILLER_132_102 ();
 b15zdnd11an1n64x5 FILLER_132_166 ();
 b15zdnd11an1n64x5 FILLER_132_230 ();
 b15zdnd11an1n64x5 FILLER_132_294 ();
 b15zdnd11an1n32x5 FILLER_132_358 ();
 b15zdnd11an1n08x5 FILLER_132_390 ();
 b15zdnd11an1n04x5 FILLER_132_398 ();
 b15zdnd00an1n02x5 FILLER_132_402 ();
 b15zdnd00an1n01x5 FILLER_132_404 ();
 b15zdnd11an1n64x5 FILLER_132_417 ();
 b15zdnd11an1n64x5 FILLER_132_481 ();
 b15zdnd11an1n64x5 FILLER_132_545 ();
 b15zdnd11an1n32x5 FILLER_132_609 ();
 b15zdnd00an1n01x5 FILLER_132_641 ();
 b15zdnd11an1n16x5 FILLER_132_645 ();
 b15zdnd11an1n04x5 FILLER_132_661 ();
 b15zdnd11an1n04x5 FILLER_132_668 ();
 b15zdnd00an1n02x5 FILLER_132_716 ();
 b15zdnd00an1n02x5 FILLER_132_726 ();
 b15zdnd11an1n64x5 FILLER_132_731 ();
 b15zdnd11an1n64x5 FILLER_132_795 ();
 b15zdnd11an1n64x5 FILLER_132_859 ();
 b15zdnd11an1n64x5 FILLER_132_923 ();
 b15zdnd11an1n64x5 FILLER_132_987 ();
 b15zdnd11an1n64x5 FILLER_132_1051 ();
 b15zdnd11an1n64x5 FILLER_132_1115 ();
 b15zdnd11an1n64x5 FILLER_132_1179 ();
 b15zdnd11an1n64x5 FILLER_132_1243 ();
 b15zdnd11an1n64x5 FILLER_132_1307 ();
 b15zdnd11an1n64x5 FILLER_132_1371 ();
 b15zdnd11an1n32x5 FILLER_132_1435 ();
 b15zdnd11an1n08x5 FILLER_132_1467 ();
 b15zdnd00an1n02x5 FILLER_132_1475 ();
 b15zdnd00an1n01x5 FILLER_132_1477 ();
 b15zdnd11an1n08x5 FILLER_132_2265 ();
 b15zdnd00an1n02x5 FILLER_132_2273 ();
 b15zdnd00an1n01x5 FILLER_132_2275 ();
 b15zdnd11an1n08x5 FILLER_133_0 ();
 b15zdnd11an1n04x5 FILLER_133_8 ();
 b15zdnd00an1n01x5 FILLER_133_12 ();
 b15zdnd11an1n64x5 FILLER_133_17 ();
 b15zdnd11an1n64x5 FILLER_133_81 ();
 b15zdnd11an1n64x5 FILLER_133_145 ();
 b15zdnd11an1n64x5 FILLER_133_209 ();
 b15zdnd11an1n64x5 FILLER_133_273 ();
 b15zdnd11an1n64x5 FILLER_133_337 ();
 b15zdnd11an1n64x5 FILLER_133_401 ();
 b15zdnd11an1n64x5 FILLER_133_465 ();
 b15zdnd11an1n64x5 FILLER_133_529 ();
 b15zdnd11an1n64x5 FILLER_133_593 ();
 b15zdnd11an1n04x5 FILLER_133_657 ();
 b15zdnd00an1n02x5 FILLER_133_661 ();
 b15zdnd00an1n01x5 FILLER_133_663 ();
 b15zdnd11an1n08x5 FILLER_133_667 ();
 b15zdnd11an1n04x5 FILLER_133_675 ();
 b15zdnd00an1n01x5 FILLER_133_679 ();
 b15zdnd11an1n04x5 FILLER_133_724 ();
 b15zdnd11an1n64x5 FILLER_133_731 ();
 b15zdnd11an1n64x5 FILLER_133_795 ();
 b15zdnd11an1n64x5 FILLER_133_859 ();
 b15zdnd11an1n64x5 FILLER_133_923 ();
 b15zdnd11an1n64x5 FILLER_133_987 ();
 b15zdnd11an1n64x5 FILLER_133_1051 ();
 b15zdnd11an1n64x5 FILLER_133_1115 ();
 b15zdnd11an1n64x5 FILLER_133_1179 ();
 b15zdnd11an1n64x5 FILLER_133_1243 ();
 b15zdnd11an1n64x5 FILLER_133_1307 ();
 b15zdnd11an1n64x5 FILLER_133_1371 ();
 b15zdnd11an1n32x5 FILLER_133_1435 ();
 b15zdnd11an1n16x5 FILLER_133_1467 ();
 b15zdnd00an1n02x5 FILLER_133_1483 ();
 b15zdnd00an1n01x5 FILLER_133_1485 ();
 b15zdnd11an1n16x5 FILLER_133_2257 ();
 b15zdnd11an1n08x5 FILLER_133_2273 ();
 b15zdnd00an1n02x5 FILLER_133_2281 ();
 b15zdnd00an1n01x5 FILLER_133_2283 ();
 b15zdnd11an1n64x5 FILLER_134_8 ();
 b15zdnd11an1n64x5 FILLER_134_72 ();
 b15zdnd11an1n04x5 FILLER_134_136 ();
 b15zdnd00an1n02x5 FILLER_134_140 ();
 b15zdnd00an1n01x5 FILLER_134_142 ();
 b15zdnd11an1n64x5 FILLER_134_165 ();
 b15zdnd11an1n04x5 FILLER_134_229 ();
 b15zdnd11an1n64x5 FILLER_134_247 ();
 b15zdnd11an1n32x5 FILLER_134_311 ();
 b15zdnd11an1n04x5 FILLER_134_343 ();
 b15zdnd11an1n64x5 FILLER_134_369 ();
 b15zdnd11an1n64x5 FILLER_134_433 ();
 b15zdnd11an1n64x5 FILLER_134_497 ();
 b15zdnd11an1n64x5 FILLER_134_561 ();
 b15zdnd11an1n64x5 FILLER_134_625 ();
 b15zdnd00an1n01x5 FILLER_134_689 ();
 b15zdnd11an1n04x5 FILLER_134_693 ();
 b15zdnd11an1n04x5 FILLER_134_700 ();
 b15zdnd11an1n04x5 FILLER_134_707 ();
 b15zdnd11an1n04x5 FILLER_134_714 ();
 b15zdnd11an1n64x5 FILLER_134_726 ();
 b15zdnd11an1n64x5 FILLER_134_790 ();
 b15zdnd11an1n64x5 FILLER_134_854 ();
 b15zdnd11an1n64x5 FILLER_134_918 ();
 b15zdnd11an1n64x5 FILLER_134_982 ();
 b15zdnd11an1n64x5 FILLER_134_1046 ();
 b15zdnd11an1n64x5 FILLER_134_1110 ();
 b15zdnd11an1n64x5 FILLER_134_1174 ();
 b15zdnd11an1n32x5 FILLER_134_1238 ();
 b15zdnd11an1n04x5 FILLER_134_1270 ();
 b15zdnd00an1n01x5 FILLER_134_1274 ();
 b15zdnd11an1n04x5 FILLER_134_1278 ();
 b15zdnd11an1n64x5 FILLER_134_1285 ();
 b15zdnd11an1n64x5 FILLER_134_1349 ();
 b15zdnd11an1n64x5 FILLER_134_1413 ();
 b15zdnd00an1n01x5 FILLER_134_1477 ();
 b15zdnd11an1n08x5 FILLER_134_2265 ();
 b15zdnd00an1n02x5 FILLER_134_2273 ();
 b15zdnd00an1n01x5 FILLER_134_2275 ();
 b15zdnd11an1n08x5 FILLER_135_0 ();
 b15zdnd00an1n02x5 FILLER_135_8 ();
 b15zdnd11an1n08x5 FILLER_135_14 ();
 b15zdnd11an1n04x5 FILLER_135_22 ();
 b15zdnd00an1n02x5 FILLER_135_26 ();
 b15zdnd11an1n04x5 FILLER_135_32 ();
 b15zdnd11an1n32x5 FILLER_135_40 ();
 b15zdnd11an1n16x5 FILLER_135_72 ();
 b15zdnd11an1n08x5 FILLER_135_88 ();
 b15zdnd00an1n01x5 FILLER_135_96 ();
 b15zdnd11an1n64x5 FILLER_135_109 ();
 b15zdnd11an1n64x5 FILLER_135_173 ();
 b15zdnd11an1n64x5 FILLER_135_237 ();
 b15zdnd11an1n64x5 FILLER_135_301 ();
 b15zdnd11an1n16x5 FILLER_135_365 ();
 b15zdnd11an1n08x5 FILLER_135_381 ();
 b15zdnd11an1n04x5 FILLER_135_389 ();
 b15zdnd11an1n04x5 FILLER_135_396 ();
 b15zdnd11an1n64x5 FILLER_135_414 ();
 b15zdnd11an1n64x5 FILLER_135_478 ();
 b15zdnd11an1n64x5 FILLER_135_542 ();
 b15zdnd11an1n64x5 FILLER_135_606 ();
 b15zdnd11an1n08x5 FILLER_135_670 ();
 b15zdnd11an1n04x5 FILLER_135_678 ();
 b15zdnd11an1n08x5 FILLER_135_691 ();
 b15zdnd00an1n02x5 FILLER_135_699 ();
 b15zdnd11an1n04x5 FILLER_135_704 ();
 b15zdnd11an1n64x5 FILLER_135_711 ();
 b15zdnd11an1n64x5 FILLER_135_775 ();
 b15zdnd11an1n64x5 FILLER_135_839 ();
 b15zdnd11an1n64x5 FILLER_135_903 ();
 b15zdnd11an1n64x5 FILLER_135_967 ();
 b15zdnd11an1n64x5 FILLER_135_1031 ();
 b15zdnd11an1n64x5 FILLER_135_1095 ();
 b15zdnd11an1n64x5 FILLER_135_1159 ();
 b15zdnd11an1n32x5 FILLER_135_1223 ();
 b15zdnd00an1n01x5 FILLER_135_1255 ();
 b15zdnd11an1n64x5 FILLER_135_1288 ();
 b15zdnd11an1n64x5 FILLER_135_1352 ();
 b15zdnd11an1n32x5 FILLER_135_1416 ();
 b15zdnd11an1n16x5 FILLER_135_1448 ();
 b15zdnd11an1n08x5 FILLER_135_1464 ();
 b15zdnd00an1n02x5 FILLER_135_1472 ();
 b15zdnd00an1n01x5 FILLER_135_1474 ();
 b15zdnd00an1n02x5 FILLER_135_1484 ();
 b15zdnd11an1n16x5 FILLER_135_2257 ();
 b15zdnd11an1n08x5 FILLER_135_2273 ();
 b15zdnd00an1n02x5 FILLER_135_2281 ();
 b15zdnd00an1n01x5 FILLER_135_2283 ();
 b15zdnd00an1n02x5 FILLER_136_8 ();
 b15zdnd11an1n04x5 FILLER_136_18 ();
 b15zdnd00an1n02x5 FILLER_136_22 ();
 b15zdnd11an1n64x5 FILLER_136_32 ();
 b15zdnd11an1n04x5 FILLER_136_96 ();
 b15zdnd00an1n02x5 FILLER_136_100 ();
 b15zdnd11an1n64x5 FILLER_136_109 ();
 b15zdnd11an1n64x5 FILLER_136_173 ();
 b15zdnd11an1n64x5 FILLER_136_237 ();
 b15zdnd11an1n32x5 FILLER_136_301 ();
 b15zdnd11an1n16x5 FILLER_136_333 ();
 b15zdnd00an1n02x5 FILLER_136_349 ();
 b15zdnd00an1n01x5 FILLER_136_351 ();
 b15zdnd11an1n64x5 FILLER_136_362 ();
 b15zdnd11an1n64x5 FILLER_136_426 ();
 b15zdnd11an1n64x5 FILLER_136_490 ();
 b15zdnd11an1n64x5 FILLER_136_554 ();
 b15zdnd11an1n64x5 FILLER_136_618 ();
 b15zdnd11an1n32x5 FILLER_136_682 ();
 b15zdnd11an1n04x5 FILLER_136_714 ();
 b15zdnd11an1n64x5 FILLER_136_726 ();
 b15zdnd11an1n64x5 FILLER_136_790 ();
 b15zdnd11an1n64x5 FILLER_136_854 ();
 b15zdnd11an1n64x5 FILLER_136_918 ();
 b15zdnd11an1n64x5 FILLER_136_982 ();
 b15zdnd11an1n64x5 FILLER_136_1046 ();
 b15zdnd11an1n64x5 FILLER_136_1110 ();
 b15zdnd11an1n64x5 FILLER_136_1174 ();
 b15zdnd11an1n32x5 FILLER_136_1238 ();
 b15zdnd11an1n16x5 FILLER_136_1270 ();
 b15zdnd11an1n64x5 FILLER_136_1289 ();
 b15zdnd11an1n64x5 FILLER_136_1353 ();
 b15zdnd11an1n32x5 FILLER_136_1417 ();
 b15zdnd11an1n16x5 FILLER_136_1449 ();
 b15zdnd11an1n08x5 FILLER_136_1465 ();
 b15zdnd11an1n04x5 FILLER_136_1473 ();
 b15zdnd00an1n01x5 FILLER_136_1477 ();
 b15zdnd11an1n08x5 FILLER_136_2265 ();
 b15zdnd00an1n02x5 FILLER_136_2273 ();
 b15zdnd00an1n01x5 FILLER_136_2275 ();
 b15zdnd11an1n64x5 FILLER_137_0 ();
 b15zdnd11an1n64x5 FILLER_137_64 ();
 b15zdnd11an1n64x5 FILLER_137_128 ();
 b15zdnd11an1n64x5 FILLER_137_192 ();
 b15zdnd11an1n64x5 FILLER_137_256 ();
 b15zdnd11an1n64x5 FILLER_137_320 ();
 b15zdnd11an1n64x5 FILLER_137_384 ();
 b15zdnd11an1n64x5 FILLER_137_448 ();
 b15zdnd11an1n64x5 FILLER_137_512 ();
 b15zdnd11an1n64x5 FILLER_137_576 ();
 b15zdnd11an1n64x5 FILLER_137_640 ();
 b15zdnd11an1n64x5 FILLER_137_704 ();
 b15zdnd11an1n64x5 FILLER_137_768 ();
 b15zdnd11an1n64x5 FILLER_137_832 ();
 b15zdnd11an1n64x5 FILLER_137_896 ();
 b15zdnd11an1n64x5 FILLER_137_960 ();
 b15zdnd11an1n64x5 FILLER_137_1024 ();
 b15zdnd11an1n64x5 FILLER_137_1088 ();
 b15zdnd11an1n64x5 FILLER_137_1152 ();
 b15zdnd11an1n64x5 FILLER_137_1216 ();
 b15zdnd11an1n64x5 FILLER_137_1280 ();
 b15zdnd11an1n64x5 FILLER_137_1344 ();
 b15zdnd11an1n64x5 FILLER_137_1408 ();
 b15zdnd11an1n08x5 FILLER_137_1472 ();
 b15zdnd11an1n04x5 FILLER_137_1480 ();
 b15zdnd00an1n02x5 FILLER_137_1484 ();
 b15zdnd11an1n16x5 FILLER_137_2257 ();
 b15zdnd11an1n08x5 FILLER_137_2273 ();
 b15zdnd00an1n02x5 FILLER_137_2281 ();
 b15zdnd00an1n01x5 FILLER_137_2283 ();
 b15zdnd11an1n04x5 FILLER_138_8 ();
 b15zdnd11an1n04x5 FILLER_138_19 ();
 b15zdnd11an1n64x5 FILLER_138_30 ();
 b15zdnd11an1n16x5 FILLER_138_94 ();
 b15zdnd00an1n02x5 FILLER_138_110 ();
 b15zdnd11an1n08x5 FILLER_138_127 ();
 b15zdnd11an1n04x5 FILLER_138_135 ();
 b15zdnd00an1n02x5 FILLER_138_139 ();
 b15zdnd00an1n01x5 FILLER_138_141 ();
 b15zdnd11an1n64x5 FILLER_138_146 ();
 b15zdnd11an1n64x5 FILLER_138_210 ();
 b15zdnd11an1n64x5 FILLER_138_274 ();
 b15zdnd11an1n64x5 FILLER_138_338 ();
 b15zdnd11an1n64x5 FILLER_138_402 ();
 b15zdnd11an1n64x5 FILLER_138_466 ();
 b15zdnd11an1n64x5 FILLER_138_530 ();
 b15zdnd11an1n64x5 FILLER_138_594 ();
 b15zdnd11an1n32x5 FILLER_138_658 ();
 b15zdnd11an1n16x5 FILLER_138_690 ();
 b15zdnd11an1n08x5 FILLER_138_706 ();
 b15zdnd11an1n04x5 FILLER_138_714 ();
 b15zdnd11an1n64x5 FILLER_138_726 ();
 b15zdnd11an1n16x5 FILLER_138_790 ();
 b15zdnd11an1n08x5 FILLER_138_806 ();
 b15zdnd00an1n02x5 FILLER_138_814 ();
 b15zdnd11an1n64x5 FILLER_138_827 ();
 b15zdnd11an1n64x5 FILLER_138_891 ();
 b15zdnd11an1n64x5 FILLER_138_955 ();
 b15zdnd11an1n64x5 FILLER_138_1019 ();
 b15zdnd11an1n64x5 FILLER_138_1083 ();
 b15zdnd11an1n64x5 FILLER_138_1147 ();
 b15zdnd11an1n64x5 FILLER_138_1211 ();
 b15zdnd11an1n64x5 FILLER_138_1275 ();
 b15zdnd11an1n64x5 FILLER_138_1339 ();
 b15zdnd11an1n64x5 FILLER_138_1403 ();
 b15zdnd11an1n08x5 FILLER_138_1467 ();
 b15zdnd00an1n02x5 FILLER_138_1475 ();
 b15zdnd00an1n01x5 FILLER_138_1477 ();
 b15zdnd00an1n02x5 FILLER_138_2265 ();
 b15zdnd00an1n02x5 FILLER_138_2274 ();
 b15zdnd11an1n64x5 FILLER_139_0 ();
 b15zdnd11an1n64x5 FILLER_139_64 ();
 b15zdnd11an1n08x5 FILLER_139_128 ();
 b15zdnd11an1n04x5 FILLER_139_136 ();
 b15zdnd00an1n02x5 FILLER_139_140 ();
 b15zdnd00an1n01x5 FILLER_139_142 ();
 b15zdnd11an1n64x5 FILLER_139_164 ();
 b15zdnd11an1n64x5 FILLER_139_228 ();
 b15zdnd11an1n64x5 FILLER_139_292 ();
 b15zdnd11an1n64x5 FILLER_139_356 ();
 b15zdnd11an1n64x5 FILLER_139_420 ();
 b15zdnd11an1n64x5 FILLER_139_484 ();
 b15zdnd11an1n64x5 FILLER_139_548 ();
 b15zdnd11an1n64x5 FILLER_139_612 ();
 b15zdnd11an1n32x5 FILLER_139_676 ();
 b15zdnd11an1n08x5 FILLER_139_708 ();
 b15zdnd00an1n01x5 FILLER_139_716 ();
 b15zdnd11an1n64x5 FILLER_139_759 ();
 b15zdnd11an1n16x5 FILLER_139_823 ();
 b15zdnd11an1n64x5 FILLER_139_881 ();
 b15zdnd11an1n64x5 FILLER_139_945 ();
 b15zdnd11an1n64x5 FILLER_139_1009 ();
 b15zdnd11an1n64x5 FILLER_139_1073 ();
 b15zdnd11an1n64x5 FILLER_139_1137 ();
 b15zdnd11an1n64x5 FILLER_139_1201 ();
 b15zdnd11an1n64x5 FILLER_139_1265 ();
 b15zdnd11an1n64x5 FILLER_139_1329 ();
 b15zdnd11an1n64x5 FILLER_139_1393 ();
 b15zdnd11an1n16x5 FILLER_139_1457 ();
 b15zdnd11an1n08x5 FILLER_139_1473 ();
 b15zdnd11an1n04x5 FILLER_139_1481 ();
 b15zdnd00an1n01x5 FILLER_139_1485 ();
 b15zdnd11an1n16x5 FILLER_139_2257 ();
 b15zdnd11an1n08x5 FILLER_139_2273 ();
 b15zdnd00an1n02x5 FILLER_139_2281 ();
 b15zdnd00an1n01x5 FILLER_139_2283 ();
 b15zdnd11an1n16x5 FILLER_140_8 ();
 b15zdnd00an1n02x5 FILLER_140_24 ();
 b15zdnd11an1n64x5 FILLER_140_34 ();
 b15zdnd11an1n64x5 FILLER_140_98 ();
 b15zdnd11an1n64x5 FILLER_140_162 ();
 b15zdnd11an1n64x5 FILLER_140_226 ();
 b15zdnd11an1n64x5 FILLER_140_290 ();
 b15zdnd11an1n64x5 FILLER_140_354 ();
 b15zdnd11an1n64x5 FILLER_140_418 ();
 b15zdnd11an1n64x5 FILLER_140_482 ();
 b15zdnd11an1n64x5 FILLER_140_546 ();
 b15zdnd11an1n64x5 FILLER_140_610 ();
 b15zdnd11an1n32x5 FILLER_140_674 ();
 b15zdnd11an1n08x5 FILLER_140_706 ();
 b15zdnd11an1n04x5 FILLER_140_714 ();
 b15zdnd11an1n64x5 FILLER_140_726 ();
 b15zdnd11an1n64x5 FILLER_140_790 ();
 b15zdnd11an1n64x5 FILLER_140_854 ();
 b15zdnd11an1n64x5 FILLER_140_918 ();
 b15zdnd11an1n64x5 FILLER_140_982 ();
 b15zdnd11an1n64x5 FILLER_140_1046 ();
 b15zdnd11an1n64x5 FILLER_140_1110 ();
 b15zdnd11an1n64x5 FILLER_140_1174 ();
 b15zdnd11an1n32x5 FILLER_140_1238 ();
 b15zdnd11an1n08x5 FILLER_140_1270 ();
 b15zdnd00an1n02x5 FILLER_140_1278 ();
 b15zdnd00an1n01x5 FILLER_140_1280 ();
 b15zdnd11an1n64x5 FILLER_140_1323 ();
 b15zdnd11an1n64x5 FILLER_140_1387 ();
 b15zdnd11an1n16x5 FILLER_140_1451 ();
 b15zdnd11an1n08x5 FILLER_140_1467 ();
 b15zdnd00an1n02x5 FILLER_140_1475 ();
 b15zdnd00an1n01x5 FILLER_140_1477 ();
 b15zdnd11an1n08x5 FILLER_140_2265 ();
 b15zdnd00an1n02x5 FILLER_140_2273 ();
 b15zdnd00an1n01x5 FILLER_140_2275 ();
 b15zdnd11an1n32x5 FILLER_141_0 ();
 b15zdnd11an1n04x5 FILLER_141_32 ();
 b15zdnd00an1n02x5 FILLER_141_36 ();
 b15zdnd00an1n01x5 FILLER_141_38 ();
 b15zdnd11an1n64x5 FILLER_141_47 ();
 b15zdnd11an1n64x5 FILLER_141_111 ();
 b15zdnd11an1n64x5 FILLER_141_175 ();
 b15zdnd11an1n16x5 FILLER_141_239 ();
 b15zdnd11an1n08x5 FILLER_141_255 ();
 b15zdnd11an1n04x5 FILLER_141_263 ();
 b15zdnd00an1n02x5 FILLER_141_267 ();
 b15zdnd11an1n64x5 FILLER_141_285 ();
 b15zdnd11an1n32x5 FILLER_141_349 ();
 b15zdnd11an1n16x5 FILLER_141_381 ();
 b15zdnd11an1n08x5 FILLER_141_397 ();
 b15zdnd11an1n04x5 FILLER_141_405 ();
 b15zdnd00an1n02x5 FILLER_141_409 ();
 b15zdnd11an1n64x5 FILLER_141_429 ();
 b15zdnd11an1n64x5 FILLER_141_493 ();
 b15zdnd11an1n64x5 FILLER_141_557 ();
 b15zdnd11an1n64x5 FILLER_141_621 ();
 b15zdnd11an1n64x5 FILLER_141_685 ();
 b15zdnd11an1n64x5 FILLER_141_749 ();
 b15zdnd11an1n64x5 FILLER_141_813 ();
 b15zdnd11an1n64x5 FILLER_141_877 ();
 b15zdnd11an1n64x5 FILLER_141_941 ();
 b15zdnd11an1n64x5 FILLER_141_1005 ();
 b15zdnd11an1n64x5 FILLER_141_1069 ();
 b15zdnd11an1n64x5 FILLER_141_1133 ();
 b15zdnd11an1n64x5 FILLER_141_1197 ();
 b15zdnd11an1n64x5 FILLER_141_1261 ();
 b15zdnd11an1n64x5 FILLER_141_1325 ();
 b15zdnd11an1n64x5 FILLER_141_1389 ();
 b15zdnd11an1n32x5 FILLER_141_1453 ();
 b15zdnd00an1n01x5 FILLER_141_1485 ();
 b15zdnd11an1n16x5 FILLER_141_2257 ();
 b15zdnd11an1n08x5 FILLER_141_2273 ();
 b15zdnd00an1n02x5 FILLER_141_2281 ();
 b15zdnd00an1n01x5 FILLER_141_2283 ();
 b15zdnd11an1n64x5 FILLER_142_8 ();
 b15zdnd11an1n64x5 FILLER_142_72 ();
 b15zdnd11an1n64x5 FILLER_142_136 ();
 b15zdnd11an1n64x5 FILLER_142_200 ();
 b15zdnd11an1n64x5 FILLER_142_264 ();
 b15zdnd11an1n16x5 FILLER_142_328 ();
 b15zdnd00an1n02x5 FILLER_142_344 ();
 b15zdnd00an1n01x5 FILLER_142_346 ();
 b15zdnd11an1n64x5 FILLER_142_389 ();
 b15zdnd11an1n64x5 FILLER_142_453 ();
 b15zdnd11an1n64x5 FILLER_142_517 ();
 b15zdnd11an1n64x5 FILLER_142_581 ();
 b15zdnd11an1n64x5 FILLER_142_645 ();
 b15zdnd11an1n08x5 FILLER_142_709 ();
 b15zdnd00an1n01x5 FILLER_142_717 ();
 b15zdnd11an1n64x5 FILLER_142_726 ();
 b15zdnd11an1n64x5 FILLER_142_790 ();
 b15zdnd11an1n64x5 FILLER_142_854 ();
 b15zdnd11an1n64x5 FILLER_142_918 ();
 b15zdnd11an1n64x5 FILLER_142_982 ();
 b15zdnd11an1n64x5 FILLER_142_1046 ();
 b15zdnd11an1n64x5 FILLER_142_1110 ();
 b15zdnd11an1n64x5 FILLER_142_1174 ();
 b15zdnd11an1n08x5 FILLER_142_1238 ();
 b15zdnd11an1n04x5 FILLER_142_1246 ();
 b15zdnd00an1n01x5 FILLER_142_1250 ();
 b15zdnd11an1n64x5 FILLER_142_1293 ();
 b15zdnd11an1n64x5 FILLER_142_1357 ();
 b15zdnd11an1n32x5 FILLER_142_1421 ();
 b15zdnd11an1n16x5 FILLER_142_1453 ();
 b15zdnd11an1n08x5 FILLER_142_1469 ();
 b15zdnd00an1n01x5 FILLER_142_1477 ();
 b15zdnd11an1n08x5 FILLER_142_2265 ();
 b15zdnd00an1n02x5 FILLER_142_2273 ();
 b15zdnd00an1n01x5 FILLER_142_2275 ();
 b15zdnd11an1n64x5 FILLER_143_0 ();
 b15zdnd11an1n64x5 FILLER_143_64 ();
 b15zdnd11an1n64x5 FILLER_143_128 ();
 b15zdnd11an1n64x5 FILLER_143_192 ();
 b15zdnd11an1n64x5 FILLER_143_256 ();
 b15zdnd11an1n64x5 FILLER_143_320 ();
 b15zdnd11an1n64x5 FILLER_143_384 ();
 b15zdnd11an1n64x5 FILLER_143_448 ();
 b15zdnd11an1n64x5 FILLER_143_512 ();
 b15zdnd11an1n64x5 FILLER_143_576 ();
 b15zdnd11an1n64x5 FILLER_143_640 ();
 b15zdnd11an1n64x5 FILLER_143_704 ();
 b15zdnd11an1n64x5 FILLER_143_768 ();
 b15zdnd11an1n64x5 FILLER_143_832 ();
 b15zdnd11an1n64x5 FILLER_143_896 ();
 b15zdnd11an1n64x5 FILLER_143_960 ();
 b15zdnd11an1n64x5 FILLER_143_1024 ();
 b15zdnd11an1n64x5 FILLER_143_1088 ();
 b15zdnd11an1n64x5 FILLER_143_1152 ();
 b15zdnd11an1n64x5 FILLER_143_1216 ();
 b15zdnd11an1n64x5 FILLER_143_1280 ();
 b15zdnd11an1n64x5 FILLER_143_1344 ();
 b15zdnd11an1n64x5 FILLER_143_1408 ();
 b15zdnd11an1n08x5 FILLER_143_1472 ();
 b15zdnd11an1n04x5 FILLER_143_1480 ();
 b15zdnd00an1n02x5 FILLER_143_1484 ();
 b15zdnd11an1n16x5 FILLER_143_2257 ();
 b15zdnd11an1n08x5 FILLER_143_2273 ();
 b15zdnd00an1n02x5 FILLER_143_2281 ();
 b15zdnd00an1n01x5 FILLER_143_2283 ();
 b15zdnd11an1n64x5 FILLER_144_8 ();
 b15zdnd11an1n64x5 FILLER_144_72 ();
 b15zdnd11an1n64x5 FILLER_144_136 ();
 b15zdnd11an1n64x5 FILLER_144_200 ();
 b15zdnd11an1n64x5 FILLER_144_264 ();
 b15zdnd11an1n64x5 FILLER_144_328 ();
 b15zdnd11an1n64x5 FILLER_144_392 ();
 b15zdnd11an1n64x5 FILLER_144_456 ();
 b15zdnd11an1n64x5 FILLER_144_520 ();
 b15zdnd11an1n64x5 FILLER_144_584 ();
 b15zdnd11an1n64x5 FILLER_144_648 ();
 b15zdnd11an1n04x5 FILLER_144_712 ();
 b15zdnd00an1n02x5 FILLER_144_716 ();
 b15zdnd11an1n64x5 FILLER_144_726 ();
 b15zdnd11an1n64x5 FILLER_144_790 ();
 b15zdnd11an1n64x5 FILLER_144_854 ();
 b15zdnd11an1n64x5 FILLER_144_918 ();
 b15zdnd11an1n64x5 FILLER_144_982 ();
 b15zdnd11an1n64x5 FILLER_144_1046 ();
 b15zdnd11an1n64x5 FILLER_144_1110 ();
 b15zdnd11an1n64x5 FILLER_144_1174 ();
 b15zdnd11an1n64x5 FILLER_144_1238 ();
 b15zdnd11an1n64x5 FILLER_144_1302 ();
 b15zdnd11an1n64x5 FILLER_144_1366 ();
 b15zdnd11an1n32x5 FILLER_144_1430 ();
 b15zdnd11an1n16x5 FILLER_144_1462 ();
 b15zdnd11an1n08x5 FILLER_144_2265 ();
 b15zdnd00an1n02x5 FILLER_144_2273 ();
 b15zdnd00an1n01x5 FILLER_144_2275 ();
 b15zdnd11an1n64x5 FILLER_145_0 ();
 b15zdnd11an1n64x5 FILLER_145_64 ();
 b15zdnd11an1n64x5 FILLER_145_128 ();
 b15zdnd11an1n64x5 FILLER_145_192 ();
 b15zdnd11an1n64x5 FILLER_145_256 ();
 b15zdnd11an1n64x5 FILLER_145_320 ();
 b15zdnd11an1n64x5 FILLER_145_384 ();
 b15zdnd11an1n64x5 FILLER_145_448 ();
 b15zdnd11an1n64x5 FILLER_145_512 ();
 b15zdnd11an1n64x5 FILLER_145_576 ();
 b15zdnd11an1n64x5 FILLER_145_640 ();
 b15zdnd11an1n64x5 FILLER_145_704 ();
 b15zdnd11an1n64x5 FILLER_145_768 ();
 b15zdnd11an1n64x5 FILLER_145_832 ();
 b15zdnd11an1n64x5 FILLER_145_896 ();
 b15zdnd11an1n64x5 FILLER_145_960 ();
 b15zdnd11an1n64x5 FILLER_145_1024 ();
 b15zdnd11an1n64x5 FILLER_145_1088 ();
 b15zdnd11an1n64x5 FILLER_145_1152 ();
 b15zdnd11an1n64x5 FILLER_145_1216 ();
 b15zdnd11an1n64x5 FILLER_145_1280 ();
 b15zdnd11an1n64x5 FILLER_145_1344 ();
 b15zdnd11an1n64x5 FILLER_145_1408 ();
 b15zdnd11an1n08x5 FILLER_145_1472 ();
 b15zdnd11an1n04x5 FILLER_145_1480 ();
 b15zdnd00an1n02x5 FILLER_145_1484 ();
 b15zdnd11an1n16x5 FILLER_145_2257 ();
 b15zdnd11an1n08x5 FILLER_145_2273 ();
 b15zdnd00an1n02x5 FILLER_145_2281 ();
 b15zdnd00an1n01x5 FILLER_145_2283 ();
 b15zdnd11an1n64x5 FILLER_146_8 ();
 b15zdnd11an1n32x5 FILLER_146_72 ();
 b15zdnd00an1n02x5 FILLER_146_104 ();
 b15zdnd11an1n64x5 FILLER_146_109 ();
 b15zdnd11an1n64x5 FILLER_146_173 ();
 b15zdnd11an1n64x5 FILLER_146_279 ();
 b15zdnd11an1n64x5 FILLER_146_343 ();
 b15zdnd11an1n64x5 FILLER_146_407 ();
 b15zdnd11an1n64x5 FILLER_146_471 ();
 b15zdnd11an1n64x5 FILLER_146_535 ();
 b15zdnd11an1n64x5 FILLER_146_599 ();
 b15zdnd11an1n32x5 FILLER_146_663 ();
 b15zdnd11an1n16x5 FILLER_146_695 ();
 b15zdnd11an1n04x5 FILLER_146_711 ();
 b15zdnd00an1n02x5 FILLER_146_715 ();
 b15zdnd00an1n01x5 FILLER_146_717 ();
 b15zdnd11an1n64x5 FILLER_146_726 ();
 b15zdnd11an1n64x5 FILLER_146_790 ();
 b15zdnd11an1n64x5 FILLER_146_854 ();
 b15zdnd11an1n64x5 FILLER_146_918 ();
 b15zdnd11an1n64x5 FILLER_146_982 ();
 b15zdnd11an1n64x5 FILLER_146_1046 ();
 b15zdnd11an1n64x5 FILLER_146_1110 ();
 b15zdnd11an1n64x5 FILLER_146_1174 ();
 b15zdnd11an1n64x5 FILLER_146_1238 ();
 b15zdnd11an1n64x5 FILLER_146_1302 ();
 b15zdnd11an1n64x5 FILLER_146_1366 ();
 b15zdnd11an1n32x5 FILLER_146_1430 ();
 b15zdnd11an1n16x5 FILLER_146_1462 ();
 b15zdnd11an1n08x5 FILLER_146_2265 ();
 b15zdnd00an1n02x5 FILLER_146_2273 ();
 b15zdnd00an1n01x5 FILLER_146_2275 ();
 b15zdnd11an1n64x5 FILLER_147_0 ();
 b15zdnd11an1n64x5 FILLER_147_64 ();
 b15zdnd11an1n64x5 FILLER_147_128 ();
 b15zdnd11an1n64x5 FILLER_147_192 ();
 b15zdnd11an1n64x5 FILLER_147_256 ();
 b15zdnd11an1n64x5 FILLER_147_320 ();
 b15zdnd11an1n64x5 FILLER_147_384 ();
 b15zdnd11an1n64x5 FILLER_147_448 ();
 b15zdnd11an1n64x5 FILLER_147_512 ();
 b15zdnd11an1n64x5 FILLER_147_576 ();
 b15zdnd11an1n64x5 FILLER_147_640 ();
 b15zdnd11an1n64x5 FILLER_147_704 ();
 b15zdnd11an1n64x5 FILLER_147_768 ();
 b15zdnd11an1n64x5 FILLER_147_832 ();
 b15zdnd11an1n64x5 FILLER_147_896 ();
 b15zdnd11an1n64x5 FILLER_147_960 ();
 b15zdnd11an1n64x5 FILLER_147_1024 ();
 b15zdnd11an1n32x5 FILLER_147_1088 ();
 b15zdnd11an1n16x5 FILLER_147_1120 ();
 b15zdnd11an1n08x5 FILLER_147_1136 ();
 b15zdnd00an1n01x5 FILLER_147_1144 ();
 b15zdnd11an1n64x5 FILLER_147_1187 ();
 b15zdnd11an1n64x5 FILLER_147_1251 ();
 b15zdnd11an1n64x5 FILLER_147_1315 ();
 b15zdnd11an1n64x5 FILLER_147_1379 ();
 b15zdnd11an1n32x5 FILLER_147_1443 ();
 b15zdnd11an1n08x5 FILLER_147_1475 ();
 b15zdnd00an1n02x5 FILLER_147_1483 ();
 b15zdnd00an1n01x5 FILLER_147_1485 ();
 b15zdnd11an1n16x5 FILLER_147_2257 ();
 b15zdnd11an1n08x5 FILLER_147_2273 ();
 b15zdnd00an1n02x5 FILLER_147_2281 ();
 b15zdnd00an1n01x5 FILLER_147_2283 ();
 b15zdnd11an1n64x5 FILLER_148_8 ();
 b15zdnd11an1n64x5 FILLER_148_72 ();
 b15zdnd11an1n64x5 FILLER_148_136 ();
 b15zdnd11an1n64x5 FILLER_148_200 ();
 b15zdnd11an1n64x5 FILLER_148_264 ();
 b15zdnd11an1n64x5 FILLER_148_328 ();
 b15zdnd11an1n32x5 FILLER_148_392 ();
 b15zdnd11an1n08x5 FILLER_148_424 ();
 b15zdnd11an1n64x5 FILLER_148_446 ();
 b15zdnd11an1n64x5 FILLER_148_510 ();
 b15zdnd11an1n64x5 FILLER_148_574 ();
 b15zdnd11an1n64x5 FILLER_148_638 ();
 b15zdnd11an1n16x5 FILLER_148_702 ();
 b15zdnd11an1n64x5 FILLER_148_726 ();
 b15zdnd11an1n64x5 FILLER_148_790 ();
 b15zdnd11an1n64x5 FILLER_148_854 ();
 b15zdnd11an1n64x5 FILLER_148_918 ();
 b15zdnd11an1n64x5 FILLER_148_982 ();
 b15zdnd11an1n64x5 FILLER_148_1046 ();
 b15zdnd11an1n64x5 FILLER_148_1110 ();
 b15zdnd11an1n64x5 FILLER_148_1174 ();
 b15zdnd11an1n64x5 FILLER_148_1238 ();
 b15zdnd11an1n64x5 FILLER_148_1302 ();
 b15zdnd11an1n64x5 FILLER_148_1366 ();
 b15zdnd11an1n32x5 FILLER_148_1430 ();
 b15zdnd11an1n16x5 FILLER_148_1462 ();
 b15zdnd00an1n02x5 FILLER_148_2265 ();
 b15zdnd00an1n02x5 FILLER_148_2274 ();
 b15zdnd11an1n64x5 FILLER_149_0 ();
 b15zdnd11an1n64x5 FILLER_149_64 ();
 b15zdnd11an1n64x5 FILLER_149_128 ();
 b15zdnd11an1n64x5 FILLER_149_192 ();
 b15zdnd11an1n64x5 FILLER_149_256 ();
 b15zdnd11an1n64x5 FILLER_149_320 ();
 b15zdnd11an1n64x5 FILLER_149_384 ();
 b15zdnd11an1n64x5 FILLER_149_448 ();
 b15zdnd11an1n64x5 FILLER_149_512 ();
 b15zdnd11an1n64x5 FILLER_149_576 ();
 b15zdnd11an1n64x5 FILLER_149_640 ();
 b15zdnd11an1n64x5 FILLER_149_704 ();
 b15zdnd11an1n64x5 FILLER_149_768 ();
 b15zdnd11an1n64x5 FILLER_149_832 ();
 b15zdnd11an1n64x5 FILLER_149_896 ();
 b15zdnd11an1n64x5 FILLER_149_960 ();
 b15zdnd11an1n64x5 FILLER_149_1024 ();
 b15zdnd11an1n64x5 FILLER_149_1088 ();
 b15zdnd11an1n64x5 FILLER_149_1152 ();
 b15zdnd11an1n32x5 FILLER_149_1216 ();
 b15zdnd11an1n16x5 FILLER_149_1248 ();
 b15zdnd11an1n04x5 FILLER_149_1264 ();
 b15zdnd00an1n02x5 FILLER_149_1268 ();
 b15zdnd00an1n01x5 FILLER_149_1270 ();
 b15zdnd11an1n64x5 FILLER_149_1280 ();
 b15zdnd11an1n64x5 FILLER_149_1344 ();
 b15zdnd11an1n64x5 FILLER_149_1408 ();
 b15zdnd11an1n08x5 FILLER_149_1472 ();
 b15zdnd11an1n04x5 FILLER_149_1480 ();
 b15zdnd00an1n02x5 FILLER_149_1484 ();
 b15zdnd11an1n16x5 FILLER_149_2257 ();
 b15zdnd11an1n08x5 FILLER_149_2273 ();
 b15zdnd00an1n02x5 FILLER_149_2281 ();
 b15zdnd00an1n01x5 FILLER_149_2283 ();
 b15zdnd11an1n64x5 FILLER_150_8 ();
 b15zdnd11an1n64x5 FILLER_150_72 ();
 b15zdnd11an1n64x5 FILLER_150_136 ();
 b15zdnd11an1n64x5 FILLER_150_200 ();
 b15zdnd11an1n64x5 FILLER_150_264 ();
 b15zdnd11an1n64x5 FILLER_150_328 ();
 b15zdnd11an1n64x5 FILLER_150_392 ();
 b15zdnd11an1n64x5 FILLER_150_456 ();
 b15zdnd11an1n64x5 FILLER_150_520 ();
 b15zdnd11an1n64x5 FILLER_150_584 ();
 b15zdnd11an1n64x5 FILLER_150_648 ();
 b15zdnd11an1n04x5 FILLER_150_712 ();
 b15zdnd00an1n02x5 FILLER_150_716 ();
 b15zdnd11an1n64x5 FILLER_150_726 ();
 b15zdnd11an1n64x5 FILLER_150_790 ();
 b15zdnd11an1n64x5 FILLER_150_854 ();
 b15zdnd11an1n64x5 FILLER_150_918 ();
 b15zdnd11an1n64x5 FILLER_150_982 ();
 b15zdnd11an1n64x5 FILLER_150_1046 ();
 b15zdnd11an1n64x5 FILLER_150_1110 ();
 b15zdnd11an1n64x5 FILLER_150_1174 ();
 b15zdnd11an1n64x5 FILLER_150_1238 ();
 b15zdnd11an1n64x5 FILLER_150_1302 ();
 b15zdnd11an1n64x5 FILLER_150_1366 ();
 b15zdnd11an1n32x5 FILLER_150_1430 ();
 b15zdnd11an1n16x5 FILLER_150_1462 ();
 b15zdnd11an1n08x5 FILLER_150_2265 ();
 b15zdnd00an1n02x5 FILLER_150_2273 ();
 b15zdnd00an1n01x5 FILLER_150_2275 ();
 b15zdnd11an1n64x5 FILLER_151_0 ();
 b15zdnd11an1n64x5 FILLER_151_64 ();
 b15zdnd11an1n64x5 FILLER_151_128 ();
 b15zdnd11an1n64x5 FILLER_151_192 ();
 b15zdnd11an1n64x5 FILLER_151_256 ();
 b15zdnd11an1n64x5 FILLER_151_320 ();
 b15zdnd11an1n64x5 FILLER_151_384 ();
 b15zdnd11an1n64x5 FILLER_151_448 ();
 b15zdnd11an1n64x5 FILLER_151_512 ();
 b15zdnd11an1n64x5 FILLER_151_576 ();
 b15zdnd11an1n64x5 FILLER_151_640 ();
 b15zdnd11an1n64x5 FILLER_151_704 ();
 b15zdnd11an1n64x5 FILLER_151_768 ();
 b15zdnd11an1n64x5 FILLER_151_832 ();
 b15zdnd11an1n64x5 FILLER_151_896 ();
 b15zdnd11an1n64x5 FILLER_151_960 ();
 b15zdnd00an1n02x5 FILLER_151_1024 ();
 b15zdnd00an1n01x5 FILLER_151_1026 ();
 b15zdnd11an1n64x5 FILLER_151_1038 ();
 b15zdnd11an1n32x5 FILLER_151_1102 ();
 b15zdnd00an1n02x5 FILLER_151_1134 ();
 b15zdnd00an1n01x5 FILLER_151_1136 ();
 b15zdnd11an1n64x5 FILLER_151_1179 ();
 b15zdnd11an1n64x5 FILLER_151_1243 ();
 b15zdnd11an1n64x5 FILLER_151_1307 ();
 b15zdnd11an1n64x5 FILLER_151_1371 ();
 b15zdnd11an1n32x5 FILLER_151_1435 ();
 b15zdnd11an1n16x5 FILLER_151_1467 ();
 b15zdnd00an1n02x5 FILLER_151_1483 ();
 b15zdnd00an1n01x5 FILLER_151_1485 ();
 b15zdnd11an1n16x5 FILLER_151_2257 ();
 b15zdnd11an1n08x5 FILLER_151_2273 ();
 b15zdnd00an1n02x5 FILLER_151_2281 ();
 b15zdnd00an1n01x5 FILLER_151_2283 ();
 b15zdnd11an1n64x5 FILLER_152_8 ();
 b15zdnd11an1n64x5 FILLER_152_72 ();
 b15zdnd11an1n64x5 FILLER_152_136 ();
 b15zdnd11an1n64x5 FILLER_152_200 ();
 b15zdnd11an1n64x5 FILLER_152_264 ();
 b15zdnd11an1n64x5 FILLER_152_328 ();
 b15zdnd11an1n64x5 FILLER_152_392 ();
 b15zdnd11an1n64x5 FILLER_152_456 ();
 b15zdnd11an1n64x5 FILLER_152_520 ();
 b15zdnd11an1n64x5 FILLER_152_584 ();
 b15zdnd11an1n64x5 FILLER_152_648 ();
 b15zdnd11an1n04x5 FILLER_152_712 ();
 b15zdnd00an1n02x5 FILLER_152_716 ();
 b15zdnd11an1n64x5 FILLER_152_726 ();
 b15zdnd11an1n64x5 FILLER_152_790 ();
 b15zdnd11an1n64x5 FILLER_152_854 ();
 b15zdnd11an1n64x5 FILLER_152_918 ();
 b15zdnd11an1n64x5 FILLER_152_982 ();
 b15zdnd11an1n64x5 FILLER_152_1046 ();
 b15zdnd11an1n64x5 FILLER_152_1110 ();
 b15zdnd11an1n64x5 FILLER_152_1174 ();
 b15zdnd11an1n64x5 FILLER_152_1238 ();
 b15zdnd11an1n64x5 FILLER_152_1302 ();
 b15zdnd11an1n64x5 FILLER_152_1366 ();
 b15zdnd11an1n32x5 FILLER_152_1430 ();
 b15zdnd11an1n16x5 FILLER_152_1462 ();
 b15zdnd11an1n08x5 FILLER_152_2265 ();
 b15zdnd00an1n02x5 FILLER_152_2273 ();
 b15zdnd00an1n01x5 FILLER_152_2275 ();
 b15zdnd11an1n64x5 FILLER_153_0 ();
 b15zdnd11an1n64x5 FILLER_153_64 ();
 b15zdnd11an1n16x5 FILLER_153_128 ();
 b15zdnd11an1n08x5 FILLER_153_144 ();
 b15zdnd00an1n02x5 FILLER_153_152 ();
 b15zdnd11an1n64x5 FILLER_153_196 ();
 b15zdnd11an1n64x5 FILLER_153_260 ();
 b15zdnd11an1n64x5 FILLER_153_324 ();
 b15zdnd11an1n04x5 FILLER_153_388 ();
 b15zdnd00an1n02x5 FILLER_153_392 ();
 b15zdnd00an1n01x5 FILLER_153_394 ();
 b15zdnd11an1n64x5 FILLER_153_426 ();
 b15zdnd11an1n64x5 FILLER_153_490 ();
 b15zdnd11an1n64x5 FILLER_153_554 ();
 b15zdnd11an1n64x5 FILLER_153_618 ();
 b15zdnd11an1n64x5 FILLER_153_682 ();
 b15zdnd11an1n64x5 FILLER_153_746 ();
 b15zdnd11an1n64x5 FILLER_153_810 ();
 b15zdnd11an1n64x5 FILLER_153_874 ();
 b15zdnd11an1n64x5 FILLER_153_938 ();
 b15zdnd11an1n64x5 FILLER_153_1002 ();
 b15zdnd11an1n64x5 FILLER_153_1066 ();
 b15zdnd11an1n64x5 FILLER_153_1130 ();
 b15zdnd11an1n64x5 FILLER_153_1194 ();
 b15zdnd11an1n64x5 FILLER_153_1258 ();
 b15zdnd11an1n64x5 FILLER_153_1322 ();
 b15zdnd11an1n16x5 FILLER_153_1386 ();
 b15zdnd11an1n08x5 FILLER_153_1402 ();
 b15zdnd00an1n02x5 FILLER_153_1410 ();
 b15zdnd00an1n01x5 FILLER_153_1412 ();
 b15zdnd11an1n16x5 FILLER_153_1455 ();
 b15zdnd11an1n08x5 FILLER_153_1471 ();
 b15zdnd11an1n04x5 FILLER_153_1479 ();
 b15zdnd00an1n02x5 FILLER_153_1483 ();
 b15zdnd00an1n01x5 FILLER_153_1485 ();
 b15zdnd11an1n16x5 FILLER_153_2257 ();
 b15zdnd11an1n08x5 FILLER_153_2273 ();
 b15zdnd00an1n02x5 FILLER_153_2281 ();
 b15zdnd00an1n01x5 FILLER_153_2283 ();
 b15zdnd00an1n02x5 FILLER_154_8 ();
 b15zdnd11an1n64x5 FILLER_154_21 ();
 b15zdnd11an1n64x5 FILLER_154_85 ();
 b15zdnd11an1n32x5 FILLER_154_149 ();
 b15zdnd11an1n16x5 FILLER_154_181 ();
 b15zdnd11an1n08x5 FILLER_154_197 ();
 b15zdnd11an1n04x5 FILLER_154_205 ();
 b15zdnd11an1n64x5 FILLER_154_229 ();
 b15zdnd11an1n64x5 FILLER_154_293 ();
 b15zdnd11an1n64x5 FILLER_154_357 ();
 b15zdnd11an1n64x5 FILLER_154_421 ();
 b15zdnd11an1n64x5 FILLER_154_485 ();
 b15zdnd11an1n64x5 FILLER_154_549 ();
 b15zdnd11an1n64x5 FILLER_154_613 ();
 b15zdnd11an1n32x5 FILLER_154_677 ();
 b15zdnd11an1n08x5 FILLER_154_709 ();
 b15zdnd00an1n01x5 FILLER_154_717 ();
 b15zdnd11an1n64x5 FILLER_154_726 ();
 b15zdnd11an1n64x5 FILLER_154_790 ();
 b15zdnd11an1n64x5 FILLER_154_854 ();
 b15zdnd11an1n32x5 FILLER_154_918 ();
 b15zdnd11an1n08x5 FILLER_154_950 ();
 b15zdnd00an1n02x5 FILLER_154_958 ();
 b15zdnd11an1n64x5 FILLER_154_969 ();
 b15zdnd11an1n64x5 FILLER_154_1033 ();
 b15zdnd11an1n64x5 FILLER_154_1097 ();
 b15zdnd11an1n16x5 FILLER_154_1161 ();
 b15zdnd11an1n04x5 FILLER_154_1177 ();
 b15zdnd11an1n64x5 FILLER_154_1223 ();
 b15zdnd11an1n64x5 FILLER_154_1287 ();
 b15zdnd11an1n64x5 FILLER_154_1351 ();
 b15zdnd11an1n32x5 FILLER_154_1415 ();
 b15zdnd11an1n16x5 FILLER_154_1447 ();
 b15zdnd11an1n08x5 FILLER_154_1463 ();
 b15zdnd11an1n04x5 FILLER_154_1471 ();
 b15zdnd00an1n02x5 FILLER_154_1475 ();
 b15zdnd00an1n01x5 FILLER_154_1477 ();
 b15zdnd11an1n08x5 FILLER_154_2265 ();
 b15zdnd00an1n02x5 FILLER_154_2273 ();
 b15zdnd00an1n01x5 FILLER_154_2275 ();
 b15zdnd11an1n64x5 FILLER_155_0 ();
 b15zdnd11an1n64x5 FILLER_155_64 ();
 b15zdnd11an1n32x5 FILLER_155_128 ();
 b15zdnd11an1n16x5 FILLER_155_160 ();
 b15zdnd11an1n08x5 FILLER_155_176 ();
 b15zdnd11an1n04x5 FILLER_155_184 ();
 b15zdnd00an1n01x5 FILLER_155_188 ();
 b15zdnd11an1n64x5 FILLER_155_211 ();
 b15zdnd11an1n64x5 FILLER_155_275 ();
 b15zdnd11an1n64x5 FILLER_155_339 ();
 b15zdnd11an1n16x5 FILLER_155_403 ();
 b15zdnd11an1n04x5 FILLER_155_419 ();
 b15zdnd00an1n02x5 FILLER_155_423 ();
 b15zdnd00an1n01x5 FILLER_155_425 ();
 b15zdnd11an1n64x5 FILLER_155_468 ();
 b15zdnd11an1n64x5 FILLER_155_532 ();
 b15zdnd11an1n64x5 FILLER_155_596 ();
 b15zdnd11an1n64x5 FILLER_155_660 ();
 b15zdnd11an1n64x5 FILLER_155_724 ();
 b15zdnd11an1n64x5 FILLER_155_788 ();
 b15zdnd11an1n64x5 FILLER_155_852 ();
 b15zdnd11an1n64x5 FILLER_155_916 ();
 b15zdnd11an1n64x5 FILLER_155_980 ();
 b15zdnd11an1n64x5 FILLER_155_1044 ();
 b15zdnd11an1n64x5 FILLER_155_1108 ();
 b15zdnd11an1n64x5 FILLER_155_1172 ();
 b15zdnd11an1n64x5 FILLER_155_1236 ();
 b15zdnd11an1n64x5 FILLER_155_1300 ();
 b15zdnd11an1n32x5 FILLER_155_1364 ();
 b15zdnd11an1n08x5 FILLER_155_1396 ();
 b15zdnd11an1n04x5 FILLER_155_1404 ();
 b15zdnd00an1n02x5 FILLER_155_1408 ();
 b15zdnd00an1n01x5 FILLER_155_1410 ();
 b15zdnd11an1n04x5 FILLER_155_1453 ();
 b15zdnd11an1n08x5 FILLER_155_1471 ();
 b15zdnd11an1n04x5 FILLER_155_1479 ();
 b15zdnd00an1n02x5 FILLER_155_1483 ();
 b15zdnd00an1n01x5 FILLER_155_1485 ();
 b15zdnd11an1n16x5 FILLER_155_2257 ();
 b15zdnd11an1n08x5 FILLER_155_2273 ();
 b15zdnd00an1n02x5 FILLER_155_2281 ();
 b15zdnd00an1n01x5 FILLER_155_2283 ();
 b15zdnd11an1n64x5 FILLER_156_8 ();
 b15zdnd11an1n64x5 FILLER_156_72 ();
 b15zdnd11an1n64x5 FILLER_156_136 ();
 b15zdnd11an1n32x5 FILLER_156_200 ();
 b15zdnd11an1n08x5 FILLER_156_232 ();
 b15zdnd11an1n04x5 FILLER_156_240 ();
 b15zdnd11an1n64x5 FILLER_156_255 ();
 b15zdnd11an1n64x5 FILLER_156_319 ();
 b15zdnd11an1n64x5 FILLER_156_383 ();
 b15zdnd11an1n64x5 FILLER_156_447 ();
 b15zdnd11an1n64x5 FILLER_156_511 ();
 b15zdnd11an1n64x5 FILLER_156_575 ();
 b15zdnd11an1n64x5 FILLER_156_639 ();
 b15zdnd11an1n08x5 FILLER_156_703 ();
 b15zdnd11an1n04x5 FILLER_156_711 ();
 b15zdnd00an1n02x5 FILLER_156_715 ();
 b15zdnd00an1n01x5 FILLER_156_717 ();
 b15zdnd11an1n64x5 FILLER_156_726 ();
 b15zdnd11an1n64x5 FILLER_156_790 ();
 b15zdnd11an1n64x5 FILLER_156_854 ();
 b15zdnd11an1n64x5 FILLER_156_918 ();
 b15zdnd11an1n64x5 FILLER_156_982 ();
 b15zdnd11an1n64x5 FILLER_156_1046 ();
 b15zdnd11an1n32x5 FILLER_156_1110 ();
 b15zdnd11an1n04x5 FILLER_156_1142 ();
 b15zdnd11an1n64x5 FILLER_156_1154 ();
 b15zdnd11an1n16x5 FILLER_156_1218 ();
 b15zdnd11an1n04x5 FILLER_156_1234 ();
 b15zdnd11an1n64x5 FILLER_156_1280 ();
 b15zdnd11an1n64x5 FILLER_156_1344 ();
 b15zdnd11an1n64x5 FILLER_156_1408 ();
 b15zdnd11an1n04x5 FILLER_156_1472 ();
 b15zdnd00an1n02x5 FILLER_156_1476 ();
 b15zdnd11an1n08x5 FILLER_156_2265 ();
 b15zdnd00an1n02x5 FILLER_156_2273 ();
 b15zdnd00an1n01x5 FILLER_156_2275 ();
 b15zdnd11an1n64x5 FILLER_157_0 ();
 b15zdnd11an1n64x5 FILLER_157_64 ();
 b15zdnd11an1n64x5 FILLER_157_128 ();
 b15zdnd11an1n64x5 FILLER_157_192 ();
 b15zdnd11an1n64x5 FILLER_157_256 ();
 b15zdnd11an1n64x5 FILLER_157_320 ();
 b15zdnd11an1n64x5 FILLER_157_384 ();
 b15zdnd11an1n64x5 FILLER_157_448 ();
 b15zdnd11an1n64x5 FILLER_157_512 ();
 b15zdnd11an1n64x5 FILLER_157_576 ();
 b15zdnd11an1n64x5 FILLER_157_640 ();
 b15zdnd11an1n64x5 FILLER_157_704 ();
 b15zdnd11an1n64x5 FILLER_157_768 ();
 b15zdnd11an1n64x5 FILLER_157_832 ();
 b15zdnd11an1n64x5 FILLER_157_896 ();
 b15zdnd11an1n64x5 FILLER_157_960 ();
 b15zdnd11an1n64x5 FILLER_157_1024 ();
 b15zdnd11an1n64x5 FILLER_157_1088 ();
 b15zdnd11an1n64x5 FILLER_157_1152 ();
 b15zdnd11an1n32x5 FILLER_157_1216 ();
 b15zdnd11an1n04x5 FILLER_157_1248 ();
 b15zdnd00an1n02x5 FILLER_157_1252 ();
 b15zdnd00an1n01x5 FILLER_157_1254 ();
 b15zdnd11an1n64x5 FILLER_157_1297 ();
 b15zdnd11an1n64x5 FILLER_157_1361 ();
 b15zdnd11an1n32x5 FILLER_157_1425 ();
 b15zdnd11an1n16x5 FILLER_157_1457 ();
 b15zdnd11an1n08x5 FILLER_157_1473 ();
 b15zdnd11an1n04x5 FILLER_157_1481 ();
 b15zdnd00an1n01x5 FILLER_157_1485 ();
 b15zdnd11an1n16x5 FILLER_157_2257 ();
 b15zdnd11an1n08x5 FILLER_157_2273 ();
 b15zdnd00an1n02x5 FILLER_157_2281 ();
 b15zdnd00an1n01x5 FILLER_157_2283 ();
 b15zdnd11an1n64x5 FILLER_158_8 ();
 b15zdnd11an1n64x5 FILLER_158_72 ();
 b15zdnd11an1n64x5 FILLER_158_136 ();
 b15zdnd11an1n64x5 FILLER_158_200 ();
 b15zdnd11an1n64x5 FILLER_158_264 ();
 b15zdnd11an1n64x5 FILLER_158_328 ();
 b15zdnd11an1n64x5 FILLER_158_392 ();
 b15zdnd11an1n64x5 FILLER_158_456 ();
 b15zdnd11an1n64x5 FILLER_158_520 ();
 b15zdnd11an1n64x5 FILLER_158_584 ();
 b15zdnd11an1n64x5 FILLER_158_648 ();
 b15zdnd11an1n04x5 FILLER_158_712 ();
 b15zdnd00an1n02x5 FILLER_158_716 ();
 b15zdnd11an1n64x5 FILLER_158_726 ();
 b15zdnd11an1n64x5 FILLER_158_790 ();
 b15zdnd11an1n64x5 FILLER_158_854 ();
 b15zdnd11an1n64x5 FILLER_158_918 ();
 b15zdnd11an1n64x5 FILLER_158_982 ();
 b15zdnd11an1n64x5 FILLER_158_1046 ();
 b15zdnd11an1n64x5 FILLER_158_1110 ();
 b15zdnd11an1n64x5 FILLER_158_1174 ();
 b15zdnd11an1n08x5 FILLER_158_1238 ();
 b15zdnd11an1n64x5 FILLER_158_1288 ();
 b15zdnd11an1n64x5 FILLER_158_1352 ();
 b15zdnd11an1n32x5 FILLER_158_1416 ();
 b15zdnd11an1n16x5 FILLER_158_1448 ();
 b15zdnd11an1n08x5 FILLER_158_1464 ();
 b15zdnd11an1n04x5 FILLER_158_1472 ();
 b15zdnd00an1n02x5 FILLER_158_1476 ();
 b15zdnd11an1n08x5 FILLER_158_2265 ();
 b15zdnd00an1n02x5 FILLER_158_2273 ();
 b15zdnd00an1n01x5 FILLER_158_2275 ();
 b15zdnd11an1n64x5 FILLER_159_0 ();
 b15zdnd11an1n64x5 FILLER_159_64 ();
 b15zdnd11an1n64x5 FILLER_159_128 ();
 b15zdnd11an1n64x5 FILLER_159_192 ();
 b15zdnd11an1n64x5 FILLER_159_256 ();
 b15zdnd11an1n64x5 FILLER_159_320 ();
 b15zdnd11an1n64x5 FILLER_159_384 ();
 b15zdnd11an1n64x5 FILLER_159_448 ();
 b15zdnd11an1n64x5 FILLER_159_512 ();
 b15zdnd11an1n64x5 FILLER_159_576 ();
 b15zdnd11an1n64x5 FILLER_159_640 ();
 b15zdnd11an1n64x5 FILLER_159_704 ();
 b15zdnd11an1n64x5 FILLER_159_768 ();
 b15zdnd11an1n64x5 FILLER_159_832 ();
 b15zdnd11an1n64x5 FILLER_159_896 ();
 b15zdnd11an1n64x5 FILLER_159_960 ();
 b15zdnd11an1n64x5 FILLER_159_1024 ();
 b15zdnd11an1n64x5 FILLER_159_1088 ();
 b15zdnd11an1n64x5 FILLER_159_1152 ();
 b15zdnd11an1n64x5 FILLER_159_1216 ();
 b15zdnd11an1n64x5 FILLER_159_1280 ();
 b15zdnd11an1n64x5 FILLER_159_1344 ();
 b15zdnd11an1n64x5 FILLER_159_1408 ();
 b15zdnd11an1n08x5 FILLER_159_1472 ();
 b15zdnd11an1n04x5 FILLER_159_1480 ();
 b15zdnd00an1n02x5 FILLER_159_1484 ();
 b15zdnd11an1n08x5 FILLER_159_2257 ();
 b15zdnd11an1n08x5 FILLER_159_2272 ();
 b15zdnd11an1n04x5 FILLER_159_2280 ();
 b15zdnd11an1n64x5 FILLER_160_8 ();
 b15zdnd11an1n64x5 FILLER_160_72 ();
 b15zdnd11an1n64x5 FILLER_160_136 ();
 b15zdnd11an1n64x5 FILLER_160_200 ();
 b15zdnd11an1n64x5 FILLER_160_264 ();
 b15zdnd11an1n64x5 FILLER_160_328 ();
 b15zdnd11an1n32x5 FILLER_160_392 ();
 b15zdnd11an1n08x5 FILLER_160_424 ();
 b15zdnd11an1n08x5 FILLER_160_448 ();
 b15zdnd11an1n04x5 FILLER_160_456 ();
 b15zdnd00an1n01x5 FILLER_160_460 ();
 b15zdnd11an1n64x5 FILLER_160_477 ();
 b15zdnd11an1n64x5 FILLER_160_541 ();
 b15zdnd11an1n64x5 FILLER_160_605 ();
 b15zdnd11an1n32x5 FILLER_160_669 ();
 b15zdnd11an1n16x5 FILLER_160_701 ();
 b15zdnd00an1n01x5 FILLER_160_717 ();
 b15zdnd11an1n64x5 FILLER_160_726 ();
 b15zdnd11an1n64x5 FILLER_160_790 ();
 b15zdnd11an1n64x5 FILLER_160_854 ();
 b15zdnd11an1n64x5 FILLER_160_918 ();
 b15zdnd11an1n64x5 FILLER_160_982 ();
 b15zdnd11an1n64x5 FILLER_160_1046 ();
 b15zdnd11an1n64x5 FILLER_160_1110 ();
 b15zdnd11an1n64x5 FILLER_160_1174 ();
 b15zdnd11an1n64x5 FILLER_160_1238 ();
 b15zdnd11an1n64x5 FILLER_160_1302 ();
 b15zdnd11an1n64x5 FILLER_160_1366 ();
 b15zdnd11an1n32x5 FILLER_160_1430 ();
 b15zdnd11an1n16x5 FILLER_160_1462 ();
 b15zdnd11an1n08x5 FILLER_160_2265 ();
 b15zdnd00an1n02x5 FILLER_160_2273 ();
 b15zdnd00an1n01x5 FILLER_160_2275 ();
 b15zdnd11an1n64x5 FILLER_161_0 ();
 b15zdnd11an1n64x5 FILLER_161_64 ();
 b15zdnd11an1n64x5 FILLER_161_128 ();
 b15zdnd11an1n64x5 FILLER_161_192 ();
 b15zdnd11an1n64x5 FILLER_161_256 ();
 b15zdnd11an1n64x5 FILLER_161_320 ();
 b15zdnd11an1n64x5 FILLER_161_384 ();
 b15zdnd11an1n64x5 FILLER_161_448 ();
 b15zdnd11an1n64x5 FILLER_161_512 ();
 b15zdnd11an1n64x5 FILLER_161_576 ();
 b15zdnd11an1n64x5 FILLER_161_640 ();
 b15zdnd11an1n64x5 FILLER_161_704 ();
 b15zdnd11an1n64x5 FILLER_161_768 ();
 b15zdnd11an1n64x5 FILLER_161_832 ();
 b15zdnd11an1n64x5 FILLER_161_896 ();
 b15zdnd11an1n64x5 FILLER_161_960 ();
 b15zdnd11an1n64x5 FILLER_161_1024 ();
 b15zdnd11an1n64x5 FILLER_161_1088 ();
 b15zdnd00an1n02x5 FILLER_161_1152 ();
 b15zdnd11an1n64x5 FILLER_161_1157 ();
 b15zdnd11an1n64x5 FILLER_161_1221 ();
 b15zdnd11an1n32x5 FILLER_161_1285 ();
 b15zdnd11an1n04x5 FILLER_161_1317 ();
 b15zdnd00an1n02x5 FILLER_161_1321 ();
 b15zdnd11an1n04x5 FILLER_161_1326 ();
 b15zdnd11an1n64x5 FILLER_161_1333 ();
 b15zdnd11an1n64x5 FILLER_161_1397 ();
 b15zdnd11an1n16x5 FILLER_161_1461 ();
 b15zdnd11an1n08x5 FILLER_161_1477 ();
 b15zdnd00an1n01x5 FILLER_161_1485 ();
 b15zdnd11an1n16x5 FILLER_161_2257 ();
 b15zdnd11an1n08x5 FILLER_161_2273 ();
 b15zdnd00an1n02x5 FILLER_161_2281 ();
 b15zdnd00an1n01x5 FILLER_161_2283 ();
 b15zdnd11an1n16x5 FILLER_162_8 ();
 b15zdnd00an1n02x5 FILLER_162_24 ();
 b15zdnd00an1n01x5 FILLER_162_26 ();
 b15zdnd11an1n04x5 FILLER_162_31 ();
 b15zdnd11an1n64x5 FILLER_162_43 ();
 b15zdnd11an1n64x5 FILLER_162_107 ();
 b15zdnd11an1n64x5 FILLER_162_171 ();
 b15zdnd11an1n64x5 FILLER_162_235 ();
 b15zdnd11an1n64x5 FILLER_162_299 ();
 b15zdnd11an1n64x5 FILLER_162_363 ();
 b15zdnd11an1n08x5 FILLER_162_427 ();
 b15zdnd11an1n04x5 FILLER_162_435 ();
 b15zdnd00an1n02x5 FILLER_162_439 ();
 b15zdnd00an1n01x5 FILLER_162_441 ();
 b15zdnd11an1n08x5 FILLER_162_456 ();
 b15zdnd00an1n01x5 FILLER_162_464 ();
 b15zdnd11an1n64x5 FILLER_162_475 ();
 b15zdnd11an1n64x5 FILLER_162_539 ();
 b15zdnd11an1n64x5 FILLER_162_603 ();
 b15zdnd11an1n32x5 FILLER_162_667 ();
 b15zdnd11an1n16x5 FILLER_162_699 ();
 b15zdnd00an1n02x5 FILLER_162_715 ();
 b15zdnd00an1n01x5 FILLER_162_717 ();
 b15zdnd11an1n64x5 FILLER_162_726 ();
 b15zdnd11an1n64x5 FILLER_162_790 ();
 b15zdnd11an1n64x5 FILLER_162_854 ();
 b15zdnd11an1n32x5 FILLER_162_918 ();
 b15zdnd11an1n08x5 FILLER_162_950 ();
 b15zdnd11an1n04x5 FILLER_162_958 ();
 b15zdnd11an1n64x5 FILLER_162_972 ();
 b15zdnd11an1n64x5 FILLER_162_1036 ();
 b15zdnd11an1n32x5 FILLER_162_1100 ();
 b15zdnd11an1n16x5 FILLER_162_1132 ();
 b15zdnd11an1n04x5 FILLER_162_1148 ();
 b15zdnd00an1n01x5 FILLER_162_1152 ();
 b15zdnd11an1n64x5 FILLER_162_1178 ();
 b15zdnd11an1n32x5 FILLER_162_1242 ();
 b15zdnd11an1n16x5 FILLER_162_1274 ();
 b15zdnd11an1n08x5 FILLER_162_1290 ();
 b15zdnd11an1n04x5 FILLER_162_1298 ();
 b15zdnd00an1n01x5 FILLER_162_1302 ();
 b15zdnd11an1n64x5 FILLER_162_1355 ();
 b15zdnd11an1n32x5 FILLER_162_1419 ();
 b15zdnd11an1n16x5 FILLER_162_1451 ();
 b15zdnd11an1n08x5 FILLER_162_1467 ();
 b15zdnd00an1n02x5 FILLER_162_1475 ();
 b15zdnd00an1n01x5 FILLER_162_1477 ();
 b15zdnd11an1n08x5 FILLER_162_2265 ();
 b15zdnd00an1n02x5 FILLER_162_2273 ();
 b15zdnd00an1n01x5 FILLER_162_2275 ();
 b15zdnd11an1n08x5 FILLER_163_0 ();
 b15zdnd00an1n01x5 FILLER_163_8 ();
 b15zdnd11an1n64x5 FILLER_163_51 ();
 b15zdnd11an1n64x5 FILLER_163_115 ();
 b15zdnd11an1n64x5 FILLER_163_179 ();
 b15zdnd11an1n64x5 FILLER_163_243 ();
 b15zdnd11an1n64x5 FILLER_163_307 ();
 b15zdnd11an1n64x5 FILLER_163_371 ();
 b15zdnd11an1n32x5 FILLER_163_435 ();
 b15zdnd11an1n04x5 FILLER_163_467 ();
 b15zdnd00an1n01x5 FILLER_163_471 ();
 b15zdnd11an1n64x5 FILLER_163_484 ();
 b15zdnd11an1n64x5 FILLER_163_548 ();
 b15zdnd11an1n64x5 FILLER_163_612 ();
 b15zdnd11an1n64x5 FILLER_163_676 ();
 b15zdnd11an1n64x5 FILLER_163_740 ();
 b15zdnd11an1n64x5 FILLER_163_804 ();
 b15zdnd11an1n64x5 FILLER_163_868 ();
 b15zdnd11an1n64x5 FILLER_163_932 ();
 b15zdnd11an1n64x5 FILLER_163_996 ();
 b15zdnd11an1n64x5 FILLER_163_1060 ();
 b15zdnd11an1n32x5 FILLER_163_1124 ();
 b15zdnd00an1n02x5 FILLER_163_1156 ();
 b15zdnd11an1n64x5 FILLER_163_1161 ();
 b15zdnd11an1n64x5 FILLER_163_1225 ();
 b15zdnd11an1n32x5 FILLER_163_1289 ();
 b15zdnd11an1n08x5 FILLER_163_1321 ();
 b15zdnd11an1n04x5 FILLER_163_1329 ();
 b15zdnd11an1n64x5 FILLER_163_1336 ();
 b15zdnd11an1n64x5 FILLER_163_1400 ();
 b15zdnd11an1n16x5 FILLER_163_1464 ();
 b15zdnd11an1n04x5 FILLER_163_1480 ();
 b15zdnd00an1n02x5 FILLER_163_1484 ();
 b15zdnd11an1n04x5 FILLER_163_2257 ();
 b15zdnd00an1n02x5 FILLER_163_2261 ();
 b15zdnd00an1n01x5 FILLER_163_2263 ();
 b15zdnd11an1n08x5 FILLER_163_2271 ();
 b15zdnd11an1n04x5 FILLER_163_2279 ();
 b15zdnd00an1n01x5 FILLER_163_2283 ();
 b15zdnd11an1n64x5 FILLER_164_8 ();
 b15zdnd11an1n64x5 FILLER_164_72 ();
 b15zdnd11an1n64x5 FILLER_164_136 ();
 b15zdnd11an1n64x5 FILLER_164_200 ();
 b15zdnd11an1n64x5 FILLER_164_264 ();
 b15zdnd11an1n64x5 FILLER_164_328 ();
 b15zdnd11an1n08x5 FILLER_164_392 ();
 b15zdnd11an1n04x5 FILLER_164_400 ();
 b15zdnd00an1n02x5 FILLER_164_404 ();
 b15zdnd00an1n01x5 FILLER_164_406 ();
 b15zdnd11an1n16x5 FILLER_164_416 ();
 b15zdnd11an1n08x5 FILLER_164_432 ();
 b15zdnd00an1n01x5 FILLER_164_440 ();
 b15zdnd11an1n64x5 FILLER_164_453 ();
 b15zdnd11an1n64x5 FILLER_164_517 ();
 b15zdnd11an1n64x5 FILLER_164_581 ();
 b15zdnd11an1n64x5 FILLER_164_645 ();
 b15zdnd11an1n08x5 FILLER_164_709 ();
 b15zdnd00an1n01x5 FILLER_164_717 ();
 b15zdnd11an1n64x5 FILLER_164_726 ();
 b15zdnd11an1n64x5 FILLER_164_790 ();
 b15zdnd11an1n64x5 FILLER_164_854 ();
 b15zdnd11an1n64x5 FILLER_164_918 ();
 b15zdnd11an1n64x5 FILLER_164_982 ();
 b15zdnd11an1n16x5 FILLER_164_1046 ();
 b15zdnd11an1n04x5 FILLER_164_1062 ();
 b15zdnd00an1n01x5 FILLER_164_1066 ();
 b15zdnd11an1n64x5 FILLER_164_1075 ();
 b15zdnd11an1n32x5 FILLER_164_1139 ();
 b15zdnd11an1n16x5 FILLER_164_1171 ();
 b15zdnd11an1n16x5 FILLER_164_1229 ();
 b15zdnd11an1n08x5 FILLER_164_1245 ();
 b15zdnd11an1n04x5 FILLER_164_1253 ();
 b15zdnd00an1n02x5 FILLER_164_1257 ();
 b15zdnd11an1n64x5 FILLER_164_1301 ();
 b15zdnd11an1n64x5 FILLER_164_1365 ();
 b15zdnd11an1n32x5 FILLER_164_1429 ();
 b15zdnd11an1n16x5 FILLER_164_1461 ();
 b15zdnd00an1n01x5 FILLER_164_1477 ();
 b15zdnd00an1n02x5 FILLER_164_2265 ();
 b15zdnd00an1n02x5 FILLER_164_2274 ();
 b15zdnd11an1n64x5 FILLER_165_0 ();
 b15zdnd11an1n64x5 FILLER_165_64 ();
 b15zdnd11an1n64x5 FILLER_165_128 ();
 b15zdnd11an1n64x5 FILLER_165_192 ();
 b15zdnd11an1n64x5 FILLER_165_256 ();
 b15zdnd11an1n64x5 FILLER_165_320 ();
 b15zdnd11an1n64x5 FILLER_165_384 ();
 b15zdnd11an1n64x5 FILLER_165_448 ();
 b15zdnd11an1n64x5 FILLER_165_512 ();
 b15zdnd11an1n64x5 FILLER_165_576 ();
 b15zdnd11an1n64x5 FILLER_165_640 ();
 b15zdnd11an1n64x5 FILLER_165_704 ();
 b15zdnd11an1n64x5 FILLER_165_768 ();
 b15zdnd11an1n64x5 FILLER_165_832 ();
 b15zdnd11an1n32x5 FILLER_165_896 ();
 b15zdnd11an1n16x5 FILLER_165_928 ();
 b15zdnd11an1n08x5 FILLER_165_944 ();
 b15zdnd00an1n01x5 FILLER_165_952 ();
 b15zdnd11an1n08x5 FILLER_165_993 ();
 b15zdnd00an1n01x5 FILLER_165_1001 ();
 b15zdnd11an1n64x5 FILLER_165_1005 ();
 b15zdnd11an1n64x5 FILLER_165_1111 ();
 b15zdnd11an1n64x5 FILLER_165_1175 ();
 b15zdnd11an1n16x5 FILLER_165_1239 ();
 b15zdnd11an1n08x5 FILLER_165_1258 ();
 b15zdnd00an1n02x5 FILLER_165_1266 ();
 b15zdnd11an1n64x5 FILLER_165_1271 ();
 b15zdnd11an1n32x5 FILLER_165_1335 ();
 b15zdnd11an1n16x5 FILLER_165_1367 ();
 b15zdnd00an1n02x5 FILLER_165_1383 ();
 b15zdnd00an1n01x5 FILLER_165_1385 ();
 b15zdnd11an1n32x5 FILLER_165_1428 ();
 b15zdnd11an1n16x5 FILLER_165_1460 ();
 b15zdnd11an1n08x5 FILLER_165_1476 ();
 b15zdnd00an1n02x5 FILLER_165_1484 ();
 b15zdnd11an1n16x5 FILLER_165_2257 ();
 b15zdnd11an1n08x5 FILLER_165_2273 ();
 b15zdnd00an1n02x5 FILLER_165_2281 ();
 b15zdnd00an1n01x5 FILLER_165_2283 ();
 b15zdnd11an1n64x5 FILLER_166_8 ();
 b15zdnd11an1n64x5 FILLER_166_72 ();
 b15zdnd11an1n64x5 FILLER_166_136 ();
 b15zdnd11an1n64x5 FILLER_166_200 ();
 b15zdnd11an1n64x5 FILLER_166_264 ();
 b15zdnd11an1n64x5 FILLER_166_328 ();
 b15zdnd11an1n32x5 FILLER_166_392 ();
 b15zdnd00an1n01x5 FILLER_166_424 ();
 b15zdnd11an1n64x5 FILLER_166_437 ();
 b15zdnd11an1n64x5 FILLER_166_501 ();
 b15zdnd11an1n64x5 FILLER_166_565 ();
 b15zdnd11an1n64x5 FILLER_166_629 ();
 b15zdnd11an1n16x5 FILLER_166_693 ();
 b15zdnd11an1n08x5 FILLER_166_709 ();
 b15zdnd00an1n01x5 FILLER_166_717 ();
 b15zdnd11an1n64x5 FILLER_166_726 ();
 b15zdnd11an1n64x5 FILLER_166_790 ();
 b15zdnd11an1n64x5 FILLER_166_854 ();
 b15zdnd11an1n32x5 FILLER_166_918 ();
 b15zdnd11an1n16x5 FILLER_166_950 ();
 b15zdnd11an1n08x5 FILLER_166_966 ();
 b15zdnd00an1n01x5 FILLER_166_974 ();
 b15zdnd11an1n32x5 FILLER_166_1017 ();
 b15zdnd11an1n04x5 FILLER_166_1049 ();
 b15zdnd00an1n01x5 FILLER_166_1053 ();
 b15zdnd11an1n08x5 FILLER_166_1062 ();
 b15zdnd00an1n01x5 FILLER_166_1070 ();
 b15zdnd11an1n64x5 FILLER_166_1079 ();
 b15zdnd11an1n64x5 FILLER_166_1143 ();
 b15zdnd11an1n16x5 FILLER_166_1207 ();
 b15zdnd11an1n08x5 FILLER_166_1223 ();
 b15zdnd00an1n01x5 FILLER_166_1231 ();
 b15zdnd11an1n64x5 FILLER_166_1284 ();
 b15zdnd11an1n64x5 FILLER_166_1348 ();
 b15zdnd11an1n64x5 FILLER_166_1412 ();
 b15zdnd00an1n02x5 FILLER_166_1476 ();
 b15zdnd11an1n08x5 FILLER_166_2265 ();
 b15zdnd00an1n02x5 FILLER_166_2273 ();
 b15zdnd00an1n01x5 FILLER_166_2275 ();
 b15zdnd11an1n64x5 FILLER_167_0 ();
 b15zdnd11an1n64x5 FILLER_167_64 ();
 b15zdnd11an1n64x5 FILLER_167_128 ();
 b15zdnd11an1n64x5 FILLER_167_192 ();
 b15zdnd11an1n64x5 FILLER_167_256 ();
 b15zdnd11an1n64x5 FILLER_167_320 ();
 b15zdnd11an1n32x5 FILLER_167_384 ();
 b15zdnd11an1n08x5 FILLER_167_416 ();
 b15zdnd00an1n02x5 FILLER_167_424 ();
 b15zdnd11an1n64x5 FILLER_167_450 ();
 b15zdnd11an1n64x5 FILLER_167_514 ();
 b15zdnd11an1n64x5 FILLER_167_578 ();
 b15zdnd11an1n64x5 FILLER_167_642 ();
 b15zdnd11an1n32x5 FILLER_167_706 ();
 b15zdnd11an1n16x5 FILLER_167_738 ();
 b15zdnd00an1n01x5 FILLER_167_754 ();
 b15zdnd11an1n64x5 FILLER_167_797 ();
 b15zdnd11an1n64x5 FILLER_167_861 ();
 b15zdnd11an1n08x5 FILLER_167_925 ();
 b15zdnd00an1n02x5 FILLER_167_933 ();
 b15zdnd11an1n16x5 FILLER_167_938 ();
 b15zdnd11an1n08x5 FILLER_167_954 ();
 b15zdnd11an1n04x5 FILLER_167_962 ();
 b15zdnd11an1n04x5 FILLER_167_1006 ();
 b15zdnd11an1n32x5 FILLER_167_1013 ();
 b15zdnd11an1n08x5 FILLER_167_1045 ();
 b15zdnd11an1n04x5 FILLER_167_1053 ();
 b15zdnd00an1n01x5 FILLER_167_1057 ();
 b15zdnd11an1n64x5 FILLER_167_1061 ();
 b15zdnd00an1n02x5 FILLER_167_1125 ();
 b15zdnd00an1n01x5 FILLER_167_1127 ();
 b15zdnd11an1n16x5 FILLER_167_1131 ();
 b15zdnd11an1n04x5 FILLER_167_1147 ();
 b15zdnd00an1n02x5 FILLER_167_1151 ();
 b15zdnd11an1n32x5 FILLER_167_1195 ();
 b15zdnd11an1n16x5 FILLER_167_1227 ();
 b15zdnd11an1n08x5 FILLER_167_1243 ();
 b15zdnd11an1n04x5 FILLER_167_1251 ();
 b15zdnd00an1n02x5 FILLER_167_1255 ();
 b15zdnd00an1n01x5 FILLER_167_1257 ();
 b15zdnd11an1n64x5 FILLER_167_1261 ();
 b15zdnd11an1n64x5 FILLER_167_1325 ();
 b15zdnd11an1n64x5 FILLER_167_1389 ();
 b15zdnd11an1n32x5 FILLER_167_1453 ();
 b15zdnd00an1n01x5 FILLER_167_1485 ();
 b15zdnd11an1n16x5 FILLER_167_2257 ();
 b15zdnd11an1n08x5 FILLER_167_2273 ();
 b15zdnd00an1n02x5 FILLER_167_2281 ();
 b15zdnd00an1n01x5 FILLER_167_2283 ();
 b15zdnd11an1n64x5 FILLER_168_8 ();
 b15zdnd11an1n64x5 FILLER_168_72 ();
 b15zdnd11an1n64x5 FILLER_168_136 ();
 b15zdnd11an1n64x5 FILLER_168_200 ();
 b15zdnd11an1n64x5 FILLER_168_264 ();
 b15zdnd11an1n64x5 FILLER_168_328 ();
 b15zdnd11an1n32x5 FILLER_168_392 ();
 b15zdnd11an1n16x5 FILLER_168_424 ();
 b15zdnd00an1n02x5 FILLER_168_440 ();
 b15zdnd11an1n08x5 FILLER_168_446 ();
 b15zdnd00an1n01x5 FILLER_168_454 ();
 b15zdnd11an1n64x5 FILLER_168_466 ();
 b15zdnd11an1n64x5 FILLER_168_530 ();
 b15zdnd11an1n64x5 FILLER_168_594 ();
 b15zdnd11an1n32x5 FILLER_168_658 ();
 b15zdnd11an1n16x5 FILLER_168_690 ();
 b15zdnd11an1n08x5 FILLER_168_706 ();
 b15zdnd11an1n04x5 FILLER_168_714 ();
 b15zdnd11an1n64x5 FILLER_168_726 ();
 b15zdnd11an1n64x5 FILLER_168_790 ();
 b15zdnd11an1n32x5 FILLER_168_854 ();
 b15zdnd11an1n16x5 FILLER_168_886 ();
 b15zdnd11an1n04x5 FILLER_168_902 ();
 b15zdnd00an1n02x5 FILLER_168_906 ();
 b15zdnd11an1n16x5 FILLER_168_960 ();
 b15zdnd11an1n08x5 FILLER_168_976 ();
 b15zdnd11an1n04x5 FILLER_168_987 ();
 b15zdnd11an1n32x5 FILLER_168_994 ();
 b15zdnd11an1n16x5 FILLER_168_1026 ();
 b15zdnd11an1n08x5 FILLER_168_1042 ();
 b15zdnd11an1n04x5 FILLER_168_1050 ();
 b15zdnd11an1n32x5 FILLER_168_1089 ();
 b15zdnd00an1n02x5 FILLER_168_1121 ();
 b15zdnd00an1n01x5 FILLER_168_1123 ();
 b15zdnd11an1n64x5 FILLER_168_1159 ();
 b15zdnd11an1n64x5 FILLER_168_1223 ();
 b15zdnd11an1n64x5 FILLER_168_1287 ();
 b15zdnd11an1n16x5 FILLER_168_1351 ();
 b15zdnd11an1n04x5 FILLER_168_1367 ();
 b15zdnd00an1n02x5 FILLER_168_1371 ();
 b15zdnd11an1n32x5 FILLER_168_1415 ();
 b15zdnd11an1n16x5 FILLER_168_1447 ();
 b15zdnd11an1n08x5 FILLER_168_1463 ();
 b15zdnd11an1n04x5 FILLER_168_1471 ();
 b15zdnd00an1n02x5 FILLER_168_1475 ();
 b15zdnd00an1n01x5 FILLER_168_1477 ();
 b15zdnd11an1n08x5 FILLER_168_2265 ();
 b15zdnd00an1n02x5 FILLER_168_2273 ();
 b15zdnd00an1n01x5 FILLER_168_2275 ();
 b15zdnd11an1n64x5 FILLER_169_0 ();
 b15zdnd11an1n64x5 FILLER_169_64 ();
 b15zdnd11an1n64x5 FILLER_169_128 ();
 b15zdnd11an1n64x5 FILLER_169_192 ();
 b15zdnd11an1n64x5 FILLER_169_256 ();
 b15zdnd11an1n64x5 FILLER_169_320 ();
 b15zdnd11an1n64x5 FILLER_169_384 ();
 b15zdnd11an1n64x5 FILLER_169_448 ();
 b15zdnd11an1n64x5 FILLER_169_512 ();
 b15zdnd11an1n64x5 FILLER_169_576 ();
 b15zdnd11an1n64x5 FILLER_169_640 ();
 b15zdnd11an1n64x5 FILLER_169_704 ();
 b15zdnd11an1n64x5 FILLER_169_768 ();
 b15zdnd11an1n64x5 FILLER_169_832 ();
 b15zdnd11an1n16x5 FILLER_169_896 ();
 b15zdnd11an1n08x5 FILLER_169_912 ();
 b15zdnd00an1n02x5 FILLER_169_920 ();
 b15zdnd00an1n01x5 FILLER_169_922 ();
 b15zdnd11an1n04x5 FILLER_169_926 ();
 b15zdnd11an1n64x5 FILLER_169_933 ();
 b15zdnd11an1n16x5 FILLER_169_997 ();
 b15zdnd11an1n08x5 FILLER_169_1013 ();
 b15zdnd11an1n04x5 FILLER_169_1021 ();
 b15zdnd11an1n08x5 FILLER_169_1041 ();
 b15zdnd11an1n04x5 FILLER_169_1049 ();
 b15zdnd11an1n64x5 FILLER_169_1056 ();
 b15zdnd11an1n04x5 FILLER_169_1120 ();
 b15zdnd11an1n64x5 FILLER_169_1127 ();
 b15zdnd11an1n64x5 FILLER_169_1191 ();
 b15zdnd11an1n64x5 FILLER_169_1255 ();
 b15zdnd11an1n64x5 FILLER_169_1319 ();
 b15zdnd11an1n64x5 FILLER_169_1383 ();
 b15zdnd11an1n32x5 FILLER_169_1447 ();
 b15zdnd11an1n04x5 FILLER_169_1479 ();
 b15zdnd00an1n02x5 FILLER_169_1483 ();
 b15zdnd00an1n01x5 FILLER_169_1485 ();
 b15zdnd11an1n16x5 FILLER_169_2257 ();
 b15zdnd11an1n08x5 FILLER_169_2273 ();
 b15zdnd00an1n02x5 FILLER_169_2281 ();
 b15zdnd00an1n01x5 FILLER_169_2283 ();
 b15zdnd11an1n64x5 FILLER_170_8 ();
 b15zdnd11an1n64x5 FILLER_170_72 ();
 b15zdnd11an1n64x5 FILLER_170_136 ();
 b15zdnd11an1n64x5 FILLER_170_200 ();
 b15zdnd11an1n64x5 FILLER_170_264 ();
 b15zdnd11an1n64x5 FILLER_170_328 ();
 b15zdnd11an1n64x5 FILLER_170_392 ();
 b15zdnd11an1n16x5 FILLER_170_456 ();
 b15zdnd11an1n04x5 FILLER_170_472 ();
 b15zdnd00an1n02x5 FILLER_170_476 ();
 b15zdnd11an1n64x5 FILLER_170_494 ();
 b15zdnd11an1n64x5 FILLER_170_558 ();
 b15zdnd11an1n32x5 FILLER_170_622 ();
 b15zdnd11an1n08x5 FILLER_170_654 ();
 b15zdnd11an1n16x5 FILLER_170_702 ();
 b15zdnd11an1n64x5 FILLER_170_726 ();
 b15zdnd11an1n64x5 FILLER_170_790 ();
 b15zdnd11an1n64x5 FILLER_170_854 ();
 b15zdnd11an1n64x5 FILLER_170_918 ();
 b15zdnd11an1n64x5 FILLER_170_982 ();
 b15zdnd11an1n64x5 FILLER_170_1046 ();
 b15zdnd11an1n64x5 FILLER_170_1110 ();
 b15zdnd11an1n16x5 FILLER_170_1174 ();
 b15zdnd00an1n02x5 FILLER_170_1190 ();
 b15zdnd00an1n01x5 FILLER_170_1192 ();
 b15zdnd11an1n64x5 FILLER_170_1235 ();
 b15zdnd11an1n64x5 FILLER_170_1299 ();
 b15zdnd11an1n64x5 FILLER_170_1363 ();
 b15zdnd11an1n32x5 FILLER_170_1427 ();
 b15zdnd11an1n16x5 FILLER_170_1459 ();
 b15zdnd00an1n02x5 FILLER_170_1475 ();
 b15zdnd00an1n01x5 FILLER_170_1477 ();
 b15zdnd11an1n08x5 FILLER_170_2265 ();
 b15zdnd00an1n02x5 FILLER_170_2273 ();
 b15zdnd00an1n01x5 FILLER_170_2275 ();
 b15zdnd11an1n64x5 FILLER_171_0 ();
 b15zdnd11an1n64x5 FILLER_171_64 ();
 b15zdnd11an1n64x5 FILLER_171_128 ();
 b15zdnd11an1n64x5 FILLER_171_192 ();
 b15zdnd11an1n16x5 FILLER_171_256 ();
 b15zdnd11an1n08x5 FILLER_171_272 ();
 b15zdnd11an1n64x5 FILLER_171_292 ();
 b15zdnd11an1n64x5 FILLER_171_356 ();
 b15zdnd11an1n64x5 FILLER_171_420 ();
 b15zdnd11an1n64x5 FILLER_171_484 ();
 b15zdnd11an1n64x5 FILLER_171_548 ();
 b15zdnd11an1n64x5 FILLER_171_612 ();
 b15zdnd11an1n16x5 FILLER_171_676 ();
 b15zdnd11an1n04x5 FILLER_171_692 ();
 b15zdnd00an1n02x5 FILLER_171_696 ();
 b15zdnd00an1n01x5 FILLER_171_698 ();
 b15zdnd11an1n64x5 FILLER_171_702 ();
 b15zdnd11an1n64x5 FILLER_171_766 ();
 b15zdnd11an1n64x5 FILLER_171_830 ();
 b15zdnd11an1n16x5 FILLER_171_894 ();
 b15zdnd11an1n04x5 FILLER_171_910 ();
 b15zdnd11an1n64x5 FILLER_171_956 ();
 b15zdnd11an1n64x5 FILLER_171_1020 ();
 b15zdnd11an1n64x5 FILLER_171_1084 ();
 b15zdnd11an1n32x5 FILLER_171_1148 ();
 b15zdnd11an1n16x5 FILLER_171_1180 ();
 b15zdnd11an1n08x5 FILLER_171_1196 ();
 b15zdnd00an1n02x5 FILLER_171_1204 ();
 b15zdnd11an1n64x5 FILLER_171_1229 ();
 b15zdnd11an1n64x5 FILLER_171_1293 ();
 b15zdnd11an1n64x5 FILLER_171_1357 ();
 b15zdnd11an1n64x5 FILLER_171_1421 ();
 b15zdnd00an1n01x5 FILLER_171_1485 ();
 b15zdnd11an1n16x5 FILLER_171_2257 ();
 b15zdnd11an1n08x5 FILLER_171_2273 ();
 b15zdnd00an1n02x5 FILLER_171_2281 ();
 b15zdnd00an1n01x5 FILLER_171_2283 ();
 b15zdnd11an1n64x5 FILLER_172_8 ();
 b15zdnd11an1n64x5 FILLER_172_72 ();
 b15zdnd11an1n64x5 FILLER_172_136 ();
 b15zdnd11an1n64x5 FILLER_172_200 ();
 b15zdnd11an1n64x5 FILLER_172_264 ();
 b15zdnd11an1n64x5 FILLER_172_328 ();
 b15zdnd11an1n64x5 FILLER_172_392 ();
 b15zdnd11an1n64x5 FILLER_172_456 ();
 b15zdnd11an1n64x5 FILLER_172_520 ();
 b15zdnd11an1n64x5 FILLER_172_584 ();
 b15zdnd11an1n64x5 FILLER_172_648 ();
 b15zdnd11an1n04x5 FILLER_172_712 ();
 b15zdnd00an1n02x5 FILLER_172_716 ();
 b15zdnd11an1n64x5 FILLER_172_726 ();
 b15zdnd11an1n64x5 FILLER_172_790 ();
 b15zdnd11an1n64x5 FILLER_172_854 ();
 b15zdnd11an1n64x5 FILLER_172_918 ();
 b15zdnd11an1n64x5 FILLER_172_982 ();
 b15zdnd11an1n08x5 FILLER_172_1046 ();
 b15zdnd11an1n04x5 FILLER_172_1054 ();
 b15zdnd00an1n02x5 FILLER_172_1058 ();
 b15zdnd11an1n64x5 FILLER_172_1076 ();
 b15zdnd11an1n64x5 FILLER_172_1140 ();
 b15zdnd11an1n64x5 FILLER_172_1204 ();
 b15zdnd11an1n64x5 FILLER_172_1268 ();
 b15zdnd11an1n64x5 FILLER_172_1332 ();
 b15zdnd11an1n64x5 FILLER_172_1396 ();
 b15zdnd11an1n16x5 FILLER_172_1460 ();
 b15zdnd00an1n02x5 FILLER_172_1476 ();
 b15zdnd11an1n08x5 FILLER_172_2265 ();
 b15zdnd00an1n02x5 FILLER_172_2273 ();
 b15zdnd00an1n01x5 FILLER_172_2275 ();
 b15zdnd11an1n64x5 FILLER_173_0 ();
 b15zdnd11an1n64x5 FILLER_173_64 ();
 b15zdnd11an1n64x5 FILLER_173_128 ();
 b15zdnd11an1n64x5 FILLER_173_192 ();
 b15zdnd11an1n64x5 FILLER_173_256 ();
 b15zdnd11an1n64x5 FILLER_173_320 ();
 b15zdnd11an1n32x5 FILLER_173_384 ();
 b15zdnd11an1n08x5 FILLER_173_416 ();
 b15zdnd00an1n02x5 FILLER_173_424 ();
 b15zdnd11an1n64x5 FILLER_173_431 ();
 b15zdnd11an1n64x5 FILLER_173_495 ();
 b15zdnd11an1n64x5 FILLER_173_559 ();
 b15zdnd11an1n32x5 FILLER_173_623 ();
 b15zdnd00an1n02x5 FILLER_173_655 ();
 b15zdnd00an1n01x5 FILLER_173_657 ();
 b15zdnd11an1n04x5 FILLER_173_698 ();
 b15zdnd11an1n16x5 FILLER_173_705 ();
 b15zdnd11an1n04x5 FILLER_173_721 ();
 b15zdnd00an1n02x5 FILLER_173_725 ();
 b15zdnd11an1n64x5 FILLER_173_730 ();
 b15zdnd11an1n64x5 FILLER_173_794 ();
 b15zdnd11an1n32x5 FILLER_173_858 ();
 b15zdnd11an1n16x5 FILLER_173_890 ();
 b15zdnd11an1n08x5 FILLER_173_906 ();
 b15zdnd00an1n02x5 FILLER_173_914 ();
 b15zdnd00an1n01x5 FILLER_173_916 ();
 b15zdnd11an1n64x5 FILLER_173_925 ();
 b15zdnd11an1n64x5 FILLER_173_989 ();
 b15zdnd11an1n64x5 FILLER_173_1053 ();
 b15zdnd11an1n64x5 FILLER_173_1117 ();
 b15zdnd11an1n32x5 FILLER_173_1181 ();
 b15zdnd11an1n08x5 FILLER_173_1213 ();
 b15zdnd00an1n02x5 FILLER_173_1221 ();
 b15zdnd00an1n01x5 FILLER_173_1223 ();
 b15zdnd11an1n64x5 FILLER_173_1244 ();
 b15zdnd11an1n64x5 FILLER_173_1308 ();
 b15zdnd11an1n64x5 FILLER_173_1372 ();
 b15zdnd11an1n32x5 FILLER_173_1436 ();
 b15zdnd11an1n16x5 FILLER_173_1468 ();
 b15zdnd00an1n02x5 FILLER_173_1484 ();
 b15zdnd11an1n16x5 FILLER_173_2257 ();
 b15zdnd11an1n08x5 FILLER_173_2273 ();
 b15zdnd00an1n02x5 FILLER_173_2281 ();
 b15zdnd00an1n01x5 FILLER_173_2283 ();
 b15zdnd11an1n64x5 FILLER_174_8 ();
 b15zdnd11an1n64x5 FILLER_174_72 ();
 b15zdnd11an1n64x5 FILLER_174_136 ();
 b15zdnd11an1n64x5 FILLER_174_200 ();
 b15zdnd11an1n64x5 FILLER_174_264 ();
 b15zdnd11an1n64x5 FILLER_174_328 ();
 b15zdnd11an1n64x5 FILLER_174_392 ();
 b15zdnd11an1n64x5 FILLER_174_456 ();
 b15zdnd11an1n64x5 FILLER_174_520 ();
 b15zdnd11an1n64x5 FILLER_174_584 ();
 b15zdnd11an1n16x5 FILLER_174_648 ();
 b15zdnd11an1n04x5 FILLER_174_704 ();
 b15zdnd11an1n04x5 FILLER_174_711 ();
 b15zdnd00an1n02x5 FILLER_174_715 ();
 b15zdnd00an1n01x5 FILLER_174_717 ();
 b15zdnd11an1n32x5 FILLER_174_726 ();
 b15zdnd11an1n16x5 FILLER_174_758 ();
 b15zdnd11an1n32x5 FILLER_174_816 ();
 b15zdnd11an1n08x5 FILLER_174_848 ();
 b15zdnd11an1n04x5 FILLER_174_856 ();
 b15zdnd00an1n02x5 FILLER_174_860 ();
 b15zdnd11an1n64x5 FILLER_174_904 ();
 b15zdnd11an1n64x5 FILLER_174_968 ();
 b15zdnd11an1n64x5 FILLER_174_1032 ();
 b15zdnd11an1n64x5 FILLER_174_1096 ();
 b15zdnd11an1n64x5 FILLER_174_1160 ();
 b15zdnd11an1n16x5 FILLER_174_1224 ();
 b15zdnd11an1n64x5 FILLER_174_1266 ();
 b15zdnd11an1n64x5 FILLER_174_1330 ();
 b15zdnd11an1n64x5 FILLER_174_1394 ();
 b15zdnd11an1n16x5 FILLER_174_1458 ();
 b15zdnd11an1n04x5 FILLER_174_1474 ();
 b15zdnd11an1n08x5 FILLER_174_2265 ();
 b15zdnd00an1n02x5 FILLER_174_2273 ();
 b15zdnd00an1n01x5 FILLER_174_2275 ();
 b15zdnd11an1n64x5 FILLER_175_0 ();
 b15zdnd11an1n64x5 FILLER_175_64 ();
 b15zdnd11an1n64x5 FILLER_175_128 ();
 b15zdnd11an1n64x5 FILLER_175_192 ();
 b15zdnd11an1n64x5 FILLER_175_256 ();
 b15zdnd11an1n64x5 FILLER_175_320 ();
 b15zdnd11an1n64x5 FILLER_175_384 ();
 b15zdnd11an1n64x5 FILLER_175_448 ();
 b15zdnd11an1n64x5 FILLER_175_512 ();
 b15zdnd11an1n64x5 FILLER_175_576 ();
 b15zdnd11an1n16x5 FILLER_175_640 ();
 b15zdnd11an1n08x5 FILLER_175_656 ();
 b15zdnd11an1n04x5 FILLER_175_664 ();
 b15zdnd11an1n04x5 FILLER_175_708 ();
 b15zdnd11an1n04x5 FILLER_175_715 ();
 b15zdnd11an1n64x5 FILLER_175_722 ();
 b15zdnd11an1n64x5 FILLER_175_786 ();
 b15zdnd11an1n64x5 FILLER_175_850 ();
 b15zdnd11an1n64x5 FILLER_175_914 ();
 b15zdnd11an1n64x5 FILLER_175_978 ();
 b15zdnd11an1n64x5 FILLER_175_1042 ();
 b15zdnd11an1n32x5 FILLER_175_1106 ();
 b15zdnd11an1n04x5 FILLER_175_1138 ();
 b15zdnd00an1n02x5 FILLER_175_1142 ();
 b15zdnd00an1n01x5 FILLER_175_1144 ();
 b15zdnd11an1n32x5 FILLER_175_1153 ();
 b15zdnd11an1n16x5 FILLER_175_1185 ();
 b15zdnd00an1n02x5 FILLER_175_1201 ();
 b15zdnd00an1n01x5 FILLER_175_1203 ();
 b15zdnd11an1n64x5 FILLER_175_1220 ();
 b15zdnd11an1n64x5 FILLER_175_1284 ();
 b15zdnd11an1n64x5 FILLER_175_1348 ();
 b15zdnd11an1n64x5 FILLER_175_1412 ();
 b15zdnd11an1n08x5 FILLER_175_1476 ();
 b15zdnd00an1n02x5 FILLER_175_1484 ();
 b15zdnd11an1n08x5 FILLER_175_2257 ();
 b15zdnd11an1n04x5 FILLER_175_2265 ();
 b15zdnd00an1n01x5 FILLER_175_2269 ();
 b15zdnd11an1n08x5 FILLER_175_2274 ();
 b15zdnd00an1n02x5 FILLER_175_2282 ();
 b15zdnd11an1n64x5 FILLER_176_8 ();
 b15zdnd11an1n64x5 FILLER_176_72 ();
 b15zdnd11an1n64x5 FILLER_176_136 ();
 b15zdnd11an1n64x5 FILLER_176_200 ();
 b15zdnd11an1n64x5 FILLER_176_264 ();
 b15zdnd11an1n64x5 FILLER_176_328 ();
 b15zdnd11an1n32x5 FILLER_176_392 ();
 b15zdnd11an1n04x5 FILLER_176_424 ();
 b15zdnd00an1n01x5 FILLER_176_428 ();
 b15zdnd11an1n64x5 FILLER_176_435 ();
 b15zdnd11an1n64x5 FILLER_176_499 ();
 b15zdnd11an1n64x5 FILLER_176_563 ();
 b15zdnd11an1n64x5 FILLER_176_627 ();
 b15zdnd11an1n04x5 FILLER_176_691 ();
 b15zdnd00an1n01x5 FILLER_176_695 ();
 b15zdnd11an1n04x5 FILLER_176_699 ();
 b15zdnd00an1n01x5 FILLER_176_703 ();
 b15zdnd11an1n08x5 FILLER_176_707 ();
 b15zdnd00an1n02x5 FILLER_176_715 ();
 b15zdnd00an1n01x5 FILLER_176_717 ();
 b15zdnd11an1n64x5 FILLER_176_726 ();
 b15zdnd11an1n64x5 FILLER_176_790 ();
 b15zdnd11an1n64x5 FILLER_176_854 ();
 b15zdnd11an1n64x5 FILLER_176_918 ();
 b15zdnd11an1n64x5 FILLER_176_982 ();
 b15zdnd11an1n64x5 FILLER_176_1046 ();
 b15zdnd11an1n64x5 FILLER_176_1110 ();
 b15zdnd11an1n08x5 FILLER_176_1174 ();
 b15zdnd11an1n64x5 FILLER_176_1198 ();
 b15zdnd11an1n64x5 FILLER_176_1262 ();
 b15zdnd11an1n64x5 FILLER_176_1326 ();
 b15zdnd11an1n64x5 FILLER_176_1390 ();
 b15zdnd11an1n16x5 FILLER_176_1454 ();
 b15zdnd11an1n08x5 FILLER_176_1470 ();
 b15zdnd11an1n08x5 FILLER_176_2265 ();
 b15zdnd00an1n02x5 FILLER_176_2273 ();
 b15zdnd00an1n01x5 FILLER_176_2275 ();
 b15zdnd11an1n64x5 FILLER_177_0 ();
 b15zdnd11an1n64x5 FILLER_177_64 ();
 b15zdnd11an1n64x5 FILLER_177_128 ();
 b15zdnd11an1n64x5 FILLER_177_192 ();
 b15zdnd11an1n64x5 FILLER_177_256 ();
 b15zdnd11an1n64x5 FILLER_177_320 ();
 b15zdnd11an1n64x5 FILLER_177_384 ();
 b15zdnd11an1n64x5 FILLER_177_448 ();
 b15zdnd11an1n64x5 FILLER_177_512 ();
 b15zdnd11an1n64x5 FILLER_177_576 ();
 b15zdnd11an1n64x5 FILLER_177_640 ();
 b15zdnd11an1n64x5 FILLER_177_704 ();
 b15zdnd11an1n64x5 FILLER_177_768 ();
 b15zdnd11an1n64x5 FILLER_177_832 ();
 b15zdnd11an1n64x5 FILLER_177_896 ();
 b15zdnd11an1n64x5 FILLER_177_960 ();
 b15zdnd11an1n64x5 FILLER_177_1024 ();
 b15zdnd11an1n64x5 FILLER_177_1088 ();
 b15zdnd11an1n64x5 FILLER_177_1152 ();
 b15zdnd11an1n64x5 FILLER_177_1216 ();
 b15zdnd11an1n32x5 FILLER_177_1280 ();
 b15zdnd11an1n16x5 FILLER_177_1312 ();
 b15zdnd11an1n04x5 FILLER_177_1328 ();
 b15zdnd11an1n64x5 FILLER_177_1348 ();
 b15zdnd11an1n64x5 FILLER_177_1412 ();
 b15zdnd11an1n08x5 FILLER_177_1476 ();
 b15zdnd00an1n02x5 FILLER_177_1484 ();
 b15zdnd11an1n16x5 FILLER_177_2257 ();
 b15zdnd11an1n08x5 FILLER_177_2273 ();
 b15zdnd00an1n02x5 FILLER_177_2281 ();
 b15zdnd00an1n01x5 FILLER_177_2283 ();
 b15zdnd11an1n64x5 FILLER_178_8 ();
 b15zdnd11an1n64x5 FILLER_178_72 ();
 b15zdnd11an1n64x5 FILLER_178_136 ();
 b15zdnd11an1n64x5 FILLER_178_200 ();
 b15zdnd11an1n64x5 FILLER_178_264 ();
 b15zdnd11an1n64x5 FILLER_178_328 ();
 b15zdnd11an1n32x5 FILLER_178_392 ();
 b15zdnd11an1n08x5 FILLER_178_424 ();
 b15zdnd11an1n04x5 FILLER_178_432 ();
 b15zdnd11an1n64x5 FILLER_178_463 ();
 b15zdnd11an1n64x5 FILLER_178_527 ();
 b15zdnd11an1n64x5 FILLER_178_591 ();
 b15zdnd11an1n32x5 FILLER_178_655 ();
 b15zdnd11an1n16x5 FILLER_178_687 ();
 b15zdnd11an1n08x5 FILLER_178_703 ();
 b15zdnd11an1n04x5 FILLER_178_711 ();
 b15zdnd00an1n02x5 FILLER_178_715 ();
 b15zdnd00an1n01x5 FILLER_178_717 ();
 b15zdnd11an1n64x5 FILLER_178_726 ();
 b15zdnd11an1n64x5 FILLER_178_790 ();
 b15zdnd11an1n64x5 FILLER_178_854 ();
 b15zdnd11an1n64x5 FILLER_178_918 ();
 b15zdnd11an1n64x5 FILLER_178_982 ();
 b15zdnd11an1n64x5 FILLER_178_1046 ();
 b15zdnd11an1n64x5 FILLER_178_1110 ();
 b15zdnd11an1n64x5 FILLER_178_1174 ();
 b15zdnd11an1n64x5 FILLER_178_1238 ();
 b15zdnd11an1n64x5 FILLER_178_1302 ();
 b15zdnd11an1n64x5 FILLER_178_1366 ();
 b15zdnd11an1n32x5 FILLER_178_1430 ();
 b15zdnd11an1n16x5 FILLER_178_1462 ();
 b15zdnd11an1n08x5 FILLER_178_2265 ();
 b15zdnd00an1n02x5 FILLER_178_2273 ();
 b15zdnd00an1n01x5 FILLER_178_2275 ();
 b15zdnd11an1n64x5 FILLER_179_0 ();
 b15zdnd11an1n64x5 FILLER_179_64 ();
 b15zdnd11an1n64x5 FILLER_179_128 ();
 b15zdnd11an1n64x5 FILLER_179_192 ();
 b15zdnd11an1n64x5 FILLER_179_256 ();
 b15zdnd11an1n64x5 FILLER_179_320 ();
 b15zdnd11an1n64x5 FILLER_179_384 ();
 b15zdnd11an1n64x5 FILLER_179_448 ();
 b15zdnd11an1n64x5 FILLER_179_512 ();
 b15zdnd11an1n64x5 FILLER_179_576 ();
 b15zdnd11an1n64x5 FILLER_179_640 ();
 b15zdnd11an1n64x5 FILLER_179_704 ();
 b15zdnd11an1n64x5 FILLER_179_768 ();
 b15zdnd11an1n64x5 FILLER_179_832 ();
 b15zdnd11an1n64x5 FILLER_179_896 ();
 b15zdnd11an1n64x5 FILLER_179_960 ();
 b15zdnd11an1n64x5 FILLER_179_1024 ();
 b15zdnd11an1n64x5 FILLER_179_1088 ();
 b15zdnd11an1n64x5 FILLER_179_1152 ();
 b15zdnd11an1n64x5 FILLER_179_1216 ();
 b15zdnd11an1n64x5 FILLER_179_1280 ();
 b15zdnd11an1n64x5 FILLER_179_1344 ();
 b15zdnd11an1n64x5 FILLER_179_1408 ();
 b15zdnd11an1n08x5 FILLER_179_1472 ();
 b15zdnd11an1n04x5 FILLER_179_1480 ();
 b15zdnd00an1n02x5 FILLER_179_1484 ();
 b15zdnd11an1n16x5 FILLER_179_2257 ();
 b15zdnd11an1n08x5 FILLER_179_2273 ();
 b15zdnd00an1n02x5 FILLER_179_2281 ();
 b15zdnd00an1n01x5 FILLER_179_2283 ();
 b15zdnd11an1n64x5 FILLER_180_8 ();
 b15zdnd11an1n64x5 FILLER_180_72 ();
 b15zdnd11an1n64x5 FILLER_180_136 ();
 b15zdnd11an1n64x5 FILLER_180_200 ();
 b15zdnd11an1n64x5 FILLER_180_264 ();
 b15zdnd11an1n64x5 FILLER_180_328 ();
 b15zdnd11an1n64x5 FILLER_180_392 ();
 b15zdnd11an1n64x5 FILLER_180_456 ();
 b15zdnd11an1n32x5 FILLER_180_520 ();
 b15zdnd11an1n04x5 FILLER_180_552 ();
 b15zdnd00an1n02x5 FILLER_180_556 ();
 b15zdnd00an1n01x5 FILLER_180_558 ();
 b15zdnd11an1n64x5 FILLER_180_601 ();
 b15zdnd11an1n32x5 FILLER_180_665 ();
 b15zdnd11an1n16x5 FILLER_180_697 ();
 b15zdnd11an1n04x5 FILLER_180_713 ();
 b15zdnd00an1n01x5 FILLER_180_717 ();
 b15zdnd11an1n64x5 FILLER_180_726 ();
 b15zdnd11an1n64x5 FILLER_180_790 ();
 b15zdnd11an1n64x5 FILLER_180_854 ();
 b15zdnd11an1n64x5 FILLER_180_918 ();
 b15zdnd11an1n64x5 FILLER_180_982 ();
 b15zdnd11an1n64x5 FILLER_180_1046 ();
 b15zdnd11an1n64x5 FILLER_180_1110 ();
 b15zdnd11an1n64x5 FILLER_180_1174 ();
 b15zdnd11an1n64x5 FILLER_180_1238 ();
 b15zdnd11an1n64x5 FILLER_180_1302 ();
 b15zdnd11an1n64x5 FILLER_180_1366 ();
 b15zdnd11an1n32x5 FILLER_180_1430 ();
 b15zdnd11an1n16x5 FILLER_180_1462 ();
 b15zdnd11an1n08x5 FILLER_180_2265 ();
 b15zdnd00an1n02x5 FILLER_180_2273 ();
 b15zdnd00an1n01x5 FILLER_180_2275 ();
 b15zdnd11an1n64x5 FILLER_181_0 ();
 b15zdnd11an1n64x5 FILLER_181_64 ();
 b15zdnd11an1n64x5 FILLER_181_128 ();
 b15zdnd11an1n64x5 FILLER_181_192 ();
 b15zdnd11an1n64x5 FILLER_181_256 ();
 b15zdnd11an1n64x5 FILLER_181_320 ();
 b15zdnd11an1n32x5 FILLER_181_384 ();
 b15zdnd11an1n08x5 FILLER_181_416 ();
 b15zdnd11an1n16x5 FILLER_181_432 ();
 b15zdnd11an1n08x5 FILLER_181_448 ();
 b15zdnd11an1n64x5 FILLER_181_481 ();
 b15zdnd11an1n64x5 FILLER_181_545 ();
 b15zdnd11an1n64x5 FILLER_181_609 ();
 b15zdnd11an1n64x5 FILLER_181_673 ();
 b15zdnd11an1n64x5 FILLER_181_737 ();
 b15zdnd11an1n64x5 FILLER_181_801 ();
 b15zdnd11an1n64x5 FILLER_181_865 ();
 b15zdnd11an1n64x5 FILLER_181_929 ();
 b15zdnd11an1n64x5 FILLER_181_993 ();
 b15zdnd11an1n64x5 FILLER_181_1057 ();
 b15zdnd11an1n64x5 FILLER_181_1121 ();
 b15zdnd11an1n64x5 FILLER_181_1185 ();
 b15zdnd11an1n64x5 FILLER_181_1249 ();
 b15zdnd11an1n64x5 FILLER_181_1313 ();
 b15zdnd11an1n64x5 FILLER_181_1377 ();
 b15zdnd11an1n32x5 FILLER_181_1441 ();
 b15zdnd11an1n08x5 FILLER_181_1473 ();
 b15zdnd11an1n04x5 FILLER_181_1481 ();
 b15zdnd00an1n01x5 FILLER_181_1485 ();
 b15zdnd00an1n02x5 FILLER_181_2257 ();
 b15zdnd11an1n04x5 FILLER_181_2263 ();
 b15zdnd11an1n08x5 FILLER_181_2271 ();
 b15zdnd11an1n04x5 FILLER_181_2279 ();
 b15zdnd00an1n01x5 FILLER_181_2283 ();
 b15zdnd11an1n64x5 FILLER_182_8 ();
 b15zdnd11an1n64x5 FILLER_182_72 ();
 b15zdnd11an1n64x5 FILLER_182_136 ();
 b15zdnd11an1n64x5 FILLER_182_200 ();
 b15zdnd11an1n64x5 FILLER_182_264 ();
 b15zdnd11an1n64x5 FILLER_182_328 ();
 b15zdnd11an1n32x5 FILLER_182_392 ();
 b15zdnd11an1n16x5 FILLER_182_424 ();
 b15zdnd11an1n64x5 FILLER_182_482 ();
 b15zdnd11an1n64x5 FILLER_182_546 ();
 b15zdnd11an1n64x5 FILLER_182_610 ();
 b15zdnd11an1n32x5 FILLER_182_674 ();
 b15zdnd11an1n08x5 FILLER_182_706 ();
 b15zdnd11an1n04x5 FILLER_182_714 ();
 b15zdnd11an1n64x5 FILLER_182_726 ();
 b15zdnd11an1n64x5 FILLER_182_790 ();
 b15zdnd11an1n64x5 FILLER_182_854 ();
 b15zdnd11an1n64x5 FILLER_182_918 ();
 b15zdnd11an1n64x5 FILLER_182_982 ();
 b15zdnd11an1n64x5 FILLER_182_1046 ();
 b15zdnd11an1n64x5 FILLER_182_1110 ();
 b15zdnd11an1n64x5 FILLER_182_1174 ();
 b15zdnd11an1n64x5 FILLER_182_1238 ();
 b15zdnd11an1n64x5 FILLER_182_1302 ();
 b15zdnd11an1n64x5 FILLER_182_1366 ();
 b15zdnd11an1n32x5 FILLER_182_1430 ();
 b15zdnd11an1n16x5 FILLER_182_1462 ();
 b15zdnd11an1n08x5 FILLER_182_2265 ();
 b15zdnd00an1n02x5 FILLER_182_2273 ();
 b15zdnd00an1n01x5 FILLER_182_2275 ();
 b15zdnd11an1n64x5 FILLER_183_0 ();
 b15zdnd11an1n64x5 FILLER_183_64 ();
 b15zdnd11an1n64x5 FILLER_183_128 ();
 b15zdnd11an1n64x5 FILLER_183_192 ();
 b15zdnd11an1n64x5 FILLER_183_256 ();
 b15zdnd11an1n64x5 FILLER_183_320 ();
 b15zdnd11an1n64x5 FILLER_183_384 ();
 b15zdnd11an1n64x5 FILLER_183_448 ();
 b15zdnd11an1n64x5 FILLER_183_512 ();
 b15zdnd11an1n64x5 FILLER_183_576 ();
 b15zdnd11an1n64x5 FILLER_183_640 ();
 b15zdnd11an1n64x5 FILLER_183_704 ();
 b15zdnd11an1n64x5 FILLER_183_768 ();
 b15zdnd11an1n64x5 FILLER_183_832 ();
 b15zdnd11an1n64x5 FILLER_183_896 ();
 b15zdnd11an1n64x5 FILLER_183_960 ();
 b15zdnd11an1n64x5 FILLER_183_1024 ();
 b15zdnd11an1n64x5 FILLER_183_1088 ();
 b15zdnd11an1n64x5 FILLER_183_1152 ();
 b15zdnd11an1n64x5 FILLER_183_1216 ();
 b15zdnd11an1n64x5 FILLER_183_1280 ();
 b15zdnd11an1n64x5 FILLER_183_1344 ();
 b15zdnd11an1n64x5 FILLER_183_1408 ();
 b15zdnd11an1n08x5 FILLER_183_1472 ();
 b15zdnd11an1n04x5 FILLER_183_1480 ();
 b15zdnd00an1n02x5 FILLER_183_1484 ();
 b15zdnd11an1n16x5 FILLER_183_2257 ();
 b15zdnd11an1n08x5 FILLER_183_2273 ();
 b15zdnd00an1n02x5 FILLER_183_2281 ();
 b15zdnd00an1n01x5 FILLER_183_2283 ();
 b15zdnd11an1n64x5 FILLER_184_8 ();
 b15zdnd11an1n64x5 FILLER_184_72 ();
 b15zdnd11an1n64x5 FILLER_184_136 ();
 b15zdnd11an1n64x5 FILLER_184_200 ();
 b15zdnd11an1n64x5 FILLER_184_264 ();
 b15zdnd11an1n64x5 FILLER_184_328 ();
 b15zdnd11an1n16x5 FILLER_184_392 ();
 b15zdnd11an1n08x5 FILLER_184_408 ();
 b15zdnd11an1n64x5 FILLER_184_420 ();
 b15zdnd11an1n64x5 FILLER_184_484 ();
 b15zdnd11an1n64x5 FILLER_184_548 ();
 b15zdnd11an1n64x5 FILLER_184_612 ();
 b15zdnd11an1n32x5 FILLER_184_676 ();
 b15zdnd11an1n08x5 FILLER_184_708 ();
 b15zdnd00an1n02x5 FILLER_184_716 ();
 b15zdnd11an1n64x5 FILLER_184_726 ();
 b15zdnd11an1n64x5 FILLER_184_790 ();
 b15zdnd11an1n64x5 FILLER_184_854 ();
 b15zdnd11an1n64x5 FILLER_184_918 ();
 b15zdnd11an1n64x5 FILLER_184_982 ();
 b15zdnd11an1n64x5 FILLER_184_1046 ();
 b15zdnd11an1n64x5 FILLER_184_1110 ();
 b15zdnd11an1n64x5 FILLER_184_1174 ();
 b15zdnd11an1n16x5 FILLER_184_1238 ();
 b15zdnd11an1n08x5 FILLER_184_1254 ();
 b15zdnd11an1n04x5 FILLER_184_1262 ();
 b15zdnd00an1n01x5 FILLER_184_1266 ();
 b15zdnd11an1n64x5 FILLER_184_1309 ();
 b15zdnd11an1n64x5 FILLER_184_1373 ();
 b15zdnd11an1n32x5 FILLER_184_1437 ();
 b15zdnd11an1n08x5 FILLER_184_1469 ();
 b15zdnd00an1n01x5 FILLER_184_1477 ();
 b15zdnd11an1n08x5 FILLER_184_2265 ();
 b15zdnd00an1n02x5 FILLER_184_2273 ();
 b15zdnd00an1n01x5 FILLER_184_2275 ();
 b15zdnd11an1n64x5 FILLER_185_0 ();
 b15zdnd11an1n64x5 FILLER_185_64 ();
 b15zdnd11an1n64x5 FILLER_185_128 ();
 b15zdnd11an1n64x5 FILLER_185_192 ();
 b15zdnd11an1n64x5 FILLER_185_256 ();
 b15zdnd11an1n64x5 FILLER_185_320 ();
 b15zdnd11an1n32x5 FILLER_185_384 ();
 b15zdnd11an1n04x5 FILLER_185_416 ();
 b15zdnd00an1n01x5 FILLER_185_420 ();
 b15zdnd11an1n64x5 FILLER_185_454 ();
 b15zdnd11an1n64x5 FILLER_185_518 ();
 b15zdnd11an1n64x5 FILLER_185_582 ();
 b15zdnd11an1n64x5 FILLER_185_646 ();
 b15zdnd11an1n64x5 FILLER_185_710 ();
 b15zdnd11an1n64x5 FILLER_185_774 ();
 b15zdnd11an1n64x5 FILLER_185_838 ();
 b15zdnd11an1n64x5 FILLER_185_902 ();
 b15zdnd11an1n64x5 FILLER_185_966 ();
 b15zdnd11an1n64x5 FILLER_185_1030 ();
 b15zdnd11an1n64x5 FILLER_185_1094 ();
 b15zdnd11an1n64x5 FILLER_185_1158 ();
 b15zdnd11an1n64x5 FILLER_185_1222 ();
 b15zdnd11an1n64x5 FILLER_185_1286 ();
 b15zdnd11an1n64x5 FILLER_185_1350 ();
 b15zdnd11an1n64x5 FILLER_185_1414 ();
 b15zdnd11an1n08x5 FILLER_185_1478 ();
 b15zdnd11an1n16x5 FILLER_185_2257 ();
 b15zdnd11an1n08x5 FILLER_185_2273 ();
 b15zdnd00an1n02x5 FILLER_185_2281 ();
 b15zdnd00an1n01x5 FILLER_185_2283 ();
 b15zdnd11an1n64x5 FILLER_186_8 ();
 b15zdnd11an1n64x5 FILLER_186_72 ();
 b15zdnd11an1n64x5 FILLER_186_136 ();
 b15zdnd11an1n64x5 FILLER_186_200 ();
 b15zdnd11an1n64x5 FILLER_186_264 ();
 b15zdnd11an1n64x5 FILLER_186_328 ();
 b15zdnd11an1n64x5 FILLER_186_392 ();
 b15zdnd11an1n08x5 FILLER_186_456 ();
 b15zdnd11an1n04x5 FILLER_186_464 ();
 b15zdnd11an1n04x5 FILLER_186_510 ();
 b15zdnd11an1n64x5 FILLER_186_534 ();
 b15zdnd11an1n64x5 FILLER_186_598 ();
 b15zdnd11an1n32x5 FILLER_186_662 ();
 b15zdnd11an1n16x5 FILLER_186_694 ();
 b15zdnd11an1n08x5 FILLER_186_710 ();
 b15zdnd11an1n64x5 FILLER_186_726 ();
 b15zdnd11an1n64x5 FILLER_186_790 ();
 b15zdnd11an1n64x5 FILLER_186_854 ();
 b15zdnd11an1n08x5 FILLER_186_918 ();
 b15zdnd11an1n04x5 FILLER_186_926 ();
 b15zdnd00an1n02x5 FILLER_186_930 ();
 b15zdnd11an1n64x5 FILLER_186_974 ();
 b15zdnd11an1n64x5 FILLER_186_1038 ();
 b15zdnd11an1n64x5 FILLER_186_1102 ();
 b15zdnd11an1n64x5 FILLER_186_1166 ();
 b15zdnd11an1n64x5 FILLER_186_1230 ();
 b15zdnd11an1n64x5 FILLER_186_1294 ();
 b15zdnd11an1n64x5 FILLER_186_1358 ();
 b15zdnd11an1n32x5 FILLER_186_1422 ();
 b15zdnd11an1n16x5 FILLER_186_1454 ();
 b15zdnd11an1n08x5 FILLER_186_1470 ();
 b15zdnd11an1n08x5 FILLER_186_2265 ();
 b15zdnd00an1n02x5 FILLER_186_2273 ();
 b15zdnd00an1n01x5 FILLER_186_2275 ();
 b15zdnd11an1n64x5 FILLER_187_0 ();
 b15zdnd11an1n64x5 FILLER_187_64 ();
 b15zdnd11an1n64x5 FILLER_187_128 ();
 b15zdnd11an1n64x5 FILLER_187_192 ();
 b15zdnd11an1n64x5 FILLER_187_256 ();
 b15zdnd11an1n64x5 FILLER_187_320 ();
 b15zdnd11an1n64x5 FILLER_187_384 ();
 b15zdnd11an1n32x5 FILLER_187_448 ();
 b15zdnd11an1n16x5 FILLER_187_480 ();
 b15zdnd11an1n08x5 FILLER_187_496 ();
 b15zdnd11an1n04x5 FILLER_187_504 ();
 b15zdnd00an1n02x5 FILLER_187_508 ();
 b15zdnd11an1n64x5 FILLER_187_530 ();
 b15zdnd11an1n64x5 FILLER_187_594 ();
 b15zdnd11an1n64x5 FILLER_187_658 ();
 b15zdnd11an1n64x5 FILLER_187_722 ();
 b15zdnd11an1n64x5 FILLER_187_786 ();
 b15zdnd11an1n64x5 FILLER_187_850 ();
 b15zdnd11an1n08x5 FILLER_187_914 ();
 b15zdnd11an1n64x5 FILLER_187_964 ();
 b15zdnd11an1n64x5 FILLER_187_1028 ();
 b15zdnd11an1n64x5 FILLER_187_1092 ();
 b15zdnd11an1n64x5 FILLER_187_1156 ();
 b15zdnd11an1n16x5 FILLER_187_1220 ();
 b15zdnd00an1n02x5 FILLER_187_1236 ();
 b15zdnd11an1n64x5 FILLER_187_1258 ();
 b15zdnd11an1n64x5 FILLER_187_1322 ();
 b15zdnd11an1n64x5 FILLER_187_1386 ();
 b15zdnd11an1n32x5 FILLER_187_1450 ();
 b15zdnd11an1n04x5 FILLER_187_1482 ();
 b15zdnd11an1n16x5 FILLER_187_2257 ();
 b15zdnd11an1n08x5 FILLER_187_2273 ();
 b15zdnd00an1n02x5 FILLER_187_2281 ();
 b15zdnd00an1n01x5 FILLER_187_2283 ();
 b15zdnd11an1n64x5 FILLER_188_8 ();
 b15zdnd11an1n64x5 FILLER_188_72 ();
 b15zdnd11an1n64x5 FILLER_188_136 ();
 b15zdnd11an1n64x5 FILLER_188_200 ();
 b15zdnd11an1n64x5 FILLER_188_264 ();
 b15zdnd11an1n64x5 FILLER_188_328 ();
 b15zdnd11an1n64x5 FILLER_188_392 ();
 b15zdnd11an1n64x5 FILLER_188_456 ();
 b15zdnd11an1n64x5 FILLER_188_520 ();
 b15zdnd11an1n64x5 FILLER_188_584 ();
 b15zdnd11an1n64x5 FILLER_188_648 ();
 b15zdnd11an1n04x5 FILLER_188_712 ();
 b15zdnd00an1n02x5 FILLER_188_716 ();
 b15zdnd11an1n64x5 FILLER_188_726 ();
 b15zdnd11an1n64x5 FILLER_188_790 ();
 b15zdnd11an1n64x5 FILLER_188_854 ();
 b15zdnd11an1n64x5 FILLER_188_918 ();
 b15zdnd11an1n64x5 FILLER_188_982 ();
 b15zdnd11an1n64x5 FILLER_188_1046 ();
 b15zdnd11an1n64x5 FILLER_188_1110 ();
 b15zdnd11an1n64x5 FILLER_188_1174 ();
 b15zdnd11an1n32x5 FILLER_188_1238 ();
 b15zdnd11an1n04x5 FILLER_188_1270 ();
 b15zdnd00an1n01x5 FILLER_188_1274 ();
 b15zdnd11an1n04x5 FILLER_188_1301 ();
 b15zdnd11an1n64x5 FILLER_188_1319 ();
 b15zdnd11an1n64x5 FILLER_188_1383 ();
 b15zdnd11an1n16x5 FILLER_188_1447 ();
 b15zdnd11an1n08x5 FILLER_188_1463 ();
 b15zdnd11an1n04x5 FILLER_188_1471 ();
 b15zdnd00an1n02x5 FILLER_188_1475 ();
 b15zdnd00an1n01x5 FILLER_188_1477 ();
 b15zdnd11an1n08x5 FILLER_188_2265 ();
 b15zdnd00an1n02x5 FILLER_188_2273 ();
 b15zdnd00an1n01x5 FILLER_188_2275 ();
 b15zdnd11an1n64x5 FILLER_189_0 ();
 b15zdnd11an1n64x5 FILLER_189_64 ();
 b15zdnd11an1n64x5 FILLER_189_128 ();
 b15zdnd11an1n64x5 FILLER_189_192 ();
 b15zdnd11an1n64x5 FILLER_189_256 ();
 b15zdnd11an1n64x5 FILLER_189_320 ();
 b15zdnd11an1n64x5 FILLER_189_384 ();
 b15zdnd11an1n64x5 FILLER_189_448 ();
 b15zdnd11an1n64x5 FILLER_189_512 ();
 b15zdnd11an1n64x5 FILLER_189_576 ();
 b15zdnd11an1n64x5 FILLER_189_640 ();
 b15zdnd11an1n64x5 FILLER_189_704 ();
 b15zdnd11an1n64x5 FILLER_189_768 ();
 b15zdnd11an1n64x5 FILLER_189_832 ();
 b15zdnd11an1n64x5 FILLER_189_896 ();
 b15zdnd11an1n64x5 FILLER_189_960 ();
 b15zdnd11an1n64x5 FILLER_189_1024 ();
 b15zdnd11an1n64x5 FILLER_189_1088 ();
 b15zdnd11an1n64x5 FILLER_189_1152 ();
 b15zdnd11an1n64x5 FILLER_189_1216 ();
 b15zdnd11an1n32x5 FILLER_189_1280 ();
 b15zdnd00an1n01x5 FILLER_189_1312 ();
 b15zdnd11an1n04x5 FILLER_189_1327 ();
 b15zdnd00an1n02x5 FILLER_189_1331 ();
 b15zdnd00an1n01x5 FILLER_189_1333 ();
 b15zdnd11an1n64x5 FILLER_189_1358 ();
 b15zdnd11an1n64x5 FILLER_189_1422 ();
 b15zdnd11an1n16x5 FILLER_189_2257 ();
 b15zdnd11an1n08x5 FILLER_189_2273 ();
 b15zdnd00an1n02x5 FILLER_189_2281 ();
 b15zdnd00an1n01x5 FILLER_189_2283 ();
 b15zdnd11an1n64x5 FILLER_190_8 ();
 b15zdnd11an1n64x5 FILLER_190_72 ();
 b15zdnd11an1n64x5 FILLER_190_136 ();
 b15zdnd11an1n64x5 FILLER_190_200 ();
 b15zdnd11an1n64x5 FILLER_190_264 ();
 b15zdnd11an1n64x5 FILLER_190_328 ();
 b15zdnd11an1n16x5 FILLER_190_392 ();
 b15zdnd11an1n08x5 FILLER_190_408 ();
 b15zdnd00an1n02x5 FILLER_190_416 ();
 b15zdnd11an1n32x5 FILLER_190_425 ();
 b15zdnd11an1n04x5 FILLER_190_457 ();
 b15zdnd11an1n64x5 FILLER_190_479 ();
 b15zdnd11an1n64x5 FILLER_190_543 ();
 b15zdnd11an1n64x5 FILLER_190_607 ();
 b15zdnd11an1n32x5 FILLER_190_671 ();
 b15zdnd11an1n08x5 FILLER_190_703 ();
 b15zdnd11an1n04x5 FILLER_190_711 ();
 b15zdnd00an1n02x5 FILLER_190_715 ();
 b15zdnd00an1n01x5 FILLER_190_717 ();
 b15zdnd11an1n64x5 FILLER_190_726 ();
 b15zdnd11an1n64x5 FILLER_190_790 ();
 b15zdnd11an1n64x5 FILLER_190_854 ();
 b15zdnd11an1n64x5 FILLER_190_918 ();
 b15zdnd11an1n64x5 FILLER_190_982 ();
 b15zdnd11an1n64x5 FILLER_190_1046 ();
 b15zdnd11an1n64x5 FILLER_190_1110 ();
 b15zdnd11an1n64x5 FILLER_190_1174 ();
 b15zdnd11an1n32x5 FILLER_190_1238 ();
 b15zdnd11an1n16x5 FILLER_190_1270 ();
 b15zdnd11an1n08x5 FILLER_190_1286 ();
 b15zdnd11an1n04x5 FILLER_190_1294 ();
 b15zdnd00an1n01x5 FILLER_190_1298 ();
 b15zdnd11an1n64x5 FILLER_190_1315 ();
 b15zdnd11an1n64x5 FILLER_190_1379 ();
 b15zdnd11an1n32x5 FILLER_190_1443 ();
 b15zdnd00an1n02x5 FILLER_190_1475 ();
 b15zdnd00an1n01x5 FILLER_190_1477 ();
 b15zdnd11an1n08x5 FILLER_190_2265 ();
 b15zdnd00an1n02x5 FILLER_190_2273 ();
 b15zdnd00an1n01x5 FILLER_190_2275 ();
 b15zdnd11an1n64x5 FILLER_191_0 ();
 b15zdnd11an1n64x5 FILLER_191_64 ();
 b15zdnd11an1n64x5 FILLER_191_128 ();
 b15zdnd11an1n64x5 FILLER_191_192 ();
 b15zdnd11an1n64x5 FILLER_191_256 ();
 b15zdnd11an1n64x5 FILLER_191_320 ();
 b15zdnd11an1n64x5 FILLER_191_384 ();
 b15zdnd11an1n64x5 FILLER_191_448 ();
 b15zdnd11an1n64x5 FILLER_191_512 ();
 b15zdnd11an1n64x5 FILLER_191_576 ();
 b15zdnd11an1n64x5 FILLER_191_640 ();
 b15zdnd11an1n64x5 FILLER_191_704 ();
 b15zdnd11an1n64x5 FILLER_191_768 ();
 b15zdnd11an1n64x5 FILLER_191_832 ();
 b15zdnd11an1n64x5 FILLER_191_896 ();
 b15zdnd11an1n64x5 FILLER_191_960 ();
 b15zdnd11an1n64x5 FILLER_191_1024 ();
 b15zdnd11an1n64x5 FILLER_191_1088 ();
 b15zdnd11an1n64x5 FILLER_191_1152 ();
 b15zdnd11an1n64x5 FILLER_191_1216 ();
 b15zdnd11an1n32x5 FILLER_191_1280 ();
 b15zdnd11an1n04x5 FILLER_191_1312 ();
 b15zdnd11an1n64x5 FILLER_191_1347 ();
 b15zdnd11an1n64x5 FILLER_191_1411 ();
 b15zdnd11an1n08x5 FILLER_191_1475 ();
 b15zdnd00an1n02x5 FILLER_191_1483 ();
 b15zdnd00an1n01x5 FILLER_191_1485 ();
 b15zdnd11an1n16x5 FILLER_191_2257 ();
 b15zdnd11an1n08x5 FILLER_191_2273 ();
 b15zdnd00an1n02x5 FILLER_191_2281 ();
 b15zdnd00an1n01x5 FILLER_191_2283 ();
 b15zdnd11an1n64x5 FILLER_192_8 ();
 b15zdnd11an1n64x5 FILLER_192_72 ();
 b15zdnd11an1n64x5 FILLER_192_136 ();
 b15zdnd11an1n64x5 FILLER_192_200 ();
 b15zdnd11an1n64x5 FILLER_192_264 ();
 b15zdnd11an1n64x5 FILLER_192_328 ();
 b15zdnd11an1n64x5 FILLER_192_392 ();
 b15zdnd11an1n16x5 FILLER_192_456 ();
 b15zdnd11an1n08x5 FILLER_192_472 ();
 b15zdnd11an1n04x5 FILLER_192_480 ();
 b15zdnd00an1n01x5 FILLER_192_484 ();
 b15zdnd11an1n64x5 FILLER_192_499 ();
 b15zdnd11an1n64x5 FILLER_192_563 ();
 b15zdnd11an1n64x5 FILLER_192_627 ();
 b15zdnd11an1n16x5 FILLER_192_691 ();
 b15zdnd11an1n08x5 FILLER_192_707 ();
 b15zdnd00an1n02x5 FILLER_192_715 ();
 b15zdnd00an1n01x5 FILLER_192_717 ();
 b15zdnd11an1n64x5 FILLER_192_726 ();
 b15zdnd11an1n64x5 FILLER_192_790 ();
 b15zdnd11an1n64x5 FILLER_192_854 ();
 b15zdnd11an1n64x5 FILLER_192_918 ();
 b15zdnd11an1n64x5 FILLER_192_982 ();
 b15zdnd11an1n64x5 FILLER_192_1046 ();
 b15zdnd11an1n64x5 FILLER_192_1110 ();
 b15zdnd11an1n64x5 FILLER_192_1174 ();
 b15zdnd11an1n64x5 FILLER_192_1238 ();
 b15zdnd11an1n64x5 FILLER_192_1302 ();
 b15zdnd11an1n64x5 FILLER_192_1366 ();
 b15zdnd11an1n32x5 FILLER_192_1430 ();
 b15zdnd11an1n16x5 FILLER_192_1462 ();
 b15zdnd11an1n08x5 FILLER_192_2265 ();
 b15zdnd00an1n02x5 FILLER_192_2273 ();
 b15zdnd00an1n01x5 FILLER_192_2275 ();
 b15zdnd11an1n64x5 FILLER_193_0 ();
 b15zdnd11an1n64x5 FILLER_193_64 ();
 b15zdnd11an1n64x5 FILLER_193_128 ();
 b15zdnd11an1n64x5 FILLER_193_192 ();
 b15zdnd11an1n64x5 FILLER_193_256 ();
 b15zdnd11an1n64x5 FILLER_193_320 ();
 b15zdnd11an1n64x5 FILLER_193_384 ();
 b15zdnd11an1n64x5 FILLER_193_448 ();
 b15zdnd11an1n64x5 FILLER_193_512 ();
 b15zdnd11an1n64x5 FILLER_193_576 ();
 b15zdnd11an1n64x5 FILLER_193_640 ();
 b15zdnd11an1n64x5 FILLER_193_704 ();
 b15zdnd11an1n64x5 FILLER_193_768 ();
 b15zdnd11an1n64x5 FILLER_193_832 ();
 b15zdnd11an1n64x5 FILLER_193_896 ();
 b15zdnd11an1n64x5 FILLER_193_960 ();
 b15zdnd11an1n64x5 FILLER_193_1024 ();
 b15zdnd11an1n64x5 FILLER_193_1088 ();
 b15zdnd11an1n64x5 FILLER_193_1152 ();
 b15zdnd11an1n64x5 FILLER_193_1216 ();
 b15zdnd11an1n64x5 FILLER_193_1280 ();
 b15zdnd11an1n64x5 FILLER_193_1344 ();
 b15zdnd11an1n64x5 FILLER_193_1408 ();
 b15zdnd11an1n08x5 FILLER_193_1472 ();
 b15zdnd11an1n04x5 FILLER_193_1480 ();
 b15zdnd00an1n02x5 FILLER_193_1484 ();
 b15zdnd11an1n16x5 FILLER_193_2257 ();
 b15zdnd11an1n08x5 FILLER_193_2273 ();
 b15zdnd00an1n02x5 FILLER_193_2281 ();
 b15zdnd00an1n01x5 FILLER_193_2283 ();
 b15zdnd11an1n64x5 FILLER_194_8 ();
 b15zdnd11an1n64x5 FILLER_194_72 ();
 b15zdnd11an1n64x5 FILLER_194_136 ();
 b15zdnd11an1n64x5 FILLER_194_200 ();
 b15zdnd11an1n64x5 FILLER_194_264 ();
 b15zdnd11an1n64x5 FILLER_194_328 ();
 b15zdnd11an1n64x5 FILLER_194_392 ();
 b15zdnd11an1n64x5 FILLER_194_456 ();
 b15zdnd11an1n64x5 FILLER_194_520 ();
 b15zdnd11an1n64x5 FILLER_194_584 ();
 b15zdnd11an1n64x5 FILLER_194_648 ();
 b15zdnd11an1n04x5 FILLER_194_712 ();
 b15zdnd00an1n02x5 FILLER_194_716 ();
 b15zdnd11an1n64x5 FILLER_194_726 ();
 b15zdnd11an1n64x5 FILLER_194_790 ();
 b15zdnd11an1n64x5 FILLER_194_854 ();
 b15zdnd11an1n64x5 FILLER_194_918 ();
 b15zdnd11an1n64x5 FILLER_194_982 ();
 b15zdnd11an1n64x5 FILLER_194_1046 ();
 b15zdnd11an1n64x5 FILLER_194_1110 ();
 b15zdnd11an1n64x5 FILLER_194_1174 ();
 b15zdnd11an1n64x5 FILLER_194_1238 ();
 b15zdnd11an1n64x5 FILLER_194_1302 ();
 b15zdnd11an1n64x5 FILLER_194_1366 ();
 b15zdnd11an1n16x5 FILLER_194_1430 ();
 b15zdnd11an1n08x5 FILLER_194_1446 ();
 b15zdnd00an1n02x5 FILLER_194_1454 ();
 b15zdnd00an1n02x5 FILLER_194_1476 ();
 b15zdnd11an1n08x5 FILLER_194_2265 ();
 b15zdnd00an1n02x5 FILLER_194_2273 ();
 b15zdnd00an1n01x5 FILLER_194_2275 ();
 b15zdnd11an1n64x5 FILLER_195_0 ();
 b15zdnd11an1n64x5 FILLER_195_64 ();
 b15zdnd11an1n64x5 FILLER_195_128 ();
 b15zdnd11an1n64x5 FILLER_195_192 ();
 b15zdnd11an1n64x5 FILLER_195_256 ();
 b15zdnd11an1n64x5 FILLER_195_320 ();
 b15zdnd11an1n64x5 FILLER_195_384 ();
 b15zdnd11an1n64x5 FILLER_195_448 ();
 b15zdnd11an1n64x5 FILLER_195_512 ();
 b15zdnd11an1n64x5 FILLER_195_576 ();
 b15zdnd11an1n64x5 FILLER_195_640 ();
 b15zdnd11an1n64x5 FILLER_195_704 ();
 b15zdnd11an1n64x5 FILLER_195_768 ();
 b15zdnd11an1n64x5 FILLER_195_832 ();
 b15zdnd11an1n64x5 FILLER_195_896 ();
 b15zdnd11an1n64x5 FILLER_195_960 ();
 b15zdnd11an1n64x5 FILLER_195_1024 ();
 b15zdnd11an1n64x5 FILLER_195_1088 ();
 b15zdnd11an1n64x5 FILLER_195_1152 ();
 b15zdnd11an1n64x5 FILLER_195_1216 ();
 b15zdnd11an1n64x5 FILLER_195_1280 ();
 b15zdnd11an1n64x5 FILLER_195_1344 ();
 b15zdnd11an1n64x5 FILLER_195_1408 ();
 b15zdnd11an1n08x5 FILLER_195_1472 ();
 b15zdnd11an1n04x5 FILLER_195_1480 ();
 b15zdnd00an1n02x5 FILLER_195_1484 ();
 b15zdnd11an1n16x5 FILLER_195_2257 ();
 b15zdnd11an1n08x5 FILLER_195_2273 ();
 b15zdnd00an1n02x5 FILLER_195_2281 ();
 b15zdnd00an1n01x5 FILLER_195_2283 ();
 b15zdnd11an1n64x5 FILLER_196_8 ();
 b15zdnd11an1n64x5 FILLER_196_72 ();
 b15zdnd11an1n64x5 FILLER_196_136 ();
 b15zdnd11an1n64x5 FILLER_196_200 ();
 b15zdnd11an1n64x5 FILLER_196_264 ();
 b15zdnd11an1n64x5 FILLER_196_328 ();
 b15zdnd11an1n64x5 FILLER_196_392 ();
 b15zdnd11an1n32x5 FILLER_196_456 ();
 b15zdnd11an1n08x5 FILLER_196_488 ();
 b15zdnd11an1n04x5 FILLER_196_496 ();
 b15zdnd00an1n02x5 FILLER_196_500 ();
 b15zdnd00an1n01x5 FILLER_196_502 ();
 b15zdnd11an1n64x5 FILLER_196_545 ();
 b15zdnd11an1n64x5 FILLER_196_609 ();
 b15zdnd11an1n32x5 FILLER_196_673 ();
 b15zdnd11an1n08x5 FILLER_196_705 ();
 b15zdnd11an1n04x5 FILLER_196_713 ();
 b15zdnd00an1n01x5 FILLER_196_717 ();
 b15zdnd11an1n64x5 FILLER_196_726 ();
 b15zdnd11an1n08x5 FILLER_196_790 ();
 b15zdnd11an1n64x5 FILLER_196_807 ();
 b15zdnd11an1n64x5 FILLER_196_871 ();
 b15zdnd11an1n64x5 FILLER_196_935 ();
 b15zdnd11an1n32x5 FILLER_196_999 ();
 b15zdnd11an1n16x5 FILLER_196_1031 ();
 b15zdnd00an1n02x5 FILLER_196_1047 ();
 b15zdnd11an1n64x5 FILLER_196_1056 ();
 b15zdnd11an1n64x5 FILLER_196_1120 ();
 b15zdnd11an1n08x5 FILLER_196_1184 ();
 b15zdnd11an1n04x5 FILLER_196_1192 ();
 b15zdnd00an1n02x5 FILLER_196_1196 ();
 b15zdnd00an1n01x5 FILLER_196_1198 ();
 b15zdnd11an1n64x5 FILLER_196_1210 ();
 b15zdnd11an1n64x5 FILLER_196_1274 ();
 b15zdnd11an1n16x5 FILLER_196_1338 ();
 b15zdnd00an1n02x5 FILLER_196_1354 ();
 b15zdnd00an1n01x5 FILLER_196_1356 ();
 b15zdnd11an1n08x5 FILLER_196_1399 ();
 b15zdnd11an1n04x5 FILLER_196_1407 ();
 b15zdnd11an1n32x5 FILLER_196_1431 ();
 b15zdnd11an1n08x5 FILLER_196_1463 ();
 b15zdnd11an1n04x5 FILLER_196_1471 ();
 b15zdnd00an1n02x5 FILLER_196_1475 ();
 b15zdnd00an1n01x5 FILLER_196_1477 ();
 b15zdnd11an1n08x5 FILLER_196_2265 ();
 b15zdnd00an1n02x5 FILLER_196_2273 ();
 b15zdnd00an1n01x5 FILLER_196_2275 ();
 b15zdnd11an1n16x5 FILLER_197_0 ();
 b15zdnd00an1n01x5 FILLER_197_16 ();
 b15zdnd11an1n04x5 FILLER_197_21 ();
 b15zdnd00an1n02x5 FILLER_197_25 ();
 b15zdnd11an1n64x5 FILLER_197_31 ();
 b15zdnd11an1n64x5 FILLER_197_95 ();
 b15zdnd11an1n64x5 FILLER_197_159 ();
 b15zdnd11an1n64x5 FILLER_197_223 ();
 b15zdnd11an1n64x5 FILLER_197_287 ();
 b15zdnd11an1n64x5 FILLER_197_351 ();
 b15zdnd11an1n64x5 FILLER_197_415 ();
 b15zdnd11an1n64x5 FILLER_197_479 ();
 b15zdnd11an1n64x5 FILLER_197_543 ();
 b15zdnd11an1n64x5 FILLER_197_607 ();
 b15zdnd11an1n64x5 FILLER_197_671 ();
 b15zdnd11an1n64x5 FILLER_197_735 ();
 b15zdnd11an1n64x5 FILLER_197_799 ();
 b15zdnd11an1n64x5 FILLER_197_863 ();
 b15zdnd11an1n64x5 FILLER_197_927 ();
 b15zdnd11an1n64x5 FILLER_197_991 ();
 b15zdnd11an1n64x5 FILLER_197_1055 ();
 b15zdnd11an1n32x5 FILLER_197_1119 ();
 b15zdnd11an1n16x5 FILLER_197_1151 ();
 b15zdnd11an1n08x5 FILLER_197_1167 ();
 b15zdnd00an1n01x5 FILLER_197_1175 ();
 b15zdnd11an1n08x5 FILLER_197_1192 ();
 b15zdnd00an1n01x5 FILLER_197_1200 ();
 b15zdnd11an1n64x5 FILLER_197_1210 ();
 b15zdnd11an1n64x5 FILLER_197_1274 ();
 b15zdnd11an1n64x5 FILLER_197_1338 ();
 b15zdnd11an1n64x5 FILLER_197_1402 ();
 b15zdnd11an1n16x5 FILLER_197_1466 ();
 b15zdnd11an1n04x5 FILLER_197_1482 ();
 b15zdnd11an1n16x5 FILLER_197_2257 ();
 b15zdnd11an1n08x5 FILLER_197_2273 ();
 b15zdnd00an1n02x5 FILLER_197_2281 ();
 b15zdnd00an1n01x5 FILLER_197_2283 ();
 b15zdnd00an1n02x5 FILLER_198_8 ();
 b15zdnd11an1n64x5 FILLER_198_52 ();
 b15zdnd11an1n64x5 FILLER_198_116 ();
 b15zdnd11an1n64x5 FILLER_198_180 ();
 b15zdnd11an1n64x5 FILLER_198_244 ();
 b15zdnd11an1n64x5 FILLER_198_308 ();
 b15zdnd11an1n64x5 FILLER_198_372 ();
 b15zdnd11an1n64x5 FILLER_198_436 ();
 b15zdnd11an1n64x5 FILLER_198_500 ();
 b15zdnd11an1n64x5 FILLER_198_564 ();
 b15zdnd11an1n64x5 FILLER_198_628 ();
 b15zdnd11an1n16x5 FILLER_198_692 ();
 b15zdnd11an1n08x5 FILLER_198_708 ();
 b15zdnd00an1n02x5 FILLER_198_716 ();
 b15zdnd11an1n64x5 FILLER_198_726 ();
 b15zdnd11an1n64x5 FILLER_198_790 ();
 b15zdnd11an1n64x5 FILLER_198_854 ();
 b15zdnd11an1n64x5 FILLER_198_918 ();
 b15zdnd11an1n64x5 FILLER_198_982 ();
 b15zdnd11an1n64x5 FILLER_198_1046 ();
 b15zdnd11an1n64x5 FILLER_198_1110 ();
 b15zdnd11an1n64x5 FILLER_198_1174 ();
 b15zdnd11an1n64x5 FILLER_198_1238 ();
 b15zdnd11an1n64x5 FILLER_198_1302 ();
 b15zdnd11an1n64x5 FILLER_198_1366 ();
 b15zdnd11an1n04x5 FILLER_198_1430 ();
 b15zdnd00an1n02x5 FILLER_198_1434 ();
 b15zdnd11an1n64x5 FILLER_198_1444 ();
 b15zdnd11an1n64x5 FILLER_198_1508 ();
 b15zdnd11an1n64x5 FILLER_198_1572 ();
 b15zdnd11an1n32x5 FILLER_198_1636 ();
 b15zdnd00an1n02x5 FILLER_198_1668 ();
 b15zdnd11an1n04x5 FILLER_198_1673 ();
 b15zdnd11an1n64x5 FILLER_198_1712 ();
 b15zdnd11an1n64x5 FILLER_198_1776 ();
 b15zdnd11an1n64x5 FILLER_198_1840 ();
 b15zdnd11an1n64x5 FILLER_198_1904 ();
 b15zdnd11an1n64x5 FILLER_198_1968 ();
 b15zdnd11an1n64x5 FILLER_198_2032 ();
 b15zdnd11an1n32x5 FILLER_198_2096 ();
 b15zdnd11an1n16x5 FILLER_198_2128 ();
 b15zdnd11an1n08x5 FILLER_198_2144 ();
 b15zdnd00an1n02x5 FILLER_198_2152 ();
 b15zdnd11an1n64x5 FILLER_198_2162 ();
 b15zdnd11an1n04x5 FILLER_198_2226 ();
 b15zdnd00an1n02x5 FILLER_198_2230 ();
 b15zdnd00an1n02x5 FILLER_198_2274 ();
 b15zdnd11an1n64x5 FILLER_199_0 ();
 b15zdnd11an1n64x5 FILLER_199_64 ();
 b15zdnd11an1n64x5 FILLER_199_128 ();
 b15zdnd11an1n64x5 FILLER_199_192 ();
 b15zdnd11an1n64x5 FILLER_199_256 ();
 b15zdnd11an1n64x5 FILLER_199_320 ();
 b15zdnd11an1n64x5 FILLER_199_384 ();
 b15zdnd11an1n64x5 FILLER_199_448 ();
 b15zdnd11an1n64x5 FILLER_199_512 ();
 b15zdnd11an1n64x5 FILLER_199_576 ();
 b15zdnd11an1n64x5 FILLER_199_640 ();
 b15zdnd11an1n64x5 FILLER_199_704 ();
 b15zdnd11an1n64x5 FILLER_199_768 ();
 b15zdnd11an1n64x5 FILLER_199_832 ();
 b15zdnd11an1n64x5 FILLER_199_896 ();
 b15zdnd11an1n64x5 FILLER_199_960 ();
 b15zdnd11an1n64x5 FILLER_199_1024 ();
 b15zdnd11an1n64x5 FILLER_199_1088 ();
 b15zdnd11an1n32x5 FILLER_199_1152 ();
 b15zdnd00an1n01x5 FILLER_199_1184 ();
 b15zdnd11an1n64x5 FILLER_199_1195 ();
 b15zdnd11an1n64x5 FILLER_199_1259 ();
 b15zdnd11an1n64x5 FILLER_199_1323 ();
 b15zdnd11an1n64x5 FILLER_199_1387 ();
 b15zdnd11an1n64x5 FILLER_199_1451 ();
 b15zdnd11an1n64x5 FILLER_199_1515 ();
 b15zdnd11an1n64x5 FILLER_199_1579 ();
 b15zdnd11an1n16x5 FILLER_199_1643 ();
 b15zdnd11an1n04x5 FILLER_199_1670 ();
 b15zdnd00an1n01x5 FILLER_199_1674 ();
 b15zdnd11an1n16x5 FILLER_199_1678 ();
 b15zdnd11an1n04x5 FILLER_199_1694 ();
 b15zdnd00an1n02x5 FILLER_199_1698 ();
 b15zdnd00an1n01x5 FILLER_199_1700 ();
 b15zdnd11an1n64x5 FILLER_199_1736 ();
 b15zdnd11an1n64x5 FILLER_199_1800 ();
 b15zdnd11an1n16x5 FILLER_199_1864 ();
 b15zdnd11an1n08x5 FILLER_199_1880 ();
 b15zdnd11an1n04x5 FILLER_199_1888 ();
 b15zdnd00an1n02x5 FILLER_199_1892 ();
 b15zdnd00an1n01x5 FILLER_199_1894 ();
 b15zdnd11an1n64x5 FILLER_199_1937 ();
 b15zdnd11an1n64x5 FILLER_199_2001 ();
 b15zdnd11an1n64x5 FILLER_199_2065 ();
 b15zdnd11an1n64x5 FILLER_199_2129 ();
 b15zdnd11an1n32x5 FILLER_199_2193 ();
 b15zdnd11an1n08x5 FILLER_199_2225 ();
 b15zdnd11an1n04x5 FILLER_199_2233 ();
 b15zdnd00an1n02x5 FILLER_199_2237 ();
 b15zdnd00an1n01x5 FILLER_199_2239 ();
 b15zdnd00an1n02x5 FILLER_199_2282 ();
 b15zdnd11an1n08x5 FILLER_200_8 ();
 b15zdnd11an1n04x5 FILLER_200_16 ();
 b15zdnd00an1n01x5 FILLER_200_20 ();
 b15zdnd11an1n64x5 FILLER_200_25 ();
 b15zdnd11an1n64x5 FILLER_200_89 ();
 b15zdnd11an1n64x5 FILLER_200_153 ();
 b15zdnd11an1n64x5 FILLER_200_217 ();
 b15zdnd11an1n64x5 FILLER_200_281 ();
 b15zdnd11an1n64x5 FILLER_200_345 ();
 b15zdnd11an1n64x5 FILLER_200_409 ();
 b15zdnd11an1n32x5 FILLER_200_473 ();
 b15zdnd11an1n16x5 FILLER_200_505 ();
 b15zdnd11an1n04x5 FILLER_200_521 ();
 b15zdnd00an1n02x5 FILLER_200_525 ();
 b15zdnd11an1n64x5 FILLER_200_538 ();
 b15zdnd11an1n64x5 FILLER_200_602 ();
 b15zdnd11an1n32x5 FILLER_200_666 ();
 b15zdnd11an1n16x5 FILLER_200_698 ();
 b15zdnd11an1n04x5 FILLER_200_714 ();
 b15zdnd11an1n64x5 FILLER_200_726 ();
 b15zdnd11an1n64x5 FILLER_200_790 ();
 b15zdnd11an1n64x5 FILLER_200_854 ();
 b15zdnd11an1n64x5 FILLER_200_918 ();
 b15zdnd11an1n64x5 FILLER_200_982 ();
 b15zdnd11an1n64x5 FILLER_200_1046 ();
 b15zdnd11an1n64x5 FILLER_200_1110 ();
 b15zdnd11an1n64x5 FILLER_200_1174 ();
 b15zdnd11an1n64x5 FILLER_200_1238 ();
 b15zdnd11an1n64x5 FILLER_200_1302 ();
 b15zdnd11an1n64x5 FILLER_200_1366 ();
 b15zdnd11an1n64x5 FILLER_200_1430 ();
 b15zdnd11an1n64x5 FILLER_200_1494 ();
 b15zdnd11an1n64x5 FILLER_200_1558 ();
 b15zdnd11an1n64x5 FILLER_200_1622 ();
 b15zdnd11an1n16x5 FILLER_200_1686 ();
 b15zdnd00an1n02x5 FILLER_200_1702 ();
 b15zdnd00an1n01x5 FILLER_200_1704 ();
 b15zdnd11an1n04x5 FILLER_200_1708 ();
 b15zdnd11an1n64x5 FILLER_200_1715 ();
 b15zdnd11an1n64x5 FILLER_200_1779 ();
 b15zdnd11an1n64x5 FILLER_200_1843 ();
 b15zdnd11an1n64x5 FILLER_200_1907 ();
 b15zdnd11an1n64x5 FILLER_200_1971 ();
 b15zdnd11an1n64x5 FILLER_200_2035 ();
 b15zdnd11an1n32x5 FILLER_200_2099 ();
 b15zdnd11an1n16x5 FILLER_200_2131 ();
 b15zdnd11an1n04x5 FILLER_200_2147 ();
 b15zdnd00an1n02x5 FILLER_200_2151 ();
 b15zdnd00an1n01x5 FILLER_200_2153 ();
 b15zdnd11an1n64x5 FILLER_200_2162 ();
 b15zdnd11an1n04x5 FILLER_200_2226 ();
 b15zdnd00an1n02x5 FILLER_200_2230 ();
 b15zdnd00an1n02x5 FILLER_200_2274 ();
 b15zdnd11an1n04x5 FILLER_201_0 ();
 b15zdnd00an1n02x5 FILLER_201_4 ();
 b15zdnd11an1n64x5 FILLER_201_48 ();
 b15zdnd11an1n64x5 FILLER_201_112 ();
 b15zdnd11an1n64x5 FILLER_201_176 ();
 b15zdnd11an1n64x5 FILLER_201_240 ();
 b15zdnd11an1n64x5 FILLER_201_304 ();
 b15zdnd11an1n64x5 FILLER_201_368 ();
 b15zdnd11an1n64x5 FILLER_201_432 ();
 b15zdnd11an1n64x5 FILLER_201_496 ();
 b15zdnd11an1n64x5 FILLER_201_560 ();
 b15zdnd11an1n32x5 FILLER_201_624 ();
 b15zdnd11an1n16x5 FILLER_201_656 ();
 b15zdnd11an1n04x5 FILLER_201_672 ();
 b15zdnd00an1n01x5 FILLER_201_676 ();
 b15zdnd11an1n64x5 FILLER_201_686 ();
 b15zdnd11an1n64x5 FILLER_201_750 ();
 b15zdnd11an1n64x5 FILLER_201_814 ();
 b15zdnd11an1n64x5 FILLER_201_878 ();
 b15zdnd11an1n32x5 FILLER_201_942 ();
 b15zdnd11an1n16x5 FILLER_201_974 ();
 b15zdnd00an1n02x5 FILLER_201_990 ();
 b15zdnd11an1n64x5 FILLER_201_1003 ();
 b15zdnd11an1n08x5 FILLER_201_1067 ();
 b15zdnd11an1n04x5 FILLER_201_1075 ();
 b15zdnd00an1n02x5 FILLER_201_1079 ();
 b15zdnd00an1n01x5 FILLER_201_1081 ();
 b15zdnd11an1n64x5 FILLER_201_1124 ();
 b15zdnd11an1n64x5 FILLER_201_1188 ();
 b15zdnd11an1n64x5 FILLER_201_1252 ();
 b15zdnd11an1n64x5 FILLER_201_1316 ();
 b15zdnd11an1n64x5 FILLER_201_1380 ();
 b15zdnd11an1n16x5 FILLER_201_1444 ();
 b15zdnd00an1n01x5 FILLER_201_1460 ();
 b15zdnd11an1n64x5 FILLER_201_1503 ();
 b15zdnd11an1n64x5 FILLER_201_1567 ();
 b15zdnd11an1n64x5 FILLER_201_1631 ();
 b15zdnd11an1n64x5 FILLER_201_1695 ();
 b15zdnd11an1n64x5 FILLER_201_1759 ();
 b15zdnd11an1n64x5 FILLER_201_1823 ();
 b15zdnd11an1n64x5 FILLER_201_1887 ();
 b15zdnd11an1n64x5 FILLER_201_1951 ();
 b15zdnd11an1n64x5 FILLER_201_2015 ();
 b15zdnd11an1n64x5 FILLER_201_2079 ();
 b15zdnd11an1n64x5 FILLER_201_2143 ();
 b15zdnd11an1n64x5 FILLER_201_2207 ();
 b15zdnd11an1n08x5 FILLER_201_2271 ();
 b15zdnd11an1n04x5 FILLER_201_2279 ();
 b15zdnd00an1n01x5 FILLER_201_2283 ();
 b15zdnd11an1n64x5 FILLER_202_8 ();
 b15zdnd11an1n64x5 FILLER_202_72 ();
 b15zdnd11an1n64x5 FILLER_202_136 ();
 b15zdnd11an1n64x5 FILLER_202_200 ();
 b15zdnd11an1n64x5 FILLER_202_264 ();
 b15zdnd11an1n64x5 FILLER_202_328 ();
 b15zdnd11an1n64x5 FILLER_202_392 ();
 b15zdnd11an1n64x5 FILLER_202_456 ();
 b15zdnd11an1n64x5 FILLER_202_520 ();
 b15zdnd11an1n64x5 FILLER_202_584 ();
 b15zdnd11an1n64x5 FILLER_202_648 ();
 b15zdnd11an1n04x5 FILLER_202_712 ();
 b15zdnd00an1n02x5 FILLER_202_716 ();
 b15zdnd11an1n64x5 FILLER_202_726 ();
 b15zdnd11an1n64x5 FILLER_202_790 ();
 b15zdnd11an1n64x5 FILLER_202_854 ();
 b15zdnd11an1n64x5 FILLER_202_918 ();
 b15zdnd11an1n64x5 FILLER_202_982 ();
 b15zdnd11an1n64x5 FILLER_202_1046 ();
 b15zdnd11an1n64x5 FILLER_202_1110 ();
 b15zdnd11an1n64x5 FILLER_202_1174 ();
 b15zdnd11an1n08x5 FILLER_202_1238 ();
 b15zdnd11an1n04x5 FILLER_202_1246 ();
 b15zdnd00an1n02x5 FILLER_202_1250 ();
 b15zdnd11an1n64x5 FILLER_202_1283 ();
 b15zdnd11an1n32x5 FILLER_202_1347 ();
 b15zdnd11an1n16x5 FILLER_202_1379 ();
 b15zdnd11an1n04x5 FILLER_202_1395 ();
 b15zdnd00an1n02x5 FILLER_202_1399 ();
 b15zdnd00an1n01x5 FILLER_202_1401 ();
 b15zdnd11an1n64x5 FILLER_202_1433 ();
 b15zdnd11an1n64x5 FILLER_202_1497 ();
 b15zdnd11an1n64x5 FILLER_202_1561 ();
 b15zdnd11an1n64x5 FILLER_202_1625 ();
 b15zdnd11an1n64x5 FILLER_202_1689 ();
 b15zdnd11an1n64x5 FILLER_202_1753 ();
 b15zdnd11an1n64x5 FILLER_202_1817 ();
 b15zdnd11an1n64x5 FILLER_202_1881 ();
 b15zdnd11an1n64x5 FILLER_202_1945 ();
 b15zdnd11an1n64x5 FILLER_202_2051 ();
 b15zdnd11an1n32x5 FILLER_202_2115 ();
 b15zdnd11an1n04x5 FILLER_202_2147 ();
 b15zdnd00an1n02x5 FILLER_202_2151 ();
 b15zdnd00an1n01x5 FILLER_202_2153 ();
 b15zdnd11an1n64x5 FILLER_202_2162 ();
 b15zdnd11an1n32x5 FILLER_202_2226 ();
 b15zdnd11an1n16x5 FILLER_202_2258 ();
 b15zdnd00an1n02x5 FILLER_202_2274 ();
 b15zdnd11an1n64x5 FILLER_203_0 ();
 b15zdnd11an1n64x5 FILLER_203_64 ();
 b15zdnd11an1n64x5 FILLER_203_128 ();
 b15zdnd11an1n64x5 FILLER_203_192 ();
 b15zdnd11an1n64x5 FILLER_203_256 ();
 b15zdnd11an1n64x5 FILLER_203_320 ();
 b15zdnd11an1n64x5 FILLER_203_384 ();
 b15zdnd11an1n64x5 FILLER_203_448 ();
 b15zdnd11an1n64x5 FILLER_203_512 ();
 b15zdnd11an1n64x5 FILLER_203_576 ();
 b15zdnd11an1n64x5 FILLER_203_640 ();
 b15zdnd11an1n64x5 FILLER_203_704 ();
 b15zdnd11an1n64x5 FILLER_203_768 ();
 b15zdnd11an1n64x5 FILLER_203_832 ();
 b15zdnd11an1n64x5 FILLER_203_896 ();
 b15zdnd11an1n64x5 FILLER_203_960 ();
 b15zdnd11an1n64x5 FILLER_203_1024 ();
 b15zdnd11an1n64x5 FILLER_203_1088 ();
 b15zdnd11an1n16x5 FILLER_203_1152 ();
 b15zdnd11an1n08x5 FILLER_203_1168 ();
 b15zdnd11an1n04x5 FILLER_203_1176 ();
 b15zdnd00an1n01x5 FILLER_203_1180 ();
 b15zdnd11an1n32x5 FILLER_203_1201 ();
 b15zdnd00an1n02x5 FILLER_203_1233 ();
 b15zdnd11an1n64x5 FILLER_203_1255 ();
 b15zdnd11an1n64x5 FILLER_203_1319 ();
 b15zdnd11an1n32x5 FILLER_203_1383 ();
 b15zdnd11an1n16x5 FILLER_203_1415 ();
 b15zdnd00an1n02x5 FILLER_203_1431 ();
 b15zdnd11an1n64x5 FILLER_203_1449 ();
 b15zdnd11an1n64x5 FILLER_203_1513 ();
 b15zdnd11an1n64x5 FILLER_203_1577 ();
 b15zdnd11an1n64x5 FILLER_203_1641 ();
 b15zdnd11an1n64x5 FILLER_203_1705 ();
 b15zdnd11an1n64x5 FILLER_203_1769 ();
 b15zdnd11an1n64x5 FILLER_203_1833 ();
 b15zdnd11an1n64x5 FILLER_203_1897 ();
 b15zdnd11an1n32x5 FILLER_203_1961 ();
 b15zdnd00an1n02x5 FILLER_203_1993 ();
 b15zdnd11an1n64x5 FILLER_203_2037 ();
 b15zdnd11an1n64x5 FILLER_203_2101 ();
 b15zdnd11an1n64x5 FILLER_203_2165 ();
 b15zdnd11an1n32x5 FILLER_203_2229 ();
 b15zdnd11an1n16x5 FILLER_203_2261 ();
 b15zdnd11an1n04x5 FILLER_203_2277 ();
 b15zdnd00an1n02x5 FILLER_203_2281 ();
 b15zdnd00an1n01x5 FILLER_203_2283 ();
 b15zdnd11an1n64x5 FILLER_204_8 ();
 b15zdnd11an1n64x5 FILLER_204_72 ();
 b15zdnd11an1n64x5 FILLER_204_136 ();
 b15zdnd11an1n64x5 FILLER_204_200 ();
 b15zdnd11an1n64x5 FILLER_204_264 ();
 b15zdnd11an1n64x5 FILLER_204_328 ();
 b15zdnd11an1n64x5 FILLER_204_392 ();
 b15zdnd11an1n64x5 FILLER_204_456 ();
 b15zdnd11an1n64x5 FILLER_204_520 ();
 b15zdnd11an1n64x5 FILLER_204_584 ();
 b15zdnd11an1n64x5 FILLER_204_648 ();
 b15zdnd11an1n04x5 FILLER_204_712 ();
 b15zdnd00an1n02x5 FILLER_204_716 ();
 b15zdnd11an1n64x5 FILLER_204_726 ();
 b15zdnd11an1n64x5 FILLER_204_790 ();
 b15zdnd11an1n32x5 FILLER_204_854 ();
 b15zdnd11an1n08x5 FILLER_204_886 ();
 b15zdnd11an1n64x5 FILLER_204_902 ();
 b15zdnd11an1n64x5 FILLER_204_966 ();
 b15zdnd11an1n64x5 FILLER_204_1030 ();
 b15zdnd11an1n64x5 FILLER_204_1094 ();
 b15zdnd11an1n32x5 FILLER_204_1158 ();
 b15zdnd11an1n16x5 FILLER_204_1190 ();
 b15zdnd11an1n08x5 FILLER_204_1206 ();
 b15zdnd11an1n04x5 FILLER_204_1214 ();
 b15zdnd00an1n01x5 FILLER_204_1218 ();
 b15zdnd11an1n32x5 FILLER_204_1239 ();
 b15zdnd11an1n16x5 FILLER_204_1271 ();
 b15zdnd11an1n08x5 FILLER_204_1287 ();
 b15zdnd00an1n02x5 FILLER_204_1295 ();
 b15zdnd00an1n01x5 FILLER_204_1297 ();
 b15zdnd11an1n64x5 FILLER_204_1314 ();
 b15zdnd11an1n64x5 FILLER_204_1378 ();
 b15zdnd11an1n64x5 FILLER_204_1442 ();
 b15zdnd11an1n64x5 FILLER_204_1506 ();
 b15zdnd11an1n64x5 FILLER_204_1570 ();
 b15zdnd11an1n64x5 FILLER_204_1634 ();
 b15zdnd11an1n64x5 FILLER_204_1698 ();
 b15zdnd11an1n64x5 FILLER_204_1762 ();
 b15zdnd11an1n64x5 FILLER_204_1826 ();
 b15zdnd11an1n64x5 FILLER_204_1890 ();
 b15zdnd11an1n64x5 FILLER_204_1954 ();
 b15zdnd11an1n64x5 FILLER_204_2018 ();
 b15zdnd11an1n64x5 FILLER_204_2082 ();
 b15zdnd11an1n08x5 FILLER_204_2146 ();
 b15zdnd11an1n64x5 FILLER_204_2162 ();
 b15zdnd11an1n32x5 FILLER_204_2226 ();
 b15zdnd11an1n16x5 FILLER_204_2258 ();
 b15zdnd00an1n02x5 FILLER_204_2274 ();
 b15zdnd11an1n64x5 FILLER_205_0 ();
 b15zdnd11an1n64x5 FILLER_205_64 ();
 b15zdnd11an1n64x5 FILLER_205_128 ();
 b15zdnd11an1n64x5 FILLER_205_192 ();
 b15zdnd11an1n64x5 FILLER_205_256 ();
 b15zdnd11an1n64x5 FILLER_205_320 ();
 b15zdnd11an1n64x5 FILLER_205_384 ();
 b15zdnd11an1n64x5 FILLER_205_448 ();
 b15zdnd11an1n64x5 FILLER_205_512 ();
 b15zdnd11an1n64x5 FILLER_205_576 ();
 b15zdnd11an1n64x5 FILLER_205_640 ();
 b15zdnd11an1n64x5 FILLER_205_704 ();
 b15zdnd11an1n64x5 FILLER_205_768 ();
 b15zdnd11an1n64x5 FILLER_205_832 ();
 b15zdnd11an1n64x5 FILLER_205_896 ();
 b15zdnd11an1n64x5 FILLER_205_960 ();
 b15zdnd11an1n64x5 FILLER_205_1024 ();
 b15zdnd11an1n64x5 FILLER_205_1088 ();
 b15zdnd11an1n32x5 FILLER_205_1152 ();
 b15zdnd00an1n01x5 FILLER_205_1184 ();
 b15zdnd11an1n16x5 FILLER_205_1196 ();
 b15zdnd00an1n02x5 FILLER_205_1212 ();
 b15zdnd11an1n08x5 FILLER_205_1240 ();
 b15zdnd11an1n04x5 FILLER_205_1248 ();
 b15zdnd00an1n01x5 FILLER_205_1252 ();
 b15zdnd11an1n64x5 FILLER_205_1267 ();
 b15zdnd11an1n64x5 FILLER_205_1331 ();
 b15zdnd11an1n64x5 FILLER_205_1395 ();
 b15zdnd11an1n64x5 FILLER_205_1459 ();
 b15zdnd11an1n64x5 FILLER_205_1523 ();
 b15zdnd11an1n64x5 FILLER_205_1587 ();
 b15zdnd11an1n64x5 FILLER_205_1651 ();
 b15zdnd11an1n64x5 FILLER_205_1715 ();
 b15zdnd11an1n64x5 FILLER_205_1779 ();
 b15zdnd11an1n64x5 FILLER_205_1843 ();
 b15zdnd11an1n64x5 FILLER_205_1907 ();
 b15zdnd11an1n64x5 FILLER_205_1971 ();
 b15zdnd11an1n64x5 FILLER_205_2035 ();
 b15zdnd11an1n64x5 FILLER_205_2099 ();
 b15zdnd11an1n64x5 FILLER_205_2163 ();
 b15zdnd11an1n16x5 FILLER_205_2227 ();
 b15zdnd11an1n04x5 FILLER_205_2243 ();
 b15zdnd11an1n32x5 FILLER_205_2252 ();
 b15zdnd11an1n64x5 FILLER_206_8 ();
 b15zdnd11an1n64x5 FILLER_206_72 ();
 b15zdnd11an1n64x5 FILLER_206_136 ();
 b15zdnd11an1n32x5 FILLER_206_200 ();
 b15zdnd11an1n16x5 FILLER_206_232 ();
 b15zdnd11an1n08x5 FILLER_206_248 ();
 b15zdnd11an1n04x5 FILLER_206_256 ();
 b15zdnd00an1n02x5 FILLER_206_260 ();
 b15zdnd00an1n01x5 FILLER_206_262 ();
 b15zdnd11an1n64x5 FILLER_206_271 ();
 b15zdnd11an1n64x5 FILLER_206_335 ();
 b15zdnd11an1n64x5 FILLER_206_399 ();
 b15zdnd11an1n64x5 FILLER_206_463 ();
 b15zdnd11an1n64x5 FILLER_206_527 ();
 b15zdnd11an1n16x5 FILLER_206_591 ();
 b15zdnd11an1n08x5 FILLER_206_607 ();
 b15zdnd00an1n02x5 FILLER_206_615 ();
 b15zdnd00an1n01x5 FILLER_206_617 ();
 b15zdnd11an1n64x5 FILLER_206_630 ();
 b15zdnd11an1n16x5 FILLER_206_694 ();
 b15zdnd11an1n08x5 FILLER_206_710 ();
 b15zdnd11an1n64x5 FILLER_206_726 ();
 b15zdnd11an1n64x5 FILLER_206_790 ();
 b15zdnd11an1n64x5 FILLER_206_854 ();
 b15zdnd11an1n64x5 FILLER_206_918 ();
 b15zdnd11an1n64x5 FILLER_206_982 ();
 b15zdnd11an1n64x5 FILLER_206_1046 ();
 b15zdnd11an1n64x5 FILLER_206_1110 ();
 b15zdnd11an1n08x5 FILLER_206_1174 ();
 b15zdnd11an1n04x5 FILLER_206_1182 ();
 b15zdnd00an1n02x5 FILLER_206_1186 ();
 b15zdnd00an1n01x5 FILLER_206_1188 ();
 b15zdnd11an1n32x5 FILLER_206_1198 ();
 b15zdnd11an1n16x5 FILLER_206_1230 ();
 b15zdnd00an1n01x5 FILLER_206_1246 ();
 b15zdnd11an1n64x5 FILLER_206_1278 ();
 b15zdnd11an1n32x5 FILLER_206_1342 ();
 b15zdnd11an1n04x5 FILLER_206_1374 ();
 b15zdnd11an1n64x5 FILLER_206_1409 ();
 b15zdnd11an1n64x5 FILLER_206_1473 ();
 b15zdnd11an1n64x5 FILLER_206_1537 ();
 b15zdnd11an1n64x5 FILLER_206_1601 ();
 b15zdnd11an1n64x5 FILLER_206_1665 ();
 b15zdnd11an1n64x5 FILLER_206_1729 ();
 b15zdnd11an1n64x5 FILLER_206_1793 ();
 b15zdnd11an1n64x5 FILLER_206_1857 ();
 b15zdnd11an1n64x5 FILLER_206_1921 ();
 b15zdnd11an1n64x5 FILLER_206_1985 ();
 b15zdnd11an1n64x5 FILLER_206_2049 ();
 b15zdnd11an1n32x5 FILLER_206_2113 ();
 b15zdnd11an1n08x5 FILLER_206_2145 ();
 b15zdnd00an1n01x5 FILLER_206_2153 ();
 b15zdnd11an1n64x5 FILLER_206_2162 ();
 b15zdnd11an1n32x5 FILLER_206_2226 ();
 b15zdnd11an1n04x5 FILLER_206_2263 ();
 b15zdnd11an1n04x5 FILLER_206_2272 ();
 b15zdnd11an1n64x5 FILLER_207_0 ();
 b15zdnd11an1n64x5 FILLER_207_64 ();
 b15zdnd11an1n64x5 FILLER_207_128 ();
 b15zdnd11an1n64x5 FILLER_207_192 ();
 b15zdnd11an1n64x5 FILLER_207_256 ();
 b15zdnd11an1n64x5 FILLER_207_320 ();
 b15zdnd11an1n64x5 FILLER_207_384 ();
 b15zdnd11an1n64x5 FILLER_207_448 ();
 b15zdnd11an1n64x5 FILLER_207_512 ();
 b15zdnd11an1n64x5 FILLER_207_576 ();
 b15zdnd11an1n16x5 FILLER_207_640 ();
 b15zdnd11an1n08x5 FILLER_207_656 ();
 b15zdnd00an1n02x5 FILLER_207_664 ();
 b15zdnd11an1n64x5 FILLER_207_686 ();
 b15zdnd11an1n64x5 FILLER_207_750 ();
 b15zdnd11an1n64x5 FILLER_207_814 ();
 b15zdnd11an1n64x5 FILLER_207_878 ();
 b15zdnd11an1n64x5 FILLER_207_942 ();
 b15zdnd11an1n64x5 FILLER_207_1006 ();
 b15zdnd11an1n64x5 FILLER_207_1070 ();
 b15zdnd11an1n64x5 FILLER_207_1134 ();
 b15zdnd11an1n04x5 FILLER_207_1198 ();
 b15zdnd00an1n02x5 FILLER_207_1202 ();
 b15zdnd11an1n16x5 FILLER_207_1220 ();
 b15zdnd11an1n08x5 FILLER_207_1236 ();
 b15zdnd00an1n01x5 FILLER_207_1244 ();
 b15zdnd11an1n64x5 FILLER_207_1271 ();
 b15zdnd11an1n64x5 FILLER_207_1335 ();
 b15zdnd11an1n64x5 FILLER_207_1399 ();
 b15zdnd11an1n64x5 FILLER_207_1463 ();
 b15zdnd11an1n16x5 FILLER_207_1527 ();
 b15zdnd00an1n02x5 FILLER_207_1543 ();
 b15zdnd11an1n64x5 FILLER_207_1587 ();
 b15zdnd11an1n64x5 FILLER_207_1651 ();
 b15zdnd11an1n64x5 FILLER_207_1715 ();
 b15zdnd11an1n64x5 FILLER_207_1779 ();
 b15zdnd11an1n64x5 FILLER_207_1843 ();
 b15zdnd11an1n64x5 FILLER_207_1907 ();
 b15zdnd11an1n64x5 FILLER_207_1971 ();
 b15zdnd11an1n64x5 FILLER_207_2035 ();
 b15zdnd11an1n64x5 FILLER_207_2099 ();
 b15zdnd11an1n64x5 FILLER_207_2163 ();
 b15zdnd11an1n08x5 FILLER_207_2227 ();
 b15zdnd11an1n04x5 FILLER_207_2235 ();
 b15zdnd00an1n02x5 FILLER_207_2239 ();
 b15zdnd11an1n04x5 FILLER_207_2246 ();
 b15zdnd11an1n08x5 FILLER_207_2255 ();
 b15zdnd11an1n04x5 FILLER_207_2263 ();
 b15zdnd00an1n02x5 FILLER_207_2267 ();
 b15zdnd11an1n04x5 FILLER_207_2277 ();
 b15zdnd00an1n02x5 FILLER_207_2281 ();
 b15zdnd00an1n01x5 FILLER_207_2283 ();
 b15zdnd11an1n64x5 FILLER_208_8 ();
 b15zdnd11an1n64x5 FILLER_208_72 ();
 b15zdnd11an1n64x5 FILLER_208_136 ();
 b15zdnd11an1n64x5 FILLER_208_200 ();
 b15zdnd11an1n64x5 FILLER_208_264 ();
 b15zdnd11an1n08x5 FILLER_208_328 ();
 b15zdnd11an1n04x5 FILLER_208_336 ();
 b15zdnd00an1n02x5 FILLER_208_340 ();
 b15zdnd11an1n64x5 FILLER_208_384 ();
 b15zdnd11an1n64x5 FILLER_208_448 ();
 b15zdnd11an1n64x5 FILLER_208_512 ();
 b15zdnd11an1n64x5 FILLER_208_576 ();
 b15zdnd11an1n64x5 FILLER_208_640 ();
 b15zdnd11an1n08x5 FILLER_208_704 ();
 b15zdnd11an1n04x5 FILLER_208_712 ();
 b15zdnd00an1n02x5 FILLER_208_716 ();
 b15zdnd11an1n64x5 FILLER_208_726 ();
 b15zdnd11an1n32x5 FILLER_208_790 ();
 b15zdnd11an1n08x5 FILLER_208_822 ();
 b15zdnd00an1n01x5 FILLER_208_830 ();
 b15zdnd11an1n64x5 FILLER_208_850 ();
 b15zdnd11an1n64x5 FILLER_208_914 ();
 b15zdnd11an1n64x5 FILLER_208_978 ();
 b15zdnd11an1n64x5 FILLER_208_1042 ();
 b15zdnd11an1n64x5 FILLER_208_1106 ();
 b15zdnd11an1n64x5 FILLER_208_1170 ();
 b15zdnd11an1n64x5 FILLER_208_1234 ();
 b15zdnd11an1n64x5 FILLER_208_1298 ();
 b15zdnd11an1n64x5 FILLER_208_1362 ();
 b15zdnd11an1n64x5 FILLER_208_1426 ();
 b15zdnd11an1n32x5 FILLER_208_1490 ();
 b15zdnd11an1n16x5 FILLER_208_1522 ();
 b15zdnd11an1n08x5 FILLER_208_1538 ();
 b15zdnd00an1n01x5 FILLER_208_1546 ();
 b15zdnd11an1n64x5 FILLER_208_1589 ();
 b15zdnd11an1n64x5 FILLER_208_1653 ();
 b15zdnd11an1n64x5 FILLER_208_1717 ();
 b15zdnd11an1n64x5 FILLER_208_1781 ();
 b15zdnd11an1n64x5 FILLER_208_1845 ();
 b15zdnd11an1n64x5 FILLER_208_1909 ();
 b15zdnd11an1n64x5 FILLER_208_1973 ();
 b15zdnd11an1n64x5 FILLER_208_2037 ();
 b15zdnd11an1n32x5 FILLER_208_2101 ();
 b15zdnd11an1n16x5 FILLER_208_2133 ();
 b15zdnd11an1n04x5 FILLER_208_2149 ();
 b15zdnd00an1n01x5 FILLER_208_2153 ();
 b15zdnd11an1n64x5 FILLER_208_2162 ();
 b15zdnd11an1n32x5 FILLER_208_2226 ();
 b15zdnd11an1n08x5 FILLER_208_2258 ();
 b15zdnd11an1n04x5 FILLER_208_2271 ();
 b15zdnd00an1n01x5 FILLER_208_2275 ();
 b15zdnd11an1n64x5 FILLER_209_0 ();
 b15zdnd11an1n64x5 FILLER_209_64 ();
 b15zdnd11an1n64x5 FILLER_209_128 ();
 b15zdnd11an1n64x5 FILLER_209_192 ();
 b15zdnd11an1n64x5 FILLER_209_256 ();
 b15zdnd11an1n16x5 FILLER_209_320 ();
 b15zdnd11an1n08x5 FILLER_209_336 ();
 b15zdnd11an1n64x5 FILLER_209_386 ();
 b15zdnd11an1n64x5 FILLER_209_450 ();
 b15zdnd11an1n64x5 FILLER_209_514 ();
 b15zdnd11an1n64x5 FILLER_209_578 ();
 b15zdnd11an1n64x5 FILLER_209_642 ();
 b15zdnd11an1n64x5 FILLER_209_706 ();
 b15zdnd11an1n64x5 FILLER_209_770 ();
 b15zdnd11an1n64x5 FILLER_209_834 ();
 b15zdnd11an1n64x5 FILLER_209_898 ();
 b15zdnd11an1n64x5 FILLER_209_962 ();
 b15zdnd11an1n64x5 FILLER_209_1026 ();
 b15zdnd11an1n64x5 FILLER_209_1090 ();
 b15zdnd11an1n64x5 FILLER_209_1154 ();
 b15zdnd11an1n64x5 FILLER_209_1218 ();
 b15zdnd11an1n64x5 FILLER_209_1282 ();
 b15zdnd11an1n64x5 FILLER_209_1346 ();
 b15zdnd11an1n64x5 FILLER_209_1410 ();
 b15zdnd11an1n64x5 FILLER_209_1474 ();
 b15zdnd11an1n64x5 FILLER_209_1538 ();
 b15zdnd11an1n64x5 FILLER_209_1602 ();
 b15zdnd11an1n64x5 FILLER_209_1666 ();
 b15zdnd11an1n64x5 FILLER_209_1730 ();
 b15zdnd11an1n64x5 FILLER_209_1794 ();
 b15zdnd11an1n64x5 FILLER_209_1858 ();
 b15zdnd11an1n64x5 FILLER_209_1922 ();
 b15zdnd11an1n64x5 FILLER_209_1986 ();
 b15zdnd11an1n64x5 FILLER_209_2050 ();
 b15zdnd11an1n64x5 FILLER_209_2114 ();
 b15zdnd11an1n64x5 FILLER_209_2178 ();
 b15zdnd11an1n08x5 FILLER_209_2242 ();
 b15zdnd11an1n04x5 FILLER_209_2250 ();
 b15zdnd00an1n01x5 FILLER_209_2254 ();
 b15zdnd11an1n16x5 FILLER_209_2260 ();
 b15zdnd11an1n08x5 FILLER_209_2276 ();
 b15zdnd11an1n64x5 FILLER_210_8 ();
 b15zdnd11an1n64x5 FILLER_210_72 ();
 b15zdnd11an1n64x5 FILLER_210_136 ();
 b15zdnd11an1n64x5 FILLER_210_200 ();
 b15zdnd11an1n64x5 FILLER_210_264 ();
 b15zdnd11an1n64x5 FILLER_210_328 ();
 b15zdnd11an1n64x5 FILLER_210_392 ();
 b15zdnd11an1n64x5 FILLER_210_456 ();
 b15zdnd11an1n64x5 FILLER_210_520 ();
 b15zdnd11an1n16x5 FILLER_210_584 ();
 b15zdnd11an1n08x5 FILLER_210_600 ();
 b15zdnd11an1n64x5 FILLER_210_650 ();
 b15zdnd11an1n04x5 FILLER_210_714 ();
 b15zdnd11an1n64x5 FILLER_210_726 ();
 b15zdnd11an1n64x5 FILLER_210_790 ();
 b15zdnd11an1n32x5 FILLER_210_854 ();
 b15zdnd00an1n02x5 FILLER_210_886 ();
 b15zdnd00an1n01x5 FILLER_210_888 ();
 b15zdnd11an1n64x5 FILLER_210_912 ();
 b15zdnd11an1n64x5 FILLER_210_976 ();
 b15zdnd11an1n64x5 FILLER_210_1040 ();
 b15zdnd11an1n64x5 FILLER_210_1104 ();
 b15zdnd11an1n64x5 FILLER_210_1168 ();
 b15zdnd11an1n64x5 FILLER_210_1232 ();
 b15zdnd11an1n64x5 FILLER_210_1296 ();
 b15zdnd11an1n64x5 FILLER_210_1360 ();
 b15zdnd11an1n64x5 FILLER_210_1424 ();
 b15zdnd11an1n64x5 FILLER_210_1488 ();
 b15zdnd11an1n64x5 FILLER_210_1552 ();
 b15zdnd11an1n64x5 FILLER_210_1616 ();
 b15zdnd11an1n64x5 FILLER_210_1680 ();
 b15zdnd11an1n64x5 FILLER_210_1744 ();
 b15zdnd11an1n64x5 FILLER_210_1808 ();
 b15zdnd11an1n64x5 FILLER_210_1872 ();
 b15zdnd11an1n64x5 FILLER_210_1936 ();
 b15zdnd11an1n64x5 FILLER_210_2000 ();
 b15zdnd11an1n64x5 FILLER_210_2064 ();
 b15zdnd11an1n16x5 FILLER_210_2128 ();
 b15zdnd11an1n08x5 FILLER_210_2144 ();
 b15zdnd00an1n02x5 FILLER_210_2152 ();
 b15zdnd11an1n64x5 FILLER_210_2162 ();
 b15zdnd11an1n32x5 FILLER_210_2226 ();
 b15zdnd11an1n16x5 FILLER_210_2258 ();
 b15zdnd00an1n02x5 FILLER_210_2274 ();
 b15zdnd11an1n64x5 FILLER_211_0 ();
 b15zdnd11an1n64x5 FILLER_211_64 ();
 b15zdnd11an1n64x5 FILLER_211_128 ();
 b15zdnd11an1n64x5 FILLER_211_192 ();
 b15zdnd11an1n64x5 FILLER_211_256 ();
 b15zdnd11an1n16x5 FILLER_211_320 ();
 b15zdnd00an1n02x5 FILLER_211_336 ();
 b15zdnd11an1n64x5 FILLER_211_380 ();
 b15zdnd11an1n64x5 FILLER_211_444 ();
 b15zdnd11an1n64x5 FILLER_211_508 ();
 b15zdnd11an1n64x5 FILLER_211_572 ();
 b15zdnd11an1n64x5 FILLER_211_636 ();
 b15zdnd11an1n64x5 FILLER_211_700 ();
 b15zdnd11an1n64x5 FILLER_211_764 ();
 b15zdnd11an1n32x5 FILLER_211_828 ();
 b15zdnd11an1n16x5 FILLER_211_860 ();
 b15zdnd11an1n08x5 FILLER_211_876 ();
 b15zdnd00an1n02x5 FILLER_211_884 ();
 b15zdnd11an1n32x5 FILLER_211_890 ();
 b15zdnd11an1n16x5 FILLER_211_922 ();
 b15zdnd00an1n02x5 FILLER_211_938 ();
 b15zdnd00an1n01x5 FILLER_211_940 ();
 b15zdnd11an1n64x5 FILLER_211_959 ();
 b15zdnd11an1n32x5 FILLER_211_1023 ();
 b15zdnd11an1n16x5 FILLER_211_1055 ();
 b15zdnd11an1n08x5 FILLER_211_1071 ();
 b15zdnd11an1n04x5 FILLER_211_1079 ();
 b15zdnd00an1n02x5 FILLER_211_1083 ();
 b15zdnd00an1n01x5 FILLER_211_1085 ();
 b15zdnd11an1n64x5 FILLER_211_1105 ();
 b15zdnd11an1n64x5 FILLER_211_1169 ();
 b15zdnd11an1n64x5 FILLER_211_1233 ();
 b15zdnd11an1n64x5 FILLER_211_1297 ();
 b15zdnd11an1n64x5 FILLER_211_1361 ();
 b15zdnd11an1n64x5 FILLER_211_1425 ();
 b15zdnd11an1n64x5 FILLER_211_1489 ();
 b15zdnd11an1n64x5 FILLER_211_1553 ();
 b15zdnd11an1n64x5 FILLER_211_1617 ();
 b15zdnd11an1n64x5 FILLER_211_1681 ();
 b15zdnd11an1n08x5 FILLER_211_1745 ();
 b15zdnd11an1n64x5 FILLER_211_1795 ();
 b15zdnd11an1n64x5 FILLER_211_1859 ();
 b15zdnd11an1n64x5 FILLER_211_1923 ();
 b15zdnd11an1n64x5 FILLER_211_1987 ();
 b15zdnd11an1n64x5 FILLER_211_2051 ();
 b15zdnd11an1n64x5 FILLER_211_2115 ();
 b15zdnd11an1n64x5 FILLER_211_2179 ();
 b15zdnd11an1n32x5 FILLER_211_2243 ();
 b15zdnd11an1n08x5 FILLER_211_2275 ();
 b15zdnd00an1n01x5 FILLER_211_2283 ();
 b15zdnd11an1n64x5 FILLER_212_8 ();
 b15zdnd11an1n64x5 FILLER_212_72 ();
 b15zdnd11an1n64x5 FILLER_212_136 ();
 b15zdnd11an1n64x5 FILLER_212_200 ();
 b15zdnd11an1n64x5 FILLER_212_264 ();
 b15zdnd11an1n64x5 FILLER_212_328 ();
 b15zdnd11an1n64x5 FILLER_212_392 ();
 b15zdnd11an1n64x5 FILLER_212_456 ();
 b15zdnd11an1n64x5 FILLER_212_520 ();
 b15zdnd11an1n64x5 FILLER_212_584 ();
 b15zdnd11an1n64x5 FILLER_212_648 ();
 b15zdnd11an1n04x5 FILLER_212_712 ();
 b15zdnd00an1n02x5 FILLER_212_716 ();
 b15zdnd11an1n64x5 FILLER_212_726 ();
 b15zdnd11an1n64x5 FILLER_212_790 ();
 b15zdnd11an1n64x5 FILLER_212_854 ();
 b15zdnd11an1n64x5 FILLER_212_918 ();
 b15zdnd11an1n64x5 FILLER_212_982 ();
 b15zdnd11an1n64x5 FILLER_212_1046 ();
 b15zdnd11an1n32x5 FILLER_212_1110 ();
 b15zdnd11an1n08x5 FILLER_212_1142 ();
 b15zdnd11an1n32x5 FILLER_212_1164 ();
 b15zdnd11an1n16x5 FILLER_212_1196 ();
 b15zdnd00an1n02x5 FILLER_212_1212 ();
 b15zdnd11an1n64x5 FILLER_212_1226 ();
 b15zdnd11an1n64x5 FILLER_212_1290 ();
 b15zdnd11an1n64x5 FILLER_212_1354 ();
 b15zdnd11an1n64x5 FILLER_212_1418 ();
 b15zdnd11an1n64x5 FILLER_212_1482 ();
 b15zdnd11an1n64x5 FILLER_212_1546 ();
 b15zdnd11an1n32x5 FILLER_212_1610 ();
 b15zdnd11an1n16x5 FILLER_212_1642 ();
 b15zdnd11an1n08x5 FILLER_212_1658 ();
 b15zdnd11an1n04x5 FILLER_212_1666 ();
 b15zdnd00an1n01x5 FILLER_212_1670 ();
 b15zdnd11an1n64x5 FILLER_212_1713 ();
 b15zdnd11an1n64x5 FILLER_212_1777 ();
 b15zdnd11an1n64x5 FILLER_212_1841 ();
 b15zdnd11an1n64x5 FILLER_212_1905 ();
 b15zdnd11an1n64x5 FILLER_212_1969 ();
 b15zdnd11an1n64x5 FILLER_212_2033 ();
 b15zdnd11an1n32x5 FILLER_212_2097 ();
 b15zdnd11an1n16x5 FILLER_212_2129 ();
 b15zdnd11an1n08x5 FILLER_212_2145 ();
 b15zdnd00an1n01x5 FILLER_212_2153 ();
 b15zdnd11an1n64x5 FILLER_212_2162 ();
 b15zdnd11an1n32x5 FILLER_212_2226 ();
 b15zdnd11an1n16x5 FILLER_212_2258 ();
 b15zdnd00an1n02x5 FILLER_212_2274 ();
 b15zdnd11an1n64x5 FILLER_213_0 ();
 b15zdnd11an1n64x5 FILLER_213_64 ();
 b15zdnd11an1n64x5 FILLER_213_128 ();
 b15zdnd11an1n64x5 FILLER_213_192 ();
 b15zdnd11an1n64x5 FILLER_213_256 ();
 b15zdnd11an1n64x5 FILLER_213_320 ();
 b15zdnd11an1n64x5 FILLER_213_384 ();
 b15zdnd11an1n64x5 FILLER_213_448 ();
 b15zdnd11an1n64x5 FILLER_213_512 ();
 b15zdnd11an1n64x5 FILLER_213_576 ();
 b15zdnd11an1n64x5 FILLER_213_640 ();
 b15zdnd11an1n64x5 FILLER_213_704 ();
 b15zdnd11an1n64x5 FILLER_213_768 ();
 b15zdnd11an1n64x5 FILLER_213_832 ();
 b15zdnd11an1n64x5 FILLER_213_896 ();
 b15zdnd11an1n64x5 FILLER_213_960 ();
 b15zdnd11an1n64x5 FILLER_213_1024 ();
 b15zdnd11an1n64x5 FILLER_213_1088 ();
 b15zdnd11an1n64x5 FILLER_213_1152 ();
 b15zdnd11an1n64x5 FILLER_213_1216 ();
 b15zdnd11an1n64x5 FILLER_213_1280 ();
 b15zdnd11an1n32x5 FILLER_213_1344 ();
 b15zdnd11an1n04x5 FILLER_213_1376 ();
 b15zdnd11an1n64x5 FILLER_213_1422 ();
 b15zdnd11an1n64x5 FILLER_213_1486 ();
 b15zdnd11an1n64x5 FILLER_213_1550 ();
 b15zdnd11an1n64x5 FILLER_213_1614 ();
 b15zdnd11an1n32x5 FILLER_213_1678 ();
 b15zdnd11an1n16x5 FILLER_213_1710 ();
 b15zdnd11an1n64x5 FILLER_213_1768 ();
 b15zdnd11an1n64x5 FILLER_213_1832 ();
 b15zdnd11an1n64x5 FILLER_213_1896 ();
 b15zdnd11an1n64x5 FILLER_213_1960 ();
 b15zdnd11an1n64x5 FILLER_213_2024 ();
 b15zdnd11an1n64x5 FILLER_213_2088 ();
 b15zdnd11an1n64x5 FILLER_213_2152 ();
 b15zdnd11an1n64x5 FILLER_213_2216 ();
 b15zdnd11an1n04x5 FILLER_213_2280 ();
 b15zdnd11an1n64x5 FILLER_214_8 ();
 b15zdnd11an1n64x5 FILLER_214_72 ();
 b15zdnd11an1n64x5 FILLER_214_136 ();
 b15zdnd11an1n64x5 FILLER_214_200 ();
 b15zdnd11an1n64x5 FILLER_214_264 ();
 b15zdnd11an1n64x5 FILLER_214_328 ();
 b15zdnd11an1n64x5 FILLER_214_392 ();
 b15zdnd11an1n64x5 FILLER_214_456 ();
 b15zdnd11an1n64x5 FILLER_214_520 ();
 b15zdnd11an1n64x5 FILLER_214_584 ();
 b15zdnd11an1n64x5 FILLER_214_648 ();
 b15zdnd11an1n04x5 FILLER_214_712 ();
 b15zdnd00an1n02x5 FILLER_214_716 ();
 b15zdnd11an1n64x5 FILLER_214_726 ();
 b15zdnd11an1n32x5 FILLER_214_790 ();
 b15zdnd11an1n16x5 FILLER_214_822 ();
 b15zdnd11an1n08x5 FILLER_214_838 ();
 b15zdnd00an1n02x5 FILLER_214_846 ();
 b15zdnd00an1n01x5 FILLER_214_848 ();
 b15zdnd11an1n64x5 FILLER_214_870 ();
 b15zdnd11an1n64x5 FILLER_214_934 ();
 b15zdnd11an1n64x5 FILLER_214_998 ();
 b15zdnd11an1n64x5 FILLER_214_1062 ();
 b15zdnd11an1n64x5 FILLER_214_1126 ();
 b15zdnd11an1n64x5 FILLER_214_1190 ();
 b15zdnd11an1n64x5 FILLER_214_1254 ();
 b15zdnd11an1n64x5 FILLER_214_1318 ();
 b15zdnd11an1n64x5 FILLER_214_1382 ();
 b15zdnd11an1n32x5 FILLER_214_1446 ();
 b15zdnd11an1n16x5 FILLER_214_1478 ();
 b15zdnd11an1n64x5 FILLER_214_1536 ();
 b15zdnd11an1n64x5 FILLER_214_1600 ();
 b15zdnd11an1n64x5 FILLER_214_1664 ();
 b15zdnd11an1n64x5 FILLER_214_1728 ();
 b15zdnd11an1n64x5 FILLER_214_1792 ();
 b15zdnd11an1n64x5 FILLER_214_1856 ();
 b15zdnd11an1n64x5 FILLER_214_1920 ();
 b15zdnd11an1n64x5 FILLER_214_1984 ();
 b15zdnd11an1n64x5 FILLER_214_2048 ();
 b15zdnd11an1n32x5 FILLER_214_2112 ();
 b15zdnd11an1n08x5 FILLER_214_2144 ();
 b15zdnd00an1n02x5 FILLER_214_2152 ();
 b15zdnd11an1n64x5 FILLER_214_2162 ();
 b15zdnd11an1n32x5 FILLER_214_2226 ();
 b15zdnd11an1n16x5 FILLER_214_2258 ();
 b15zdnd00an1n02x5 FILLER_214_2274 ();
 b15zdnd11an1n64x5 FILLER_215_0 ();
 b15zdnd11an1n64x5 FILLER_215_64 ();
 b15zdnd11an1n64x5 FILLER_215_128 ();
 b15zdnd11an1n64x5 FILLER_215_192 ();
 b15zdnd11an1n64x5 FILLER_215_256 ();
 b15zdnd11an1n64x5 FILLER_215_320 ();
 b15zdnd11an1n64x5 FILLER_215_384 ();
 b15zdnd11an1n64x5 FILLER_215_448 ();
 b15zdnd11an1n64x5 FILLER_215_512 ();
 b15zdnd11an1n64x5 FILLER_215_576 ();
 b15zdnd11an1n64x5 FILLER_215_640 ();
 b15zdnd11an1n64x5 FILLER_215_704 ();
 b15zdnd11an1n64x5 FILLER_215_768 ();
 b15zdnd11an1n64x5 FILLER_215_832 ();
 b15zdnd11an1n64x5 FILLER_215_896 ();
 b15zdnd11an1n16x5 FILLER_215_960 ();
 b15zdnd11an1n64x5 FILLER_215_995 ();
 b15zdnd11an1n64x5 FILLER_215_1059 ();
 b15zdnd11an1n64x5 FILLER_215_1123 ();
 b15zdnd11an1n16x5 FILLER_215_1187 ();
 b15zdnd11an1n08x5 FILLER_215_1203 ();
 b15zdnd11an1n04x5 FILLER_215_1211 ();
 b15zdnd00an1n02x5 FILLER_215_1215 ();
 b15zdnd11an1n64x5 FILLER_215_1237 ();
 b15zdnd11an1n64x5 FILLER_215_1301 ();
 b15zdnd11an1n64x5 FILLER_215_1365 ();
 b15zdnd11an1n64x5 FILLER_215_1429 ();
 b15zdnd11an1n64x5 FILLER_215_1493 ();
 b15zdnd11an1n64x5 FILLER_215_1557 ();
 b15zdnd11an1n32x5 FILLER_215_1621 ();
 b15zdnd11an1n64x5 FILLER_215_1695 ();
 b15zdnd11an1n64x5 FILLER_215_1759 ();
 b15zdnd11an1n64x5 FILLER_215_1823 ();
 b15zdnd11an1n64x5 FILLER_215_1887 ();
 b15zdnd11an1n64x5 FILLER_215_1951 ();
 b15zdnd11an1n64x5 FILLER_215_2015 ();
 b15zdnd11an1n64x5 FILLER_215_2079 ();
 b15zdnd11an1n16x5 FILLER_215_2143 ();
 b15zdnd11an1n64x5 FILLER_215_2175 ();
 b15zdnd11an1n32x5 FILLER_215_2239 ();
 b15zdnd11an1n08x5 FILLER_215_2271 ();
 b15zdnd11an1n04x5 FILLER_215_2279 ();
 b15zdnd00an1n01x5 FILLER_215_2283 ();
 b15zdnd11an1n64x5 FILLER_216_8 ();
 b15zdnd11an1n64x5 FILLER_216_72 ();
 b15zdnd11an1n64x5 FILLER_216_136 ();
 b15zdnd11an1n64x5 FILLER_216_200 ();
 b15zdnd11an1n64x5 FILLER_216_264 ();
 b15zdnd11an1n64x5 FILLER_216_328 ();
 b15zdnd11an1n64x5 FILLER_216_392 ();
 b15zdnd11an1n64x5 FILLER_216_456 ();
 b15zdnd11an1n64x5 FILLER_216_520 ();
 b15zdnd11an1n64x5 FILLER_216_584 ();
 b15zdnd11an1n64x5 FILLER_216_648 ();
 b15zdnd11an1n04x5 FILLER_216_712 ();
 b15zdnd00an1n02x5 FILLER_216_716 ();
 b15zdnd11an1n64x5 FILLER_216_726 ();
 b15zdnd11an1n16x5 FILLER_216_790 ();
 b15zdnd00an1n02x5 FILLER_216_806 ();
 b15zdnd00an1n01x5 FILLER_216_808 ();
 b15zdnd11an1n64x5 FILLER_216_851 ();
 b15zdnd11an1n64x5 FILLER_216_915 ();
 b15zdnd11an1n64x5 FILLER_216_979 ();
 b15zdnd11an1n64x5 FILLER_216_1043 ();
 b15zdnd11an1n64x5 FILLER_216_1107 ();
 b15zdnd11an1n64x5 FILLER_216_1171 ();
 b15zdnd11an1n64x5 FILLER_216_1235 ();
 b15zdnd11an1n64x5 FILLER_216_1299 ();
 b15zdnd11an1n64x5 FILLER_216_1363 ();
 b15zdnd11an1n64x5 FILLER_216_1427 ();
 b15zdnd11an1n64x5 FILLER_216_1491 ();
 b15zdnd11an1n64x5 FILLER_216_1555 ();
 b15zdnd11an1n64x5 FILLER_216_1619 ();
 b15zdnd11an1n64x5 FILLER_216_1683 ();
 b15zdnd11an1n64x5 FILLER_216_1747 ();
 b15zdnd11an1n64x5 FILLER_216_1811 ();
 b15zdnd11an1n64x5 FILLER_216_1875 ();
 b15zdnd11an1n64x5 FILLER_216_1939 ();
 b15zdnd11an1n64x5 FILLER_216_2003 ();
 b15zdnd11an1n64x5 FILLER_216_2067 ();
 b15zdnd11an1n16x5 FILLER_216_2131 ();
 b15zdnd11an1n04x5 FILLER_216_2147 ();
 b15zdnd00an1n02x5 FILLER_216_2151 ();
 b15zdnd00an1n01x5 FILLER_216_2153 ();
 b15zdnd11an1n64x5 FILLER_216_2162 ();
 b15zdnd11an1n32x5 FILLER_216_2226 ();
 b15zdnd11an1n16x5 FILLER_216_2258 ();
 b15zdnd00an1n02x5 FILLER_216_2274 ();
 b15zdnd11an1n64x5 FILLER_217_0 ();
 b15zdnd11an1n64x5 FILLER_217_64 ();
 b15zdnd11an1n64x5 FILLER_217_128 ();
 b15zdnd11an1n64x5 FILLER_217_192 ();
 b15zdnd11an1n64x5 FILLER_217_256 ();
 b15zdnd11an1n64x5 FILLER_217_320 ();
 b15zdnd11an1n64x5 FILLER_217_384 ();
 b15zdnd11an1n64x5 FILLER_217_448 ();
 b15zdnd11an1n64x5 FILLER_217_512 ();
 b15zdnd11an1n64x5 FILLER_217_576 ();
 b15zdnd11an1n32x5 FILLER_217_640 ();
 b15zdnd11an1n08x5 FILLER_217_672 ();
 b15zdnd00an1n02x5 FILLER_217_680 ();
 b15zdnd11an1n04x5 FILLER_217_694 ();
 b15zdnd00an1n01x5 FILLER_217_698 ();
 b15zdnd11an1n64x5 FILLER_217_741 ();
 b15zdnd11an1n64x5 FILLER_217_805 ();
 b15zdnd11an1n16x5 FILLER_217_869 ();
 b15zdnd11an1n08x5 FILLER_217_885 ();
 b15zdnd11an1n32x5 FILLER_217_935 ();
 b15zdnd11an1n16x5 FILLER_217_967 ();
 b15zdnd11an1n08x5 FILLER_217_983 ();
 b15zdnd00an1n02x5 FILLER_217_991 ();
 b15zdnd00an1n01x5 FILLER_217_993 ();
 b15zdnd11an1n64x5 FILLER_217_1013 ();
 b15zdnd11an1n64x5 FILLER_217_1077 ();
 b15zdnd11an1n64x5 FILLER_217_1141 ();
 b15zdnd11an1n64x5 FILLER_217_1205 ();
 b15zdnd11an1n64x5 FILLER_217_1269 ();
 b15zdnd11an1n64x5 FILLER_217_1333 ();
 b15zdnd11an1n64x5 FILLER_217_1397 ();
 b15zdnd11an1n64x5 FILLER_217_1461 ();
 b15zdnd11an1n64x5 FILLER_217_1525 ();
 b15zdnd11an1n64x5 FILLER_217_1589 ();
 b15zdnd11an1n64x5 FILLER_217_1653 ();
 b15zdnd11an1n64x5 FILLER_217_1717 ();
 b15zdnd11an1n64x5 FILLER_217_1781 ();
 b15zdnd11an1n64x5 FILLER_217_1845 ();
 b15zdnd11an1n64x5 FILLER_217_1909 ();
 b15zdnd11an1n64x5 FILLER_217_1973 ();
 b15zdnd11an1n64x5 FILLER_217_2037 ();
 b15zdnd11an1n64x5 FILLER_217_2101 ();
 b15zdnd11an1n64x5 FILLER_217_2165 ();
 b15zdnd11an1n32x5 FILLER_217_2229 ();
 b15zdnd11an1n16x5 FILLER_217_2261 ();
 b15zdnd11an1n04x5 FILLER_217_2277 ();
 b15zdnd00an1n02x5 FILLER_217_2281 ();
 b15zdnd00an1n01x5 FILLER_217_2283 ();
 b15zdnd11an1n64x5 FILLER_218_8 ();
 b15zdnd11an1n64x5 FILLER_218_72 ();
 b15zdnd11an1n64x5 FILLER_218_136 ();
 b15zdnd11an1n64x5 FILLER_218_200 ();
 b15zdnd11an1n64x5 FILLER_218_264 ();
 b15zdnd11an1n64x5 FILLER_218_328 ();
 b15zdnd11an1n64x5 FILLER_218_392 ();
 b15zdnd11an1n64x5 FILLER_218_456 ();
 b15zdnd11an1n64x5 FILLER_218_520 ();
 b15zdnd11an1n16x5 FILLER_218_584 ();
 b15zdnd11an1n04x5 FILLER_218_600 ();
 b15zdnd11an1n32x5 FILLER_218_620 ();
 b15zdnd00an1n02x5 FILLER_218_652 ();
 b15zdnd11an1n04x5 FILLER_218_668 ();
 b15zdnd11an1n08x5 FILLER_218_693 ();
 b15zdnd00an1n02x5 FILLER_218_701 ();
 b15zdnd00an1n01x5 FILLER_218_703 ();
 b15zdnd00an1n02x5 FILLER_218_716 ();
 b15zdnd11an1n64x5 FILLER_218_726 ();
 b15zdnd11an1n64x5 FILLER_218_790 ();
 b15zdnd11an1n64x5 FILLER_218_854 ();
 b15zdnd11an1n64x5 FILLER_218_918 ();
 b15zdnd11an1n04x5 FILLER_218_982 ();
 b15zdnd00an1n02x5 FILLER_218_986 ();
 b15zdnd00an1n01x5 FILLER_218_988 ();
 b15zdnd11an1n64x5 FILLER_218_1008 ();
 b15zdnd11an1n64x5 FILLER_218_1072 ();
 b15zdnd11an1n64x5 FILLER_218_1136 ();
 b15zdnd11an1n64x5 FILLER_218_1200 ();
 b15zdnd11an1n64x5 FILLER_218_1264 ();
 b15zdnd11an1n64x5 FILLER_218_1328 ();
 b15zdnd11an1n64x5 FILLER_218_1392 ();
 b15zdnd11an1n64x5 FILLER_218_1456 ();
 b15zdnd11an1n64x5 FILLER_218_1520 ();
 b15zdnd11an1n64x5 FILLER_218_1584 ();
 b15zdnd11an1n64x5 FILLER_218_1648 ();
 b15zdnd11an1n64x5 FILLER_218_1712 ();
 b15zdnd11an1n64x5 FILLER_218_1776 ();
 b15zdnd11an1n64x5 FILLER_218_1840 ();
 b15zdnd11an1n64x5 FILLER_218_1904 ();
 b15zdnd11an1n64x5 FILLER_218_1968 ();
 b15zdnd11an1n64x5 FILLER_218_2032 ();
 b15zdnd11an1n32x5 FILLER_218_2096 ();
 b15zdnd11an1n16x5 FILLER_218_2128 ();
 b15zdnd11an1n08x5 FILLER_218_2144 ();
 b15zdnd00an1n02x5 FILLER_218_2152 ();
 b15zdnd11an1n64x5 FILLER_218_2162 ();
 b15zdnd11an1n16x5 FILLER_218_2226 ();
 b15zdnd00an1n02x5 FILLER_218_2242 ();
 b15zdnd00an1n01x5 FILLER_218_2244 ();
 b15zdnd11an1n08x5 FILLER_218_2249 ();
 b15zdnd11an1n04x5 FILLER_218_2257 ();
 b15zdnd11an1n08x5 FILLER_218_2265 ();
 b15zdnd00an1n02x5 FILLER_218_2273 ();
 b15zdnd00an1n01x5 FILLER_218_2275 ();
 b15zdnd11an1n08x5 FILLER_219_0 ();
 b15zdnd11an1n04x5 FILLER_219_8 ();
 b15zdnd00an1n02x5 FILLER_219_12 ();
 b15zdnd00an1n01x5 FILLER_219_14 ();
 b15zdnd11an1n64x5 FILLER_219_22 ();
 b15zdnd11an1n64x5 FILLER_219_86 ();
 b15zdnd11an1n64x5 FILLER_219_150 ();
 b15zdnd11an1n64x5 FILLER_219_214 ();
 b15zdnd11an1n64x5 FILLER_219_278 ();
 b15zdnd11an1n64x5 FILLER_219_342 ();
 b15zdnd11an1n64x5 FILLER_219_406 ();
 b15zdnd11an1n64x5 FILLER_219_470 ();
 b15zdnd11an1n64x5 FILLER_219_534 ();
 b15zdnd11an1n32x5 FILLER_219_598 ();
 b15zdnd11an1n16x5 FILLER_219_630 ();
 b15zdnd11an1n04x5 FILLER_219_646 ();
 b15zdnd00an1n01x5 FILLER_219_650 ();
 b15zdnd11an1n32x5 FILLER_219_667 ();
 b15zdnd11an1n16x5 FILLER_219_699 ();
 b15zdnd11an1n04x5 FILLER_219_757 ();
 b15zdnd11an1n16x5 FILLER_219_803 ();
 b15zdnd11an1n08x5 FILLER_219_819 ();
 b15zdnd11an1n04x5 FILLER_219_827 ();
 b15zdnd00an1n02x5 FILLER_219_831 ();
 b15zdnd11an1n04x5 FILLER_219_837 ();
 b15zdnd11an1n64x5 FILLER_219_849 ();
 b15zdnd11an1n64x5 FILLER_219_913 ();
 b15zdnd11an1n64x5 FILLER_219_977 ();
 b15zdnd11an1n64x5 FILLER_219_1041 ();
 b15zdnd11an1n64x5 FILLER_219_1105 ();
 b15zdnd11an1n64x5 FILLER_219_1169 ();
 b15zdnd11an1n32x5 FILLER_219_1233 ();
 b15zdnd00an1n02x5 FILLER_219_1265 ();
 b15zdnd00an1n01x5 FILLER_219_1267 ();
 b15zdnd11an1n64x5 FILLER_219_1310 ();
 b15zdnd11an1n64x5 FILLER_219_1374 ();
 b15zdnd11an1n64x5 FILLER_219_1438 ();
 b15zdnd11an1n64x5 FILLER_219_1502 ();
 b15zdnd11an1n64x5 FILLER_219_1566 ();
 b15zdnd11an1n64x5 FILLER_219_1630 ();
 b15zdnd11an1n64x5 FILLER_219_1694 ();
 b15zdnd11an1n64x5 FILLER_219_1758 ();
 b15zdnd11an1n64x5 FILLER_219_1822 ();
 b15zdnd11an1n64x5 FILLER_219_1886 ();
 b15zdnd11an1n64x5 FILLER_219_1950 ();
 b15zdnd11an1n64x5 FILLER_219_2014 ();
 b15zdnd11an1n32x5 FILLER_219_2078 ();
 b15zdnd11an1n08x5 FILLER_219_2110 ();
 b15zdnd00an1n02x5 FILLER_219_2118 ();
 b15zdnd00an1n01x5 FILLER_219_2120 ();
 b15zdnd11an1n64x5 FILLER_219_2133 ();
 b15zdnd11an1n32x5 FILLER_219_2197 ();
 b15zdnd11an1n08x5 FILLER_219_2229 ();
 b15zdnd00an1n02x5 FILLER_219_2237 ();
 b15zdnd00an1n01x5 FILLER_219_2239 ();
 b15zdnd00an1n02x5 FILLER_219_2282 ();
 b15zdnd00an1n02x5 FILLER_220_8 ();
 b15zdnd11an1n04x5 FILLER_220_18 ();
 b15zdnd11an1n64x5 FILLER_220_42 ();
 b15zdnd11an1n64x5 FILLER_220_106 ();
 b15zdnd11an1n64x5 FILLER_220_170 ();
 b15zdnd11an1n64x5 FILLER_220_234 ();
 b15zdnd11an1n64x5 FILLER_220_298 ();
 b15zdnd11an1n64x5 FILLER_220_362 ();
 b15zdnd11an1n64x5 FILLER_220_426 ();
 b15zdnd11an1n64x5 FILLER_220_490 ();
 b15zdnd11an1n64x5 FILLER_220_554 ();
 b15zdnd11an1n16x5 FILLER_220_618 ();
 b15zdnd11an1n08x5 FILLER_220_634 ();
 b15zdnd11an1n04x5 FILLER_220_642 ();
 b15zdnd11an1n04x5 FILLER_220_651 ();
 b15zdnd11an1n32x5 FILLER_220_667 ();
 b15zdnd11an1n16x5 FILLER_220_699 ();
 b15zdnd00an1n02x5 FILLER_220_715 ();
 b15zdnd00an1n01x5 FILLER_220_717 ();
 b15zdnd11an1n16x5 FILLER_220_726 ();
 b15zdnd11an1n08x5 FILLER_220_742 ();
 b15zdnd11an1n32x5 FILLER_220_792 ();
 b15zdnd11an1n16x5 FILLER_220_824 ();
 b15zdnd11an1n08x5 FILLER_220_840 ();
 b15zdnd11an1n04x5 FILLER_220_848 ();
 b15zdnd00an1n02x5 FILLER_220_852 ();
 b15zdnd11an1n64x5 FILLER_220_876 ();
 b15zdnd11an1n64x5 FILLER_220_940 ();
 b15zdnd11an1n64x5 FILLER_220_1004 ();
 b15zdnd11an1n64x5 FILLER_220_1068 ();
 b15zdnd11an1n64x5 FILLER_220_1132 ();
 b15zdnd11an1n64x5 FILLER_220_1196 ();
 b15zdnd11an1n64x5 FILLER_220_1260 ();
 b15zdnd11an1n64x5 FILLER_220_1324 ();
 b15zdnd11an1n64x5 FILLER_220_1388 ();
 b15zdnd11an1n64x5 FILLER_220_1452 ();
 b15zdnd11an1n64x5 FILLER_220_1516 ();
 b15zdnd11an1n64x5 FILLER_220_1580 ();
 b15zdnd11an1n64x5 FILLER_220_1644 ();
 b15zdnd11an1n64x5 FILLER_220_1708 ();
 b15zdnd11an1n64x5 FILLER_220_1772 ();
 b15zdnd11an1n64x5 FILLER_220_1836 ();
 b15zdnd11an1n64x5 FILLER_220_1900 ();
 b15zdnd11an1n64x5 FILLER_220_1964 ();
 b15zdnd11an1n64x5 FILLER_220_2028 ();
 b15zdnd11an1n04x5 FILLER_220_2134 ();
 b15zdnd11an1n04x5 FILLER_220_2150 ();
 b15zdnd11an1n64x5 FILLER_220_2162 ();
 b15zdnd11an1n32x5 FILLER_220_2226 ();
 b15zdnd11an1n16x5 FILLER_220_2258 ();
 b15zdnd00an1n02x5 FILLER_220_2274 ();
 b15zdnd11an1n64x5 FILLER_221_0 ();
 b15zdnd11an1n64x5 FILLER_221_64 ();
 b15zdnd11an1n64x5 FILLER_221_128 ();
 b15zdnd11an1n64x5 FILLER_221_192 ();
 b15zdnd11an1n64x5 FILLER_221_256 ();
 b15zdnd11an1n64x5 FILLER_221_320 ();
 b15zdnd11an1n64x5 FILLER_221_384 ();
 b15zdnd11an1n64x5 FILLER_221_448 ();
 b15zdnd11an1n64x5 FILLER_221_512 ();
 b15zdnd11an1n64x5 FILLER_221_576 ();
 b15zdnd11an1n32x5 FILLER_221_640 ();
 b15zdnd11an1n08x5 FILLER_221_672 ();
 b15zdnd11an1n04x5 FILLER_221_680 ();
 b15zdnd00an1n01x5 FILLER_221_684 ();
 b15zdnd11an1n64x5 FILLER_221_727 ();
 b15zdnd11an1n64x5 FILLER_221_791 ();
 b15zdnd11an1n64x5 FILLER_221_855 ();
 b15zdnd11an1n64x5 FILLER_221_919 ();
 b15zdnd11an1n64x5 FILLER_221_983 ();
 b15zdnd11an1n64x5 FILLER_221_1047 ();
 b15zdnd11an1n64x5 FILLER_221_1111 ();
 b15zdnd11an1n32x5 FILLER_221_1175 ();
 b15zdnd11an1n08x5 FILLER_221_1207 ();
 b15zdnd11an1n04x5 FILLER_221_1215 ();
 b15zdnd00an1n02x5 FILLER_221_1219 ();
 b15zdnd11an1n64x5 FILLER_221_1225 ();
 b15zdnd11an1n64x5 FILLER_221_1289 ();
 b15zdnd11an1n32x5 FILLER_221_1353 ();
 b15zdnd11an1n16x5 FILLER_221_1385 ();
 b15zdnd11an1n08x5 FILLER_221_1401 ();
 b15zdnd00an1n02x5 FILLER_221_1409 ();
 b15zdnd00an1n01x5 FILLER_221_1411 ();
 b15zdnd11an1n04x5 FILLER_221_1443 ();
 b15zdnd11an1n16x5 FILLER_221_1467 ();
 b15zdnd11an1n08x5 FILLER_221_1483 ();
 b15zdnd11an1n04x5 FILLER_221_1491 ();
 b15zdnd00an1n02x5 FILLER_221_1495 ();
 b15zdnd11an1n64x5 FILLER_221_1513 ();
 b15zdnd11an1n64x5 FILLER_221_1577 ();
 b15zdnd11an1n64x5 FILLER_221_1641 ();
 b15zdnd11an1n64x5 FILLER_221_1705 ();
 b15zdnd11an1n64x5 FILLER_221_1769 ();
 b15zdnd11an1n64x5 FILLER_221_1833 ();
 b15zdnd11an1n64x5 FILLER_221_1897 ();
 b15zdnd11an1n64x5 FILLER_221_1961 ();
 b15zdnd11an1n32x5 FILLER_221_2025 ();
 b15zdnd11an1n16x5 FILLER_221_2057 ();
 b15zdnd11an1n04x5 FILLER_221_2073 ();
 b15zdnd00an1n02x5 FILLER_221_2077 ();
 b15zdnd11an1n04x5 FILLER_221_2121 ();
 b15zdnd11an1n64x5 FILLER_221_2141 ();
 b15zdnd11an1n64x5 FILLER_221_2205 ();
 b15zdnd11an1n08x5 FILLER_221_2269 ();
 b15zdnd11an1n04x5 FILLER_221_2277 ();
 b15zdnd00an1n02x5 FILLER_221_2281 ();
 b15zdnd00an1n01x5 FILLER_221_2283 ();
 b15zdnd11an1n64x5 FILLER_222_8 ();
 b15zdnd11an1n64x5 FILLER_222_72 ();
 b15zdnd11an1n64x5 FILLER_222_136 ();
 b15zdnd11an1n64x5 FILLER_222_200 ();
 b15zdnd11an1n64x5 FILLER_222_264 ();
 b15zdnd11an1n64x5 FILLER_222_328 ();
 b15zdnd11an1n64x5 FILLER_222_392 ();
 b15zdnd11an1n64x5 FILLER_222_456 ();
 b15zdnd11an1n64x5 FILLER_222_520 ();
 b15zdnd11an1n64x5 FILLER_222_584 ();
 b15zdnd11an1n64x5 FILLER_222_648 ();
 b15zdnd11an1n04x5 FILLER_222_712 ();
 b15zdnd00an1n02x5 FILLER_222_716 ();
 b15zdnd11an1n64x5 FILLER_222_726 ();
 b15zdnd11an1n64x5 FILLER_222_790 ();
 b15zdnd11an1n64x5 FILLER_222_854 ();
 b15zdnd11an1n64x5 FILLER_222_918 ();
 b15zdnd11an1n64x5 FILLER_222_982 ();
 b15zdnd11an1n64x5 FILLER_222_1046 ();
 b15zdnd11an1n64x5 FILLER_222_1110 ();
 b15zdnd11an1n04x5 FILLER_222_1174 ();
 b15zdnd00an1n01x5 FILLER_222_1178 ();
 b15zdnd11an1n64x5 FILLER_222_1221 ();
 b15zdnd11an1n64x5 FILLER_222_1285 ();
 b15zdnd11an1n32x5 FILLER_222_1349 ();
 b15zdnd11an1n08x5 FILLER_222_1381 ();
 b15zdnd11an1n04x5 FILLER_222_1389 ();
 b15zdnd00an1n01x5 FILLER_222_1393 ();
 b15zdnd11an1n16x5 FILLER_222_1425 ();
 b15zdnd11an1n04x5 FILLER_222_1441 ();
 b15zdnd00an1n02x5 FILLER_222_1445 ();
 b15zdnd11an1n32x5 FILLER_222_1467 ();
 b15zdnd11an1n08x5 FILLER_222_1499 ();
 b15zdnd11an1n04x5 FILLER_222_1507 ();
 b15zdnd00an1n02x5 FILLER_222_1511 ();
 b15zdnd11an1n16x5 FILLER_222_1525 ();
 b15zdnd11an1n64x5 FILLER_222_1557 ();
 b15zdnd11an1n64x5 FILLER_222_1621 ();
 b15zdnd11an1n64x5 FILLER_222_1685 ();
 b15zdnd11an1n64x5 FILLER_222_1749 ();
 b15zdnd11an1n64x5 FILLER_222_1813 ();
 b15zdnd11an1n32x5 FILLER_222_1877 ();
 b15zdnd11an1n08x5 FILLER_222_1909 ();
 b15zdnd00an1n01x5 FILLER_222_1917 ();
 b15zdnd11an1n04x5 FILLER_222_1926 ();
 b15zdnd11an1n64x5 FILLER_222_1940 ();
 b15zdnd11an1n64x5 FILLER_222_2004 ();
 b15zdnd11an1n16x5 FILLER_222_2068 ();
 b15zdnd11an1n04x5 FILLER_222_2084 ();
 b15zdnd00an1n01x5 FILLER_222_2088 ();
 b15zdnd11an1n04x5 FILLER_222_2101 ();
 b15zdnd11an1n04x5 FILLER_222_2115 ();
 b15zdnd00an1n02x5 FILLER_222_2119 ();
 b15zdnd11an1n16x5 FILLER_222_2133 ();
 b15zdnd11an1n04x5 FILLER_222_2149 ();
 b15zdnd00an1n01x5 FILLER_222_2153 ();
 b15zdnd11an1n64x5 FILLER_222_2162 ();
 b15zdnd11an1n32x5 FILLER_222_2226 ();
 b15zdnd11an1n16x5 FILLER_222_2258 ();
 b15zdnd00an1n02x5 FILLER_222_2274 ();
 b15zdnd11an1n64x5 FILLER_223_0 ();
 b15zdnd11an1n64x5 FILLER_223_64 ();
 b15zdnd11an1n64x5 FILLER_223_128 ();
 b15zdnd11an1n64x5 FILLER_223_192 ();
 b15zdnd11an1n64x5 FILLER_223_256 ();
 b15zdnd11an1n64x5 FILLER_223_320 ();
 b15zdnd11an1n64x5 FILLER_223_384 ();
 b15zdnd11an1n64x5 FILLER_223_448 ();
 b15zdnd11an1n64x5 FILLER_223_512 ();
 b15zdnd11an1n64x5 FILLER_223_576 ();
 b15zdnd11an1n64x5 FILLER_223_640 ();
 b15zdnd11an1n64x5 FILLER_223_704 ();
 b15zdnd11an1n16x5 FILLER_223_768 ();
 b15zdnd11an1n64x5 FILLER_223_800 ();
 b15zdnd11an1n64x5 FILLER_223_864 ();
 b15zdnd11an1n64x5 FILLER_223_928 ();
 b15zdnd11an1n64x5 FILLER_223_992 ();
 b15zdnd11an1n64x5 FILLER_223_1056 ();
 b15zdnd11an1n64x5 FILLER_223_1120 ();
 b15zdnd11an1n64x5 FILLER_223_1184 ();
 b15zdnd11an1n64x5 FILLER_223_1248 ();
 b15zdnd11an1n64x5 FILLER_223_1312 ();
 b15zdnd11an1n64x5 FILLER_223_1376 ();
 b15zdnd11an1n64x5 FILLER_223_1440 ();
 b15zdnd11an1n08x5 FILLER_223_1504 ();
 b15zdnd11an1n04x5 FILLER_223_1512 ();
 b15zdnd11an1n64x5 FILLER_223_1536 ();
 b15zdnd11an1n32x5 FILLER_223_1600 ();
 b15zdnd11an1n16x5 FILLER_223_1632 ();
 b15zdnd11an1n08x5 FILLER_223_1648 ();
 b15zdnd00an1n02x5 FILLER_223_1656 ();
 b15zdnd00an1n01x5 FILLER_223_1658 ();
 b15zdnd11an1n64x5 FILLER_223_1701 ();
 b15zdnd11an1n64x5 FILLER_223_1765 ();
 b15zdnd11an1n32x5 FILLER_223_1829 ();
 b15zdnd11an1n16x5 FILLER_223_1861 ();
 b15zdnd11an1n08x5 FILLER_223_1877 ();
 b15zdnd00an1n02x5 FILLER_223_1885 ();
 b15zdnd11an1n04x5 FILLER_223_1903 ();
 b15zdnd11an1n08x5 FILLER_223_1918 ();
 b15zdnd00an1n01x5 FILLER_223_1926 ();
 b15zdnd11an1n64x5 FILLER_223_1939 ();
 b15zdnd11an1n64x5 FILLER_223_2003 ();
 b15zdnd11an1n32x5 FILLER_223_2067 ();
 b15zdnd11an1n08x5 FILLER_223_2099 ();
 b15zdnd11an1n04x5 FILLER_223_2117 ();
 b15zdnd11an1n64x5 FILLER_223_2131 ();
 b15zdnd11an1n64x5 FILLER_223_2195 ();
 b15zdnd11an1n16x5 FILLER_223_2259 ();
 b15zdnd11an1n08x5 FILLER_223_2275 ();
 b15zdnd00an1n01x5 FILLER_223_2283 ();
 b15zdnd11an1n64x5 FILLER_224_8 ();
 b15zdnd11an1n64x5 FILLER_224_72 ();
 b15zdnd11an1n64x5 FILLER_224_136 ();
 b15zdnd11an1n64x5 FILLER_224_200 ();
 b15zdnd11an1n64x5 FILLER_224_264 ();
 b15zdnd11an1n64x5 FILLER_224_328 ();
 b15zdnd11an1n64x5 FILLER_224_392 ();
 b15zdnd11an1n64x5 FILLER_224_456 ();
 b15zdnd11an1n64x5 FILLER_224_520 ();
 b15zdnd11an1n64x5 FILLER_224_584 ();
 b15zdnd11an1n64x5 FILLER_224_648 ();
 b15zdnd11an1n04x5 FILLER_224_712 ();
 b15zdnd00an1n02x5 FILLER_224_716 ();
 b15zdnd11an1n64x5 FILLER_224_726 ();
 b15zdnd11an1n64x5 FILLER_224_790 ();
 b15zdnd11an1n64x5 FILLER_224_854 ();
 b15zdnd11an1n64x5 FILLER_224_918 ();
 b15zdnd11an1n64x5 FILLER_224_982 ();
 b15zdnd11an1n64x5 FILLER_224_1046 ();
 b15zdnd11an1n64x5 FILLER_224_1110 ();
 b15zdnd11an1n64x5 FILLER_224_1174 ();
 b15zdnd11an1n64x5 FILLER_224_1238 ();
 b15zdnd11an1n64x5 FILLER_224_1302 ();
 b15zdnd11an1n64x5 FILLER_224_1366 ();
 b15zdnd11an1n64x5 FILLER_224_1430 ();
 b15zdnd11an1n16x5 FILLER_224_1494 ();
 b15zdnd00an1n02x5 FILLER_224_1510 ();
 b15zdnd11an1n64x5 FILLER_224_1523 ();
 b15zdnd11an1n64x5 FILLER_224_1587 ();
 b15zdnd11an1n04x5 FILLER_224_1651 ();
 b15zdnd00an1n02x5 FILLER_224_1655 ();
 b15zdnd00an1n01x5 FILLER_224_1657 ();
 b15zdnd11an1n16x5 FILLER_224_1700 ();
 b15zdnd11an1n16x5 FILLER_224_1726 ();
 b15zdnd11an1n08x5 FILLER_224_1742 ();
 b15zdnd00an1n02x5 FILLER_224_1750 ();
 b15zdnd00an1n01x5 FILLER_224_1752 ();
 b15zdnd11an1n04x5 FILLER_224_1765 ();
 b15zdnd00an1n02x5 FILLER_224_1769 ();
 b15zdnd00an1n01x5 FILLER_224_1771 ();
 b15zdnd11an1n64x5 FILLER_224_1795 ();
 b15zdnd11an1n16x5 FILLER_224_1859 ();
 b15zdnd11an1n08x5 FILLER_224_1875 ();
 b15zdnd00an1n02x5 FILLER_224_1883 ();
 b15zdnd11an1n32x5 FILLER_224_1895 ();
 b15zdnd11an1n04x5 FILLER_224_1927 ();
 b15zdnd00an1n02x5 FILLER_224_1931 ();
 b15zdnd11an1n64x5 FILLER_224_1949 ();
 b15zdnd11an1n64x5 FILLER_224_2013 ();
 b15zdnd11an1n64x5 FILLER_224_2077 ();
 b15zdnd11an1n08x5 FILLER_224_2141 ();
 b15zdnd11an1n04x5 FILLER_224_2149 ();
 b15zdnd00an1n01x5 FILLER_224_2153 ();
 b15zdnd11an1n64x5 FILLER_224_2162 ();
 b15zdnd11an1n32x5 FILLER_224_2226 ();
 b15zdnd11an1n16x5 FILLER_224_2258 ();
 b15zdnd00an1n02x5 FILLER_224_2274 ();
 b15zdnd11an1n64x5 FILLER_225_0 ();
 b15zdnd11an1n64x5 FILLER_225_64 ();
 b15zdnd11an1n64x5 FILLER_225_128 ();
 b15zdnd11an1n64x5 FILLER_225_192 ();
 b15zdnd11an1n64x5 FILLER_225_256 ();
 b15zdnd11an1n64x5 FILLER_225_320 ();
 b15zdnd11an1n64x5 FILLER_225_384 ();
 b15zdnd11an1n64x5 FILLER_225_448 ();
 b15zdnd11an1n64x5 FILLER_225_512 ();
 b15zdnd11an1n64x5 FILLER_225_576 ();
 b15zdnd11an1n32x5 FILLER_225_640 ();
 b15zdnd00an1n02x5 FILLER_225_672 ();
 b15zdnd00an1n01x5 FILLER_225_674 ();
 b15zdnd11an1n64x5 FILLER_225_678 ();
 b15zdnd11an1n64x5 FILLER_225_742 ();
 b15zdnd11an1n64x5 FILLER_225_806 ();
 b15zdnd11an1n64x5 FILLER_225_870 ();
 b15zdnd11an1n64x5 FILLER_225_934 ();
 b15zdnd11an1n64x5 FILLER_225_998 ();
 b15zdnd11an1n64x5 FILLER_225_1062 ();
 b15zdnd11an1n64x5 FILLER_225_1126 ();
 b15zdnd11an1n04x5 FILLER_225_1190 ();
 b15zdnd11an1n64x5 FILLER_225_1198 ();
 b15zdnd11an1n64x5 FILLER_225_1262 ();
 b15zdnd11an1n64x5 FILLER_225_1326 ();
 b15zdnd11an1n64x5 FILLER_225_1390 ();
 b15zdnd11an1n64x5 FILLER_225_1454 ();
 b15zdnd11an1n64x5 FILLER_225_1518 ();
 b15zdnd11an1n16x5 FILLER_225_1582 ();
 b15zdnd00an1n02x5 FILLER_225_1598 ();
 b15zdnd00an1n01x5 FILLER_225_1600 ();
 b15zdnd11an1n04x5 FILLER_225_1617 ();
 b15zdnd11an1n08x5 FILLER_225_1637 ();
 b15zdnd11an1n04x5 FILLER_225_1645 ();
 b15zdnd00an1n02x5 FILLER_225_1649 ();
 b15zdnd00an1n01x5 FILLER_225_1651 ();
 b15zdnd11an1n64x5 FILLER_225_1694 ();
 b15zdnd11an1n64x5 FILLER_225_1758 ();
 b15zdnd11an1n16x5 FILLER_225_1822 ();
 b15zdnd11an1n04x5 FILLER_225_1838 ();
 b15zdnd00an1n02x5 FILLER_225_1842 ();
 b15zdnd00an1n01x5 FILLER_225_1844 ();
 b15zdnd11an1n64x5 FILLER_225_1861 ();
 b15zdnd11an1n64x5 FILLER_225_1925 ();
 b15zdnd11an1n64x5 FILLER_225_1989 ();
 b15zdnd11an1n16x5 FILLER_225_2053 ();
 b15zdnd11an1n04x5 FILLER_225_2069 ();
 b15zdnd00an1n02x5 FILLER_225_2073 ();
 b15zdnd11an1n64x5 FILLER_225_2117 ();
 b15zdnd11an1n64x5 FILLER_225_2181 ();
 b15zdnd11an1n04x5 FILLER_225_2245 ();
 b15zdnd00an1n02x5 FILLER_225_2249 ();
 b15zdnd00an1n01x5 FILLER_225_2251 ();
 b15zdnd11an1n16x5 FILLER_225_2256 ();
 b15zdnd11an1n08x5 FILLER_225_2272 ();
 b15zdnd11an1n04x5 FILLER_225_2280 ();
 b15zdnd11an1n64x5 FILLER_226_8 ();
 b15zdnd11an1n64x5 FILLER_226_72 ();
 b15zdnd11an1n64x5 FILLER_226_136 ();
 b15zdnd11an1n64x5 FILLER_226_200 ();
 b15zdnd11an1n64x5 FILLER_226_264 ();
 b15zdnd11an1n64x5 FILLER_226_328 ();
 b15zdnd11an1n64x5 FILLER_226_392 ();
 b15zdnd11an1n64x5 FILLER_226_456 ();
 b15zdnd11an1n64x5 FILLER_226_520 ();
 b15zdnd11an1n64x5 FILLER_226_584 ();
 b15zdnd11an1n64x5 FILLER_226_648 ();
 b15zdnd11an1n04x5 FILLER_226_712 ();
 b15zdnd00an1n02x5 FILLER_226_716 ();
 b15zdnd11an1n64x5 FILLER_226_726 ();
 b15zdnd11an1n64x5 FILLER_226_790 ();
 b15zdnd11an1n64x5 FILLER_226_854 ();
 b15zdnd11an1n04x5 FILLER_226_918 ();
 b15zdnd00an1n02x5 FILLER_226_922 ();
 b15zdnd11an1n64x5 FILLER_226_966 ();
 b15zdnd11an1n64x5 FILLER_226_1030 ();
 b15zdnd11an1n64x5 FILLER_226_1094 ();
 b15zdnd11an1n64x5 FILLER_226_1158 ();
 b15zdnd11an1n64x5 FILLER_226_1222 ();
 b15zdnd11an1n64x5 FILLER_226_1286 ();
 b15zdnd11an1n64x5 FILLER_226_1350 ();
 b15zdnd11an1n64x5 FILLER_226_1414 ();
 b15zdnd11an1n64x5 FILLER_226_1478 ();
 b15zdnd11an1n64x5 FILLER_226_1542 ();
 b15zdnd11an1n16x5 FILLER_226_1606 ();
 b15zdnd11an1n08x5 FILLER_226_1622 ();
 b15zdnd00an1n01x5 FILLER_226_1630 ();
 b15zdnd11an1n16x5 FILLER_226_1673 ();
 b15zdnd11an1n04x5 FILLER_226_1689 ();
 b15zdnd00an1n02x5 FILLER_226_1693 ();
 b15zdnd11an1n64x5 FILLER_226_1718 ();
 b15zdnd11an1n64x5 FILLER_226_1782 ();
 b15zdnd11an1n08x5 FILLER_226_1846 ();
 b15zdnd11an1n04x5 FILLER_226_1854 ();
 b15zdnd00an1n01x5 FILLER_226_1858 ();
 b15zdnd11an1n64x5 FILLER_226_1867 ();
 b15zdnd11an1n64x5 FILLER_226_1931 ();
 b15zdnd11an1n64x5 FILLER_226_1995 ();
 b15zdnd11an1n32x5 FILLER_226_2101 ();
 b15zdnd11an1n16x5 FILLER_226_2133 ();
 b15zdnd11an1n04x5 FILLER_226_2149 ();
 b15zdnd00an1n01x5 FILLER_226_2153 ();
 b15zdnd11an1n64x5 FILLER_226_2162 ();
 b15zdnd11an1n04x5 FILLER_226_2226 ();
 b15zdnd00an1n02x5 FILLER_226_2230 ();
 b15zdnd00an1n02x5 FILLER_226_2274 ();
 b15zdnd11an1n64x5 FILLER_227_0 ();
 b15zdnd11an1n64x5 FILLER_227_64 ();
 b15zdnd11an1n64x5 FILLER_227_128 ();
 b15zdnd11an1n64x5 FILLER_227_192 ();
 b15zdnd11an1n64x5 FILLER_227_256 ();
 b15zdnd11an1n64x5 FILLER_227_320 ();
 b15zdnd11an1n64x5 FILLER_227_384 ();
 b15zdnd11an1n64x5 FILLER_227_448 ();
 b15zdnd11an1n64x5 FILLER_227_512 ();
 b15zdnd11an1n64x5 FILLER_227_576 ();
 b15zdnd11an1n64x5 FILLER_227_640 ();
 b15zdnd11an1n64x5 FILLER_227_704 ();
 b15zdnd11an1n64x5 FILLER_227_768 ();
 b15zdnd11an1n16x5 FILLER_227_832 ();
 b15zdnd11an1n04x5 FILLER_227_848 ();
 b15zdnd00an1n02x5 FILLER_227_852 ();
 b15zdnd00an1n01x5 FILLER_227_854 ();
 b15zdnd11an1n64x5 FILLER_227_871 ();
 b15zdnd11an1n64x5 FILLER_227_935 ();
 b15zdnd11an1n64x5 FILLER_227_999 ();
 b15zdnd11an1n64x5 FILLER_227_1063 ();
 b15zdnd11an1n64x5 FILLER_227_1127 ();
 b15zdnd11an1n64x5 FILLER_227_1191 ();
 b15zdnd11an1n64x5 FILLER_227_1255 ();
 b15zdnd11an1n64x5 FILLER_227_1319 ();
 b15zdnd11an1n64x5 FILLER_227_1383 ();
 b15zdnd11an1n64x5 FILLER_227_1447 ();
 b15zdnd11an1n64x5 FILLER_227_1511 ();
 b15zdnd11an1n64x5 FILLER_227_1575 ();
 b15zdnd11an1n64x5 FILLER_227_1639 ();
 b15zdnd11an1n64x5 FILLER_227_1703 ();
 b15zdnd11an1n64x5 FILLER_227_1767 ();
 b15zdnd11an1n16x5 FILLER_227_1831 ();
 b15zdnd11an1n08x5 FILLER_227_1847 ();
 b15zdnd11an1n04x5 FILLER_227_1855 ();
 b15zdnd00an1n02x5 FILLER_227_1859 ();
 b15zdnd11an1n16x5 FILLER_227_1869 ();
 b15zdnd11an1n64x5 FILLER_227_1893 ();
 b15zdnd11an1n64x5 FILLER_227_1957 ();
 b15zdnd11an1n32x5 FILLER_227_2021 ();
 b15zdnd11an1n08x5 FILLER_227_2053 ();
 b15zdnd11an1n04x5 FILLER_227_2061 ();
 b15zdnd00an1n02x5 FILLER_227_2065 ();
 b15zdnd00an1n01x5 FILLER_227_2067 ();
 b15zdnd11an1n64x5 FILLER_227_2110 ();
 b15zdnd11an1n64x5 FILLER_227_2174 ();
 b15zdnd11an1n16x5 FILLER_227_2238 ();
 b15zdnd00an1n02x5 FILLER_227_2254 ();
 b15zdnd00an1n01x5 FILLER_227_2256 ();
 b15zdnd11an1n04x5 FILLER_227_2261 ();
 b15zdnd00an1n02x5 FILLER_227_2265 ();
 b15zdnd00an1n01x5 FILLER_227_2267 ();
 b15zdnd11an1n04x5 FILLER_227_2272 ();
 b15zdnd11an1n04x5 FILLER_227_2280 ();
 b15zdnd11an1n64x5 FILLER_228_8 ();
 b15zdnd11an1n64x5 FILLER_228_72 ();
 b15zdnd11an1n64x5 FILLER_228_136 ();
 b15zdnd11an1n64x5 FILLER_228_200 ();
 b15zdnd11an1n64x5 FILLER_228_264 ();
 b15zdnd11an1n64x5 FILLER_228_328 ();
 b15zdnd11an1n64x5 FILLER_228_392 ();
 b15zdnd11an1n64x5 FILLER_228_456 ();
 b15zdnd11an1n64x5 FILLER_228_520 ();
 b15zdnd11an1n64x5 FILLER_228_584 ();
 b15zdnd11an1n64x5 FILLER_228_648 ();
 b15zdnd11an1n04x5 FILLER_228_712 ();
 b15zdnd00an1n02x5 FILLER_228_716 ();
 b15zdnd11an1n64x5 FILLER_228_726 ();
 b15zdnd11an1n64x5 FILLER_228_790 ();
 b15zdnd11an1n64x5 FILLER_228_854 ();
 b15zdnd11an1n64x5 FILLER_228_918 ();
 b15zdnd11an1n64x5 FILLER_228_982 ();
 b15zdnd00an1n02x5 FILLER_228_1046 ();
 b15zdnd00an1n01x5 FILLER_228_1048 ();
 b15zdnd11an1n64x5 FILLER_228_1091 ();
 b15zdnd11an1n64x5 FILLER_228_1155 ();
 b15zdnd11an1n64x5 FILLER_228_1219 ();
 b15zdnd11an1n64x5 FILLER_228_1283 ();
 b15zdnd11an1n64x5 FILLER_228_1347 ();
 b15zdnd11an1n64x5 FILLER_228_1411 ();
 b15zdnd11an1n64x5 FILLER_228_1475 ();
 b15zdnd11an1n64x5 FILLER_228_1539 ();
 b15zdnd11an1n64x5 FILLER_228_1603 ();
 b15zdnd11an1n64x5 FILLER_228_1667 ();
 b15zdnd11an1n64x5 FILLER_228_1731 ();
 b15zdnd11an1n64x5 FILLER_228_1795 ();
 b15zdnd11an1n64x5 FILLER_228_1859 ();
 b15zdnd11an1n64x5 FILLER_228_1923 ();
 b15zdnd11an1n64x5 FILLER_228_1987 ();
 b15zdnd00an1n02x5 FILLER_228_2051 ();
 b15zdnd00an1n01x5 FILLER_228_2053 ();
 b15zdnd11an1n32x5 FILLER_228_2096 ();
 b15zdnd11an1n16x5 FILLER_228_2128 ();
 b15zdnd11an1n08x5 FILLER_228_2144 ();
 b15zdnd00an1n02x5 FILLER_228_2152 ();
 b15zdnd11an1n64x5 FILLER_228_2162 ();
 b15zdnd11an1n04x5 FILLER_228_2226 ();
 b15zdnd00an1n02x5 FILLER_228_2230 ();
 b15zdnd00an1n02x5 FILLER_228_2274 ();
 b15zdnd11an1n64x5 FILLER_229_0 ();
 b15zdnd11an1n64x5 FILLER_229_64 ();
 b15zdnd11an1n64x5 FILLER_229_128 ();
 b15zdnd11an1n64x5 FILLER_229_192 ();
 b15zdnd11an1n64x5 FILLER_229_256 ();
 b15zdnd11an1n64x5 FILLER_229_320 ();
 b15zdnd11an1n64x5 FILLER_229_384 ();
 b15zdnd11an1n64x5 FILLER_229_448 ();
 b15zdnd11an1n64x5 FILLER_229_512 ();
 b15zdnd11an1n64x5 FILLER_229_576 ();
 b15zdnd11an1n64x5 FILLER_229_640 ();
 b15zdnd11an1n64x5 FILLER_229_704 ();
 b15zdnd11an1n64x5 FILLER_229_768 ();
 b15zdnd11an1n16x5 FILLER_229_832 ();
 b15zdnd11an1n04x5 FILLER_229_848 ();
 b15zdnd00an1n01x5 FILLER_229_852 ();
 b15zdnd11an1n64x5 FILLER_229_895 ();
 b15zdnd11an1n64x5 FILLER_229_959 ();
 b15zdnd11an1n64x5 FILLER_229_1023 ();
 b15zdnd11an1n32x5 FILLER_229_1087 ();
 b15zdnd11an1n16x5 FILLER_229_1119 ();
 b15zdnd11an1n08x5 FILLER_229_1135 ();
 b15zdnd00an1n02x5 FILLER_229_1143 ();
 b15zdnd00an1n01x5 FILLER_229_1145 ();
 b15zdnd11an1n32x5 FILLER_229_1162 ();
 b15zdnd11an1n16x5 FILLER_229_1194 ();
 b15zdnd11an1n08x5 FILLER_229_1210 ();
 b15zdnd11an1n04x5 FILLER_229_1218 ();
 b15zdnd11an1n64x5 FILLER_229_1253 ();
 b15zdnd11an1n64x5 FILLER_229_1317 ();
 b15zdnd11an1n64x5 FILLER_229_1381 ();
 b15zdnd11an1n64x5 FILLER_229_1445 ();
 b15zdnd11an1n64x5 FILLER_229_1509 ();
 b15zdnd11an1n64x5 FILLER_229_1573 ();
 b15zdnd11an1n64x5 FILLER_229_1637 ();
 b15zdnd00an1n01x5 FILLER_229_1701 ();
 b15zdnd11an1n16x5 FILLER_229_1718 ();
 b15zdnd11an1n04x5 FILLER_229_1734 ();
 b15zdnd00an1n01x5 FILLER_229_1738 ();
 b15zdnd11an1n64x5 FILLER_229_1759 ();
 b15zdnd00an1n02x5 FILLER_229_1823 ();
 b15zdnd11an1n64x5 FILLER_229_1833 ();
 b15zdnd11an1n08x5 FILLER_229_1897 ();
 b15zdnd11an1n04x5 FILLER_229_1905 ();
 b15zdnd00an1n02x5 FILLER_229_1909 ();
 b15zdnd00an1n01x5 FILLER_229_1911 ();
 b15zdnd11an1n64x5 FILLER_229_1928 ();
 b15zdnd11an1n64x5 FILLER_229_1992 ();
 b15zdnd11an1n64x5 FILLER_229_2056 ();
 b15zdnd11an1n64x5 FILLER_229_2120 ();
 b15zdnd11an1n64x5 FILLER_229_2184 ();
 b15zdnd11an1n32x5 FILLER_229_2248 ();
 b15zdnd11an1n04x5 FILLER_229_2280 ();
 b15zdnd11an1n64x5 FILLER_230_8 ();
 b15zdnd11an1n64x5 FILLER_230_72 ();
 b15zdnd11an1n64x5 FILLER_230_136 ();
 b15zdnd11an1n64x5 FILLER_230_200 ();
 b15zdnd11an1n64x5 FILLER_230_264 ();
 b15zdnd11an1n64x5 FILLER_230_328 ();
 b15zdnd11an1n64x5 FILLER_230_392 ();
 b15zdnd11an1n64x5 FILLER_230_456 ();
 b15zdnd11an1n64x5 FILLER_230_520 ();
 b15zdnd11an1n64x5 FILLER_230_584 ();
 b15zdnd11an1n64x5 FILLER_230_648 ();
 b15zdnd11an1n04x5 FILLER_230_712 ();
 b15zdnd00an1n02x5 FILLER_230_716 ();
 b15zdnd11an1n64x5 FILLER_230_726 ();
 b15zdnd11an1n64x5 FILLER_230_790 ();
 b15zdnd11an1n16x5 FILLER_230_854 ();
 b15zdnd11an1n04x5 FILLER_230_870 ();
 b15zdnd11an1n64x5 FILLER_230_886 ();
 b15zdnd11an1n64x5 FILLER_230_950 ();
 b15zdnd11an1n64x5 FILLER_230_1014 ();
 b15zdnd11an1n64x5 FILLER_230_1078 ();
 b15zdnd11an1n64x5 FILLER_230_1142 ();
 b15zdnd11an1n64x5 FILLER_230_1206 ();
 b15zdnd11an1n64x5 FILLER_230_1270 ();
 b15zdnd11an1n08x5 FILLER_230_1334 ();
 b15zdnd11an1n04x5 FILLER_230_1342 ();
 b15zdnd00an1n02x5 FILLER_230_1346 ();
 b15zdnd00an1n01x5 FILLER_230_1348 ();
 b15zdnd11an1n64x5 FILLER_230_1365 ();
 b15zdnd11an1n64x5 FILLER_230_1429 ();
 b15zdnd11an1n64x5 FILLER_230_1493 ();
 b15zdnd11an1n64x5 FILLER_230_1557 ();
 b15zdnd11an1n64x5 FILLER_230_1621 ();
 b15zdnd11an1n04x5 FILLER_230_1685 ();
 b15zdnd00an1n02x5 FILLER_230_1689 ();
 b15zdnd00an1n01x5 FILLER_230_1691 ();
 b15zdnd11an1n64x5 FILLER_230_1704 ();
 b15zdnd11an1n64x5 FILLER_230_1768 ();
 b15zdnd11an1n64x5 FILLER_230_1832 ();
 b15zdnd11an1n32x5 FILLER_230_1896 ();
 b15zdnd11an1n16x5 FILLER_230_1928 ();
 b15zdnd00an1n02x5 FILLER_230_1944 ();
 b15zdnd00an1n01x5 FILLER_230_1946 ();
 b15zdnd11an1n64x5 FILLER_230_1959 ();
 b15zdnd11an1n64x5 FILLER_230_2023 ();
 b15zdnd11an1n64x5 FILLER_230_2087 ();
 b15zdnd00an1n02x5 FILLER_230_2151 ();
 b15zdnd00an1n01x5 FILLER_230_2153 ();
 b15zdnd11an1n64x5 FILLER_230_2162 ();
 b15zdnd11an1n32x5 FILLER_230_2226 ();
 b15zdnd11an1n16x5 FILLER_230_2258 ();
 b15zdnd00an1n02x5 FILLER_230_2274 ();
 b15zdnd11an1n64x5 FILLER_231_0 ();
 b15zdnd11an1n64x5 FILLER_231_64 ();
 b15zdnd11an1n64x5 FILLER_231_128 ();
 b15zdnd11an1n64x5 FILLER_231_192 ();
 b15zdnd11an1n64x5 FILLER_231_256 ();
 b15zdnd11an1n64x5 FILLER_231_320 ();
 b15zdnd11an1n64x5 FILLER_231_384 ();
 b15zdnd11an1n64x5 FILLER_231_448 ();
 b15zdnd11an1n64x5 FILLER_231_512 ();
 b15zdnd11an1n64x5 FILLER_231_576 ();
 b15zdnd11an1n64x5 FILLER_231_640 ();
 b15zdnd11an1n64x5 FILLER_231_704 ();
 b15zdnd11an1n64x5 FILLER_231_768 ();
 b15zdnd11an1n16x5 FILLER_231_832 ();
 b15zdnd11an1n08x5 FILLER_231_848 ();
 b15zdnd11an1n64x5 FILLER_231_898 ();
 b15zdnd11an1n64x5 FILLER_231_962 ();
 b15zdnd11an1n64x5 FILLER_231_1026 ();
 b15zdnd11an1n64x5 FILLER_231_1090 ();
 b15zdnd11an1n04x5 FILLER_231_1154 ();
 b15zdnd00an1n02x5 FILLER_231_1158 ();
 b15zdnd11an1n64x5 FILLER_231_1173 ();
 b15zdnd11an1n16x5 FILLER_231_1237 ();
 b15zdnd11an1n04x5 FILLER_231_1253 ();
 b15zdnd00an1n02x5 FILLER_231_1257 ();
 b15zdnd11an1n64x5 FILLER_231_1275 ();
 b15zdnd11an1n64x5 FILLER_231_1339 ();
 b15zdnd11an1n64x5 FILLER_231_1403 ();
 b15zdnd11an1n64x5 FILLER_231_1467 ();
 b15zdnd11an1n64x5 FILLER_231_1531 ();
 b15zdnd11an1n64x5 FILLER_231_1595 ();
 b15zdnd11an1n32x5 FILLER_231_1659 ();
 b15zdnd11an1n16x5 FILLER_231_1691 ();
 b15zdnd00an1n02x5 FILLER_231_1707 ();
 b15zdnd11an1n64x5 FILLER_231_1729 ();
 b15zdnd11an1n64x5 FILLER_231_1793 ();
 b15zdnd11an1n64x5 FILLER_231_1857 ();
 b15zdnd11an1n64x5 FILLER_231_1921 ();
 b15zdnd11an1n64x5 FILLER_231_1985 ();
 b15zdnd11an1n64x5 FILLER_231_2049 ();
 b15zdnd11an1n64x5 FILLER_231_2113 ();
 b15zdnd11an1n64x5 FILLER_231_2177 ();
 b15zdnd11an1n32x5 FILLER_231_2241 ();
 b15zdnd11an1n08x5 FILLER_231_2273 ();
 b15zdnd00an1n02x5 FILLER_231_2281 ();
 b15zdnd00an1n01x5 FILLER_231_2283 ();
 b15zdnd11an1n64x5 FILLER_232_8 ();
 b15zdnd11an1n64x5 FILLER_232_72 ();
 b15zdnd11an1n64x5 FILLER_232_136 ();
 b15zdnd11an1n64x5 FILLER_232_200 ();
 b15zdnd11an1n64x5 FILLER_232_264 ();
 b15zdnd11an1n64x5 FILLER_232_328 ();
 b15zdnd11an1n64x5 FILLER_232_392 ();
 b15zdnd11an1n64x5 FILLER_232_456 ();
 b15zdnd11an1n64x5 FILLER_232_520 ();
 b15zdnd11an1n64x5 FILLER_232_584 ();
 b15zdnd11an1n64x5 FILLER_232_648 ();
 b15zdnd11an1n04x5 FILLER_232_712 ();
 b15zdnd00an1n02x5 FILLER_232_716 ();
 b15zdnd11an1n64x5 FILLER_232_726 ();
 b15zdnd11an1n64x5 FILLER_232_790 ();
 b15zdnd11an1n64x5 FILLER_232_854 ();
 b15zdnd11an1n64x5 FILLER_232_918 ();
 b15zdnd11an1n64x5 FILLER_232_982 ();
 b15zdnd11an1n64x5 FILLER_232_1046 ();
 b15zdnd11an1n32x5 FILLER_232_1110 ();
 b15zdnd11an1n16x5 FILLER_232_1142 ();
 b15zdnd11an1n08x5 FILLER_232_1158 ();
 b15zdnd11an1n64x5 FILLER_232_1179 ();
 b15zdnd11an1n08x5 FILLER_232_1243 ();
 b15zdnd11an1n04x5 FILLER_232_1251 ();
 b15zdnd11an1n32x5 FILLER_232_1275 ();
 b15zdnd11an1n04x5 FILLER_232_1307 ();
 b15zdnd11an1n64x5 FILLER_232_1353 ();
 b15zdnd11an1n64x5 FILLER_232_1417 ();
 b15zdnd11an1n64x5 FILLER_232_1481 ();
 b15zdnd11an1n64x5 FILLER_232_1545 ();
 b15zdnd11an1n64x5 FILLER_232_1609 ();
 b15zdnd11an1n64x5 FILLER_232_1673 ();
 b15zdnd11an1n64x5 FILLER_232_1737 ();
 b15zdnd11an1n64x5 FILLER_232_1801 ();
 b15zdnd11an1n64x5 FILLER_232_1865 ();
 b15zdnd11an1n64x5 FILLER_232_1929 ();
 b15zdnd11an1n64x5 FILLER_232_1993 ();
 b15zdnd11an1n64x5 FILLER_232_2057 ();
 b15zdnd11an1n32x5 FILLER_232_2121 ();
 b15zdnd00an1n01x5 FILLER_232_2153 ();
 b15zdnd11an1n64x5 FILLER_232_2162 ();
 b15zdnd11an1n32x5 FILLER_232_2226 ();
 b15zdnd11an1n16x5 FILLER_232_2258 ();
 b15zdnd00an1n02x5 FILLER_232_2274 ();
 b15zdnd11an1n64x5 FILLER_233_0 ();
 b15zdnd11an1n64x5 FILLER_233_64 ();
 b15zdnd11an1n64x5 FILLER_233_128 ();
 b15zdnd11an1n64x5 FILLER_233_192 ();
 b15zdnd11an1n64x5 FILLER_233_256 ();
 b15zdnd11an1n64x5 FILLER_233_320 ();
 b15zdnd11an1n64x5 FILLER_233_384 ();
 b15zdnd11an1n64x5 FILLER_233_448 ();
 b15zdnd11an1n64x5 FILLER_233_512 ();
 b15zdnd11an1n64x5 FILLER_233_576 ();
 b15zdnd11an1n64x5 FILLER_233_640 ();
 b15zdnd11an1n64x5 FILLER_233_704 ();
 b15zdnd11an1n64x5 FILLER_233_768 ();
 b15zdnd11an1n64x5 FILLER_233_832 ();
 b15zdnd11an1n64x5 FILLER_233_896 ();
 b15zdnd11an1n64x5 FILLER_233_960 ();
 b15zdnd11an1n64x5 FILLER_233_1024 ();
 b15zdnd11an1n64x5 FILLER_233_1088 ();
 b15zdnd11an1n64x5 FILLER_233_1152 ();
 b15zdnd11an1n64x5 FILLER_233_1216 ();
 b15zdnd11an1n64x5 FILLER_233_1280 ();
 b15zdnd11an1n64x5 FILLER_233_1344 ();
 b15zdnd11an1n64x5 FILLER_233_1408 ();
 b15zdnd11an1n64x5 FILLER_233_1472 ();
 b15zdnd11an1n64x5 FILLER_233_1536 ();
 b15zdnd11an1n64x5 FILLER_233_1600 ();
 b15zdnd11an1n64x5 FILLER_233_1664 ();
 b15zdnd11an1n64x5 FILLER_233_1728 ();
 b15zdnd11an1n64x5 FILLER_233_1792 ();
 b15zdnd11an1n64x5 FILLER_233_1856 ();
 b15zdnd11an1n64x5 FILLER_233_1920 ();
 b15zdnd11an1n64x5 FILLER_233_1984 ();
 b15zdnd11an1n64x5 FILLER_233_2048 ();
 b15zdnd11an1n64x5 FILLER_233_2112 ();
 b15zdnd11an1n64x5 FILLER_233_2176 ();
 b15zdnd11an1n32x5 FILLER_233_2240 ();
 b15zdnd11an1n08x5 FILLER_233_2272 ();
 b15zdnd11an1n04x5 FILLER_233_2280 ();
 b15zdnd11an1n64x5 FILLER_234_8 ();
 b15zdnd11an1n64x5 FILLER_234_72 ();
 b15zdnd11an1n64x5 FILLER_234_136 ();
 b15zdnd11an1n64x5 FILLER_234_200 ();
 b15zdnd11an1n64x5 FILLER_234_264 ();
 b15zdnd11an1n64x5 FILLER_234_328 ();
 b15zdnd11an1n64x5 FILLER_234_392 ();
 b15zdnd11an1n64x5 FILLER_234_456 ();
 b15zdnd11an1n64x5 FILLER_234_520 ();
 b15zdnd11an1n64x5 FILLER_234_584 ();
 b15zdnd11an1n64x5 FILLER_234_648 ();
 b15zdnd11an1n04x5 FILLER_234_712 ();
 b15zdnd00an1n02x5 FILLER_234_716 ();
 b15zdnd11an1n64x5 FILLER_234_726 ();
 b15zdnd11an1n32x5 FILLER_234_790 ();
 b15zdnd11an1n16x5 FILLER_234_822 ();
 b15zdnd11an1n08x5 FILLER_234_838 ();
 b15zdnd00an1n01x5 FILLER_234_846 ();
 b15zdnd11an1n64x5 FILLER_234_854 ();
 b15zdnd11an1n64x5 FILLER_234_918 ();
 b15zdnd11an1n64x5 FILLER_234_982 ();
 b15zdnd11an1n64x5 FILLER_234_1046 ();
 b15zdnd11an1n64x5 FILLER_234_1110 ();
 b15zdnd11an1n64x5 FILLER_234_1174 ();
 b15zdnd11an1n64x5 FILLER_234_1238 ();
 b15zdnd11an1n64x5 FILLER_234_1302 ();
 b15zdnd11an1n64x5 FILLER_234_1366 ();
 b15zdnd11an1n64x5 FILLER_234_1430 ();
 b15zdnd11an1n64x5 FILLER_234_1494 ();
 b15zdnd11an1n64x5 FILLER_234_1558 ();
 b15zdnd11an1n64x5 FILLER_234_1622 ();
 b15zdnd11an1n64x5 FILLER_234_1686 ();
 b15zdnd11an1n64x5 FILLER_234_1750 ();
 b15zdnd11an1n64x5 FILLER_234_1814 ();
 b15zdnd11an1n64x5 FILLER_234_1878 ();
 b15zdnd11an1n64x5 FILLER_234_1942 ();
 b15zdnd11an1n64x5 FILLER_234_2006 ();
 b15zdnd11an1n64x5 FILLER_234_2070 ();
 b15zdnd11an1n16x5 FILLER_234_2134 ();
 b15zdnd11an1n04x5 FILLER_234_2150 ();
 b15zdnd11an1n64x5 FILLER_234_2162 ();
 b15zdnd11an1n32x5 FILLER_234_2226 ();
 b15zdnd11an1n16x5 FILLER_234_2258 ();
 b15zdnd00an1n02x5 FILLER_234_2274 ();
 b15zdnd11an1n64x5 FILLER_235_0 ();
 b15zdnd11an1n64x5 FILLER_235_64 ();
 b15zdnd11an1n64x5 FILLER_235_128 ();
 b15zdnd11an1n64x5 FILLER_235_192 ();
 b15zdnd11an1n64x5 FILLER_235_256 ();
 b15zdnd11an1n64x5 FILLER_235_320 ();
 b15zdnd11an1n64x5 FILLER_235_384 ();
 b15zdnd11an1n64x5 FILLER_235_448 ();
 b15zdnd11an1n64x5 FILLER_235_512 ();
 b15zdnd11an1n64x5 FILLER_235_576 ();
 b15zdnd11an1n64x5 FILLER_235_640 ();
 b15zdnd11an1n64x5 FILLER_235_704 ();
 b15zdnd11an1n64x5 FILLER_235_768 ();
 b15zdnd11an1n64x5 FILLER_235_832 ();
 b15zdnd11an1n64x5 FILLER_235_896 ();
 b15zdnd11an1n64x5 FILLER_235_960 ();
 b15zdnd11an1n64x5 FILLER_235_1024 ();
 b15zdnd11an1n64x5 FILLER_235_1088 ();
 b15zdnd11an1n08x5 FILLER_235_1152 ();
 b15zdnd11an1n04x5 FILLER_235_1160 ();
 b15zdnd00an1n02x5 FILLER_235_1164 ();
 b15zdnd00an1n01x5 FILLER_235_1166 ();
 b15zdnd11an1n64x5 FILLER_235_1180 ();
 b15zdnd11an1n64x5 FILLER_235_1244 ();
 b15zdnd11an1n64x5 FILLER_235_1308 ();
 b15zdnd11an1n64x5 FILLER_235_1372 ();
 b15zdnd11an1n64x5 FILLER_235_1436 ();
 b15zdnd11an1n64x5 FILLER_235_1500 ();
 b15zdnd11an1n64x5 FILLER_235_1564 ();
 b15zdnd11an1n64x5 FILLER_235_1628 ();
 b15zdnd11an1n64x5 FILLER_235_1692 ();
 b15zdnd11an1n64x5 FILLER_235_1756 ();
 b15zdnd11an1n64x5 FILLER_235_1820 ();
 b15zdnd11an1n64x5 FILLER_235_1884 ();
 b15zdnd11an1n64x5 FILLER_235_1948 ();
 b15zdnd11an1n64x5 FILLER_235_2012 ();
 b15zdnd11an1n64x5 FILLER_235_2076 ();
 b15zdnd11an1n64x5 FILLER_235_2140 ();
 b15zdnd11an1n64x5 FILLER_235_2204 ();
 b15zdnd11an1n16x5 FILLER_235_2268 ();
 b15zdnd11an1n64x5 FILLER_236_8 ();
 b15zdnd11an1n64x5 FILLER_236_72 ();
 b15zdnd11an1n64x5 FILLER_236_136 ();
 b15zdnd11an1n64x5 FILLER_236_200 ();
 b15zdnd11an1n64x5 FILLER_236_264 ();
 b15zdnd11an1n64x5 FILLER_236_328 ();
 b15zdnd11an1n64x5 FILLER_236_392 ();
 b15zdnd11an1n64x5 FILLER_236_456 ();
 b15zdnd11an1n64x5 FILLER_236_520 ();
 b15zdnd11an1n64x5 FILLER_236_584 ();
 b15zdnd11an1n64x5 FILLER_236_648 ();
 b15zdnd11an1n04x5 FILLER_236_712 ();
 b15zdnd00an1n02x5 FILLER_236_716 ();
 b15zdnd11an1n64x5 FILLER_236_726 ();
 b15zdnd11an1n64x5 FILLER_236_790 ();
 b15zdnd11an1n64x5 FILLER_236_854 ();
 b15zdnd11an1n64x5 FILLER_236_918 ();
 b15zdnd11an1n64x5 FILLER_236_982 ();
 b15zdnd11an1n64x5 FILLER_236_1046 ();
 b15zdnd11an1n64x5 FILLER_236_1110 ();
 b15zdnd11an1n64x5 FILLER_236_1174 ();
 b15zdnd11an1n64x5 FILLER_236_1238 ();
 b15zdnd11an1n64x5 FILLER_236_1302 ();
 b15zdnd11an1n64x5 FILLER_236_1366 ();
 b15zdnd11an1n64x5 FILLER_236_1430 ();
 b15zdnd11an1n64x5 FILLER_236_1494 ();
 b15zdnd11an1n64x5 FILLER_236_1558 ();
 b15zdnd11an1n64x5 FILLER_236_1622 ();
 b15zdnd11an1n64x5 FILLER_236_1686 ();
 b15zdnd11an1n64x5 FILLER_236_1750 ();
 b15zdnd11an1n64x5 FILLER_236_1814 ();
 b15zdnd11an1n64x5 FILLER_236_1878 ();
 b15zdnd11an1n64x5 FILLER_236_1942 ();
 b15zdnd11an1n64x5 FILLER_236_2006 ();
 b15zdnd11an1n64x5 FILLER_236_2070 ();
 b15zdnd11an1n16x5 FILLER_236_2134 ();
 b15zdnd11an1n04x5 FILLER_236_2150 ();
 b15zdnd11an1n64x5 FILLER_236_2162 ();
 b15zdnd11an1n32x5 FILLER_236_2226 ();
 b15zdnd11an1n16x5 FILLER_236_2258 ();
 b15zdnd00an1n02x5 FILLER_236_2274 ();
 b15zdnd11an1n64x5 FILLER_237_0 ();
 b15zdnd11an1n64x5 FILLER_237_64 ();
 b15zdnd11an1n64x5 FILLER_237_128 ();
 b15zdnd11an1n64x5 FILLER_237_192 ();
 b15zdnd11an1n64x5 FILLER_237_256 ();
 b15zdnd11an1n64x5 FILLER_237_320 ();
 b15zdnd11an1n64x5 FILLER_237_384 ();
 b15zdnd11an1n64x5 FILLER_237_448 ();
 b15zdnd11an1n64x5 FILLER_237_512 ();
 b15zdnd11an1n64x5 FILLER_237_576 ();
 b15zdnd11an1n64x5 FILLER_237_640 ();
 b15zdnd11an1n64x5 FILLER_237_704 ();
 b15zdnd11an1n64x5 FILLER_237_768 ();
 b15zdnd11an1n16x5 FILLER_237_832 ();
 b15zdnd11an1n08x5 FILLER_237_848 ();
 b15zdnd00an1n02x5 FILLER_237_856 ();
 b15zdnd00an1n01x5 FILLER_237_858 ();
 b15zdnd11an1n64x5 FILLER_237_871 ();
 b15zdnd11an1n64x5 FILLER_237_935 ();
 b15zdnd11an1n16x5 FILLER_237_999 ();
 b15zdnd00an1n02x5 FILLER_237_1015 ();
 b15zdnd00an1n01x5 FILLER_237_1017 ();
 b15zdnd11an1n64x5 FILLER_237_1060 ();
 b15zdnd11an1n64x5 FILLER_237_1124 ();
 b15zdnd11an1n64x5 FILLER_237_1188 ();
 b15zdnd11an1n64x5 FILLER_237_1252 ();
 b15zdnd11an1n64x5 FILLER_237_1316 ();
 b15zdnd11an1n64x5 FILLER_237_1380 ();
 b15zdnd11an1n64x5 FILLER_237_1444 ();
 b15zdnd11an1n64x5 FILLER_237_1508 ();
 b15zdnd11an1n64x5 FILLER_237_1572 ();
 b15zdnd11an1n64x5 FILLER_237_1636 ();
 b15zdnd11an1n64x5 FILLER_237_1700 ();
 b15zdnd11an1n64x5 FILLER_237_1764 ();
 b15zdnd11an1n64x5 FILLER_237_1828 ();
 b15zdnd11an1n64x5 FILLER_237_1892 ();
 b15zdnd11an1n64x5 FILLER_237_1956 ();
 b15zdnd11an1n64x5 FILLER_237_2020 ();
 b15zdnd11an1n64x5 FILLER_237_2084 ();
 b15zdnd11an1n64x5 FILLER_237_2148 ();
 b15zdnd11an1n64x5 FILLER_237_2212 ();
 b15zdnd11an1n08x5 FILLER_237_2276 ();
 b15zdnd11an1n64x5 FILLER_238_8 ();
 b15zdnd11an1n64x5 FILLER_238_72 ();
 b15zdnd11an1n64x5 FILLER_238_136 ();
 b15zdnd11an1n64x5 FILLER_238_200 ();
 b15zdnd11an1n64x5 FILLER_238_264 ();
 b15zdnd11an1n64x5 FILLER_238_328 ();
 b15zdnd11an1n64x5 FILLER_238_392 ();
 b15zdnd11an1n64x5 FILLER_238_456 ();
 b15zdnd11an1n64x5 FILLER_238_520 ();
 b15zdnd11an1n64x5 FILLER_238_584 ();
 b15zdnd11an1n64x5 FILLER_238_648 ();
 b15zdnd11an1n04x5 FILLER_238_712 ();
 b15zdnd00an1n02x5 FILLER_238_716 ();
 b15zdnd11an1n64x5 FILLER_238_726 ();
 b15zdnd11an1n64x5 FILLER_238_790 ();
 b15zdnd11an1n64x5 FILLER_238_854 ();
 b15zdnd11an1n64x5 FILLER_238_918 ();
 b15zdnd11an1n64x5 FILLER_238_982 ();
 b15zdnd11an1n64x5 FILLER_238_1046 ();
 b15zdnd11an1n64x5 FILLER_238_1110 ();
 b15zdnd11an1n64x5 FILLER_238_1174 ();
 b15zdnd11an1n64x5 FILLER_238_1238 ();
 b15zdnd11an1n64x5 FILLER_238_1302 ();
 b15zdnd11an1n64x5 FILLER_238_1366 ();
 b15zdnd11an1n64x5 FILLER_238_1430 ();
 b15zdnd11an1n64x5 FILLER_238_1494 ();
 b15zdnd11an1n64x5 FILLER_238_1558 ();
 b15zdnd11an1n64x5 FILLER_238_1622 ();
 b15zdnd11an1n64x5 FILLER_238_1686 ();
 b15zdnd11an1n64x5 FILLER_238_1750 ();
 b15zdnd11an1n64x5 FILLER_238_1814 ();
 b15zdnd11an1n64x5 FILLER_238_1878 ();
 b15zdnd11an1n64x5 FILLER_238_1942 ();
 b15zdnd11an1n64x5 FILLER_238_2006 ();
 b15zdnd11an1n64x5 FILLER_238_2070 ();
 b15zdnd11an1n16x5 FILLER_238_2134 ();
 b15zdnd11an1n04x5 FILLER_238_2150 ();
 b15zdnd11an1n64x5 FILLER_238_2162 ();
 b15zdnd11an1n32x5 FILLER_238_2226 ();
 b15zdnd11an1n16x5 FILLER_238_2258 ();
 b15zdnd00an1n02x5 FILLER_238_2274 ();
 b15zdnd11an1n64x5 FILLER_239_0 ();
 b15zdnd11an1n64x5 FILLER_239_64 ();
 b15zdnd11an1n64x5 FILLER_239_128 ();
 b15zdnd11an1n64x5 FILLER_239_192 ();
 b15zdnd11an1n64x5 FILLER_239_256 ();
 b15zdnd11an1n64x5 FILLER_239_320 ();
 b15zdnd11an1n64x5 FILLER_239_384 ();
 b15zdnd11an1n64x5 FILLER_239_448 ();
 b15zdnd11an1n64x5 FILLER_239_512 ();
 b15zdnd11an1n64x5 FILLER_239_576 ();
 b15zdnd11an1n64x5 FILLER_239_640 ();
 b15zdnd11an1n64x5 FILLER_239_704 ();
 b15zdnd11an1n64x5 FILLER_239_768 ();
 b15zdnd11an1n64x5 FILLER_239_832 ();
 b15zdnd11an1n64x5 FILLER_239_896 ();
 b15zdnd11an1n64x5 FILLER_239_960 ();
 b15zdnd11an1n64x5 FILLER_239_1024 ();
 b15zdnd11an1n64x5 FILLER_239_1088 ();
 b15zdnd11an1n64x5 FILLER_239_1152 ();
 b15zdnd11an1n64x5 FILLER_239_1216 ();
 b15zdnd11an1n64x5 FILLER_239_1280 ();
 b15zdnd11an1n64x5 FILLER_239_1344 ();
 b15zdnd11an1n64x5 FILLER_239_1408 ();
 b15zdnd11an1n64x5 FILLER_239_1472 ();
 b15zdnd11an1n64x5 FILLER_239_1536 ();
 b15zdnd11an1n64x5 FILLER_239_1600 ();
 b15zdnd11an1n64x5 FILLER_239_1664 ();
 b15zdnd11an1n64x5 FILLER_239_1728 ();
 b15zdnd11an1n64x5 FILLER_239_1792 ();
 b15zdnd11an1n64x5 FILLER_239_1856 ();
 b15zdnd11an1n64x5 FILLER_239_1920 ();
 b15zdnd11an1n64x5 FILLER_239_1984 ();
 b15zdnd11an1n64x5 FILLER_239_2048 ();
 b15zdnd11an1n64x5 FILLER_239_2112 ();
 b15zdnd11an1n64x5 FILLER_239_2176 ();
 b15zdnd11an1n32x5 FILLER_239_2240 ();
 b15zdnd11an1n08x5 FILLER_239_2272 ();
 b15zdnd11an1n04x5 FILLER_239_2280 ();
 b15zdnd11an1n64x5 FILLER_240_8 ();
 b15zdnd11an1n64x5 FILLER_240_72 ();
 b15zdnd11an1n64x5 FILLER_240_136 ();
 b15zdnd11an1n64x5 FILLER_240_200 ();
 b15zdnd11an1n64x5 FILLER_240_264 ();
 b15zdnd11an1n64x5 FILLER_240_328 ();
 b15zdnd11an1n64x5 FILLER_240_392 ();
 b15zdnd11an1n64x5 FILLER_240_456 ();
 b15zdnd11an1n64x5 FILLER_240_520 ();
 b15zdnd11an1n64x5 FILLER_240_584 ();
 b15zdnd11an1n64x5 FILLER_240_648 ();
 b15zdnd11an1n04x5 FILLER_240_712 ();
 b15zdnd00an1n02x5 FILLER_240_716 ();
 b15zdnd11an1n64x5 FILLER_240_726 ();
 b15zdnd11an1n64x5 FILLER_240_790 ();
 b15zdnd11an1n64x5 FILLER_240_854 ();
 b15zdnd11an1n64x5 FILLER_240_918 ();
 b15zdnd11an1n64x5 FILLER_240_982 ();
 b15zdnd11an1n64x5 FILLER_240_1046 ();
 b15zdnd11an1n64x5 FILLER_240_1110 ();
 b15zdnd11an1n64x5 FILLER_240_1174 ();
 b15zdnd11an1n64x5 FILLER_240_1238 ();
 b15zdnd11an1n64x5 FILLER_240_1302 ();
 b15zdnd11an1n64x5 FILLER_240_1366 ();
 b15zdnd11an1n64x5 FILLER_240_1430 ();
 b15zdnd11an1n64x5 FILLER_240_1494 ();
 b15zdnd11an1n64x5 FILLER_240_1558 ();
 b15zdnd11an1n64x5 FILLER_240_1622 ();
 b15zdnd11an1n64x5 FILLER_240_1686 ();
 b15zdnd11an1n64x5 FILLER_240_1750 ();
 b15zdnd11an1n64x5 FILLER_240_1814 ();
 b15zdnd11an1n64x5 FILLER_240_1878 ();
 b15zdnd11an1n64x5 FILLER_240_1942 ();
 b15zdnd11an1n64x5 FILLER_240_2006 ();
 b15zdnd11an1n32x5 FILLER_240_2070 ();
 b15zdnd11an1n04x5 FILLER_240_2102 ();
 b15zdnd11an1n32x5 FILLER_240_2122 ();
 b15zdnd11an1n64x5 FILLER_240_2162 ();
 b15zdnd11an1n32x5 FILLER_240_2226 ();
 b15zdnd11an1n16x5 FILLER_240_2258 ();
 b15zdnd00an1n02x5 FILLER_240_2274 ();
 b15zdnd11an1n64x5 FILLER_241_0 ();
 b15zdnd11an1n64x5 FILLER_241_64 ();
 b15zdnd11an1n64x5 FILLER_241_128 ();
 b15zdnd11an1n64x5 FILLER_241_192 ();
 b15zdnd11an1n64x5 FILLER_241_256 ();
 b15zdnd11an1n64x5 FILLER_241_320 ();
 b15zdnd11an1n64x5 FILLER_241_384 ();
 b15zdnd11an1n64x5 FILLER_241_448 ();
 b15zdnd11an1n64x5 FILLER_241_512 ();
 b15zdnd11an1n64x5 FILLER_241_576 ();
 b15zdnd11an1n64x5 FILLER_241_640 ();
 b15zdnd11an1n64x5 FILLER_241_704 ();
 b15zdnd11an1n64x5 FILLER_241_768 ();
 b15zdnd11an1n64x5 FILLER_241_832 ();
 b15zdnd11an1n64x5 FILLER_241_896 ();
 b15zdnd11an1n64x5 FILLER_241_960 ();
 b15zdnd11an1n64x5 FILLER_241_1024 ();
 b15zdnd11an1n64x5 FILLER_241_1088 ();
 b15zdnd11an1n64x5 FILLER_241_1152 ();
 b15zdnd11an1n64x5 FILLER_241_1216 ();
 b15zdnd11an1n64x5 FILLER_241_1280 ();
 b15zdnd11an1n64x5 FILLER_241_1344 ();
 b15zdnd11an1n64x5 FILLER_241_1408 ();
 b15zdnd11an1n64x5 FILLER_241_1472 ();
 b15zdnd11an1n64x5 FILLER_241_1536 ();
 b15zdnd11an1n64x5 FILLER_241_1600 ();
 b15zdnd11an1n64x5 FILLER_241_1664 ();
 b15zdnd11an1n64x5 FILLER_241_1728 ();
 b15zdnd11an1n64x5 FILLER_241_1792 ();
 b15zdnd11an1n64x5 FILLER_241_1856 ();
 b15zdnd11an1n64x5 FILLER_241_1920 ();
 b15zdnd11an1n64x5 FILLER_241_1984 ();
 b15zdnd11an1n64x5 FILLER_241_2048 ();
 b15zdnd11an1n64x5 FILLER_241_2112 ();
 b15zdnd11an1n64x5 FILLER_241_2176 ();
 b15zdnd11an1n32x5 FILLER_241_2240 ();
 b15zdnd11an1n08x5 FILLER_241_2272 ();
 b15zdnd11an1n04x5 FILLER_241_2280 ();
 b15zdnd11an1n64x5 FILLER_242_8 ();
 b15zdnd11an1n64x5 FILLER_242_72 ();
 b15zdnd11an1n64x5 FILLER_242_136 ();
 b15zdnd11an1n64x5 FILLER_242_200 ();
 b15zdnd11an1n64x5 FILLER_242_264 ();
 b15zdnd11an1n64x5 FILLER_242_328 ();
 b15zdnd11an1n64x5 FILLER_242_392 ();
 b15zdnd11an1n64x5 FILLER_242_456 ();
 b15zdnd11an1n64x5 FILLER_242_520 ();
 b15zdnd11an1n64x5 FILLER_242_584 ();
 b15zdnd11an1n64x5 FILLER_242_648 ();
 b15zdnd11an1n04x5 FILLER_242_712 ();
 b15zdnd00an1n02x5 FILLER_242_716 ();
 b15zdnd11an1n64x5 FILLER_242_726 ();
 b15zdnd11an1n64x5 FILLER_242_790 ();
 b15zdnd11an1n64x5 FILLER_242_854 ();
 b15zdnd11an1n64x5 FILLER_242_918 ();
 b15zdnd11an1n64x5 FILLER_242_982 ();
 b15zdnd11an1n64x5 FILLER_242_1046 ();
 b15zdnd11an1n64x5 FILLER_242_1110 ();
 b15zdnd11an1n64x5 FILLER_242_1174 ();
 b15zdnd11an1n64x5 FILLER_242_1238 ();
 b15zdnd11an1n64x5 FILLER_242_1302 ();
 b15zdnd11an1n64x5 FILLER_242_1366 ();
 b15zdnd11an1n64x5 FILLER_242_1430 ();
 b15zdnd11an1n64x5 FILLER_242_1494 ();
 b15zdnd11an1n64x5 FILLER_242_1558 ();
 b15zdnd11an1n64x5 FILLER_242_1622 ();
 b15zdnd11an1n64x5 FILLER_242_1686 ();
 b15zdnd11an1n64x5 FILLER_242_1750 ();
 b15zdnd11an1n64x5 FILLER_242_1814 ();
 b15zdnd11an1n64x5 FILLER_242_1878 ();
 b15zdnd11an1n64x5 FILLER_242_1942 ();
 b15zdnd11an1n64x5 FILLER_242_2006 ();
 b15zdnd11an1n64x5 FILLER_242_2070 ();
 b15zdnd11an1n16x5 FILLER_242_2134 ();
 b15zdnd11an1n04x5 FILLER_242_2150 ();
 b15zdnd11an1n64x5 FILLER_242_2162 ();
 b15zdnd11an1n32x5 FILLER_242_2226 ();
 b15zdnd11an1n16x5 FILLER_242_2258 ();
 b15zdnd00an1n02x5 FILLER_242_2274 ();
 b15zdnd11an1n64x5 FILLER_243_0 ();
 b15zdnd11an1n64x5 FILLER_243_64 ();
 b15zdnd11an1n64x5 FILLER_243_128 ();
 b15zdnd11an1n64x5 FILLER_243_192 ();
 b15zdnd11an1n64x5 FILLER_243_256 ();
 b15zdnd11an1n64x5 FILLER_243_320 ();
 b15zdnd11an1n64x5 FILLER_243_384 ();
 b15zdnd11an1n64x5 FILLER_243_448 ();
 b15zdnd11an1n64x5 FILLER_243_512 ();
 b15zdnd11an1n64x5 FILLER_243_576 ();
 b15zdnd11an1n64x5 FILLER_243_640 ();
 b15zdnd11an1n64x5 FILLER_243_704 ();
 b15zdnd11an1n64x5 FILLER_243_768 ();
 b15zdnd11an1n64x5 FILLER_243_832 ();
 b15zdnd11an1n64x5 FILLER_243_896 ();
 b15zdnd11an1n64x5 FILLER_243_960 ();
 b15zdnd11an1n64x5 FILLER_243_1024 ();
 b15zdnd11an1n64x5 FILLER_243_1088 ();
 b15zdnd11an1n64x5 FILLER_243_1152 ();
 b15zdnd11an1n64x5 FILLER_243_1216 ();
 b15zdnd11an1n64x5 FILLER_243_1280 ();
 b15zdnd11an1n64x5 FILLER_243_1344 ();
 b15zdnd11an1n64x5 FILLER_243_1408 ();
 b15zdnd11an1n64x5 FILLER_243_1472 ();
 b15zdnd11an1n64x5 FILLER_243_1536 ();
 b15zdnd11an1n64x5 FILLER_243_1600 ();
 b15zdnd11an1n64x5 FILLER_243_1664 ();
 b15zdnd11an1n64x5 FILLER_243_1728 ();
 b15zdnd11an1n64x5 FILLER_243_1792 ();
 b15zdnd11an1n64x5 FILLER_243_1856 ();
 b15zdnd11an1n64x5 FILLER_243_1920 ();
 b15zdnd11an1n64x5 FILLER_243_1984 ();
 b15zdnd11an1n64x5 FILLER_243_2048 ();
 b15zdnd11an1n64x5 FILLER_243_2112 ();
 b15zdnd11an1n64x5 FILLER_243_2176 ();
 b15zdnd11an1n32x5 FILLER_243_2240 ();
 b15zdnd11an1n08x5 FILLER_243_2272 ();
 b15zdnd11an1n04x5 FILLER_243_2280 ();
 b15zdnd11an1n64x5 FILLER_244_8 ();
 b15zdnd11an1n64x5 FILLER_244_72 ();
 b15zdnd11an1n64x5 FILLER_244_136 ();
 b15zdnd11an1n64x5 FILLER_244_200 ();
 b15zdnd11an1n64x5 FILLER_244_264 ();
 b15zdnd11an1n64x5 FILLER_244_328 ();
 b15zdnd11an1n64x5 FILLER_244_392 ();
 b15zdnd11an1n64x5 FILLER_244_456 ();
 b15zdnd11an1n64x5 FILLER_244_520 ();
 b15zdnd11an1n64x5 FILLER_244_584 ();
 b15zdnd11an1n64x5 FILLER_244_648 ();
 b15zdnd11an1n04x5 FILLER_244_712 ();
 b15zdnd00an1n02x5 FILLER_244_716 ();
 b15zdnd11an1n64x5 FILLER_244_726 ();
 b15zdnd11an1n64x5 FILLER_244_790 ();
 b15zdnd11an1n64x5 FILLER_244_854 ();
 b15zdnd11an1n64x5 FILLER_244_918 ();
 b15zdnd11an1n64x5 FILLER_244_982 ();
 b15zdnd11an1n64x5 FILLER_244_1046 ();
 b15zdnd11an1n64x5 FILLER_244_1110 ();
 b15zdnd11an1n64x5 FILLER_244_1174 ();
 b15zdnd11an1n64x5 FILLER_244_1238 ();
 b15zdnd11an1n64x5 FILLER_244_1302 ();
 b15zdnd11an1n64x5 FILLER_244_1366 ();
 b15zdnd11an1n64x5 FILLER_244_1430 ();
 b15zdnd11an1n64x5 FILLER_244_1494 ();
 b15zdnd11an1n64x5 FILLER_244_1558 ();
 b15zdnd11an1n64x5 FILLER_244_1622 ();
 b15zdnd11an1n64x5 FILLER_244_1686 ();
 b15zdnd11an1n64x5 FILLER_244_1750 ();
 b15zdnd11an1n64x5 FILLER_244_1814 ();
 b15zdnd11an1n64x5 FILLER_244_1878 ();
 b15zdnd11an1n64x5 FILLER_244_1942 ();
 b15zdnd11an1n64x5 FILLER_244_2006 ();
 b15zdnd11an1n64x5 FILLER_244_2070 ();
 b15zdnd11an1n16x5 FILLER_244_2134 ();
 b15zdnd11an1n04x5 FILLER_244_2150 ();
 b15zdnd11an1n64x5 FILLER_244_2162 ();
 b15zdnd11an1n32x5 FILLER_244_2226 ();
 b15zdnd11an1n16x5 FILLER_244_2258 ();
 b15zdnd00an1n02x5 FILLER_244_2274 ();
 b15zdnd11an1n64x5 FILLER_245_0 ();
 b15zdnd11an1n64x5 FILLER_245_64 ();
 b15zdnd11an1n64x5 FILLER_245_128 ();
 b15zdnd11an1n64x5 FILLER_245_192 ();
 b15zdnd11an1n64x5 FILLER_245_256 ();
 b15zdnd11an1n64x5 FILLER_245_320 ();
 b15zdnd11an1n64x5 FILLER_245_384 ();
 b15zdnd11an1n64x5 FILLER_245_448 ();
 b15zdnd11an1n64x5 FILLER_245_512 ();
 b15zdnd11an1n64x5 FILLER_245_576 ();
 b15zdnd11an1n64x5 FILLER_245_640 ();
 b15zdnd11an1n64x5 FILLER_245_704 ();
 b15zdnd11an1n64x5 FILLER_245_768 ();
 b15zdnd11an1n64x5 FILLER_245_832 ();
 b15zdnd11an1n64x5 FILLER_245_896 ();
 b15zdnd11an1n64x5 FILLER_245_960 ();
 b15zdnd11an1n64x5 FILLER_245_1024 ();
 b15zdnd11an1n64x5 FILLER_245_1088 ();
 b15zdnd11an1n64x5 FILLER_245_1152 ();
 b15zdnd11an1n64x5 FILLER_245_1216 ();
 b15zdnd11an1n64x5 FILLER_245_1280 ();
 b15zdnd11an1n64x5 FILLER_245_1344 ();
 b15zdnd11an1n64x5 FILLER_245_1408 ();
 b15zdnd11an1n64x5 FILLER_245_1472 ();
 b15zdnd11an1n64x5 FILLER_245_1536 ();
 b15zdnd11an1n64x5 FILLER_245_1600 ();
 b15zdnd11an1n64x5 FILLER_245_1664 ();
 b15zdnd11an1n64x5 FILLER_245_1728 ();
 b15zdnd11an1n64x5 FILLER_245_1792 ();
 b15zdnd11an1n64x5 FILLER_245_1856 ();
 b15zdnd11an1n64x5 FILLER_245_1920 ();
 b15zdnd11an1n64x5 FILLER_245_1984 ();
 b15zdnd11an1n64x5 FILLER_245_2048 ();
 b15zdnd11an1n64x5 FILLER_245_2112 ();
 b15zdnd11an1n64x5 FILLER_245_2176 ();
 b15zdnd11an1n32x5 FILLER_245_2240 ();
 b15zdnd11an1n08x5 FILLER_245_2272 ();
 b15zdnd11an1n04x5 FILLER_245_2280 ();
 b15zdnd11an1n64x5 FILLER_246_8 ();
 b15zdnd11an1n64x5 FILLER_246_72 ();
 b15zdnd11an1n64x5 FILLER_246_136 ();
 b15zdnd11an1n64x5 FILLER_246_200 ();
 b15zdnd11an1n64x5 FILLER_246_264 ();
 b15zdnd11an1n64x5 FILLER_246_328 ();
 b15zdnd11an1n64x5 FILLER_246_392 ();
 b15zdnd11an1n64x5 FILLER_246_456 ();
 b15zdnd11an1n64x5 FILLER_246_520 ();
 b15zdnd11an1n64x5 FILLER_246_584 ();
 b15zdnd11an1n64x5 FILLER_246_648 ();
 b15zdnd11an1n04x5 FILLER_246_712 ();
 b15zdnd00an1n02x5 FILLER_246_716 ();
 b15zdnd11an1n64x5 FILLER_246_726 ();
 b15zdnd11an1n64x5 FILLER_246_790 ();
 b15zdnd11an1n64x5 FILLER_246_854 ();
 b15zdnd11an1n64x5 FILLER_246_918 ();
 b15zdnd11an1n64x5 FILLER_246_982 ();
 b15zdnd11an1n64x5 FILLER_246_1046 ();
 b15zdnd11an1n64x5 FILLER_246_1110 ();
 b15zdnd11an1n64x5 FILLER_246_1174 ();
 b15zdnd11an1n64x5 FILLER_246_1238 ();
 b15zdnd11an1n64x5 FILLER_246_1302 ();
 b15zdnd11an1n64x5 FILLER_246_1366 ();
 b15zdnd11an1n64x5 FILLER_246_1430 ();
 b15zdnd11an1n64x5 FILLER_246_1494 ();
 b15zdnd11an1n64x5 FILLER_246_1558 ();
 b15zdnd11an1n64x5 FILLER_246_1622 ();
 b15zdnd11an1n64x5 FILLER_246_1686 ();
 b15zdnd11an1n64x5 FILLER_246_1750 ();
 b15zdnd11an1n64x5 FILLER_246_1814 ();
 b15zdnd11an1n64x5 FILLER_246_1878 ();
 b15zdnd11an1n64x5 FILLER_246_1942 ();
 b15zdnd11an1n64x5 FILLER_246_2006 ();
 b15zdnd11an1n64x5 FILLER_246_2070 ();
 b15zdnd11an1n16x5 FILLER_246_2134 ();
 b15zdnd11an1n04x5 FILLER_246_2150 ();
 b15zdnd11an1n64x5 FILLER_246_2162 ();
 b15zdnd11an1n32x5 FILLER_246_2226 ();
 b15zdnd11an1n16x5 FILLER_246_2258 ();
 b15zdnd00an1n02x5 FILLER_246_2274 ();
 b15zdnd11an1n64x5 FILLER_247_0 ();
 b15zdnd11an1n64x5 FILLER_247_64 ();
 b15zdnd11an1n64x5 FILLER_247_128 ();
 b15zdnd11an1n64x5 FILLER_247_192 ();
 b15zdnd11an1n64x5 FILLER_247_256 ();
 b15zdnd11an1n64x5 FILLER_247_320 ();
 b15zdnd11an1n64x5 FILLER_247_384 ();
 b15zdnd11an1n64x5 FILLER_247_448 ();
 b15zdnd11an1n64x5 FILLER_247_512 ();
 b15zdnd11an1n64x5 FILLER_247_576 ();
 b15zdnd11an1n64x5 FILLER_247_640 ();
 b15zdnd11an1n64x5 FILLER_247_704 ();
 b15zdnd11an1n64x5 FILLER_247_768 ();
 b15zdnd11an1n64x5 FILLER_247_832 ();
 b15zdnd11an1n64x5 FILLER_247_896 ();
 b15zdnd11an1n64x5 FILLER_247_960 ();
 b15zdnd11an1n64x5 FILLER_247_1024 ();
 b15zdnd11an1n64x5 FILLER_247_1088 ();
 b15zdnd11an1n64x5 FILLER_247_1152 ();
 b15zdnd11an1n64x5 FILLER_247_1216 ();
 b15zdnd11an1n64x5 FILLER_247_1280 ();
 b15zdnd11an1n64x5 FILLER_247_1344 ();
 b15zdnd11an1n64x5 FILLER_247_1408 ();
 b15zdnd11an1n64x5 FILLER_247_1472 ();
 b15zdnd11an1n64x5 FILLER_247_1536 ();
 b15zdnd11an1n64x5 FILLER_247_1600 ();
 b15zdnd11an1n64x5 FILLER_247_1664 ();
 b15zdnd11an1n64x5 FILLER_247_1728 ();
 b15zdnd11an1n64x5 FILLER_247_1792 ();
 b15zdnd11an1n64x5 FILLER_247_1856 ();
 b15zdnd11an1n64x5 FILLER_247_1920 ();
 b15zdnd11an1n64x5 FILLER_247_1984 ();
 b15zdnd11an1n32x5 FILLER_247_2048 ();
 b15zdnd11an1n16x5 FILLER_247_2080 ();
 b15zdnd11an1n08x5 FILLER_247_2096 ();
 b15zdnd00an1n02x5 FILLER_247_2104 ();
 b15zdnd00an1n01x5 FILLER_247_2106 ();
 b15zdnd11an1n64x5 FILLER_247_2123 ();
 b15zdnd11an1n64x5 FILLER_247_2187 ();
 b15zdnd11an1n32x5 FILLER_247_2251 ();
 b15zdnd00an1n01x5 FILLER_247_2283 ();
 b15zdnd11an1n64x5 FILLER_248_8 ();
 b15zdnd11an1n64x5 FILLER_248_72 ();
 b15zdnd11an1n64x5 FILLER_248_136 ();
 b15zdnd11an1n64x5 FILLER_248_200 ();
 b15zdnd11an1n64x5 FILLER_248_264 ();
 b15zdnd11an1n64x5 FILLER_248_328 ();
 b15zdnd11an1n64x5 FILLER_248_392 ();
 b15zdnd11an1n64x5 FILLER_248_456 ();
 b15zdnd11an1n64x5 FILLER_248_520 ();
 b15zdnd11an1n64x5 FILLER_248_584 ();
 b15zdnd11an1n64x5 FILLER_248_648 ();
 b15zdnd11an1n04x5 FILLER_248_712 ();
 b15zdnd00an1n02x5 FILLER_248_716 ();
 b15zdnd11an1n64x5 FILLER_248_726 ();
 b15zdnd11an1n64x5 FILLER_248_790 ();
 b15zdnd11an1n64x5 FILLER_248_854 ();
 b15zdnd11an1n64x5 FILLER_248_918 ();
 b15zdnd11an1n64x5 FILLER_248_982 ();
 b15zdnd11an1n64x5 FILLER_248_1046 ();
 b15zdnd11an1n64x5 FILLER_248_1110 ();
 b15zdnd11an1n64x5 FILLER_248_1174 ();
 b15zdnd11an1n64x5 FILLER_248_1238 ();
 b15zdnd11an1n64x5 FILLER_248_1302 ();
 b15zdnd11an1n64x5 FILLER_248_1366 ();
 b15zdnd11an1n64x5 FILLER_248_1430 ();
 b15zdnd11an1n64x5 FILLER_248_1494 ();
 b15zdnd11an1n64x5 FILLER_248_1558 ();
 b15zdnd11an1n64x5 FILLER_248_1622 ();
 b15zdnd11an1n64x5 FILLER_248_1686 ();
 b15zdnd11an1n64x5 FILLER_248_1750 ();
 b15zdnd11an1n64x5 FILLER_248_1814 ();
 b15zdnd11an1n64x5 FILLER_248_1878 ();
 b15zdnd11an1n64x5 FILLER_248_1942 ();
 b15zdnd11an1n64x5 FILLER_248_2006 ();
 b15zdnd11an1n64x5 FILLER_248_2070 ();
 b15zdnd11an1n16x5 FILLER_248_2134 ();
 b15zdnd11an1n04x5 FILLER_248_2150 ();
 b15zdnd11an1n64x5 FILLER_248_2162 ();
 b15zdnd11an1n32x5 FILLER_248_2226 ();
 b15zdnd11an1n16x5 FILLER_248_2258 ();
 b15zdnd00an1n02x5 FILLER_248_2274 ();
 b15zdnd11an1n64x5 FILLER_249_0 ();
 b15zdnd11an1n64x5 FILLER_249_64 ();
 b15zdnd11an1n64x5 FILLER_249_128 ();
 b15zdnd11an1n64x5 FILLER_249_192 ();
 b15zdnd11an1n64x5 FILLER_249_256 ();
 b15zdnd11an1n64x5 FILLER_249_320 ();
 b15zdnd11an1n64x5 FILLER_249_384 ();
 b15zdnd11an1n64x5 FILLER_249_448 ();
 b15zdnd11an1n64x5 FILLER_249_512 ();
 b15zdnd11an1n64x5 FILLER_249_576 ();
 b15zdnd11an1n64x5 FILLER_249_640 ();
 b15zdnd11an1n64x5 FILLER_249_704 ();
 b15zdnd11an1n64x5 FILLER_249_768 ();
 b15zdnd11an1n64x5 FILLER_249_832 ();
 b15zdnd11an1n64x5 FILLER_249_896 ();
 b15zdnd11an1n64x5 FILLER_249_960 ();
 b15zdnd11an1n64x5 FILLER_249_1024 ();
 b15zdnd11an1n64x5 FILLER_249_1088 ();
 b15zdnd11an1n64x5 FILLER_249_1152 ();
 b15zdnd11an1n64x5 FILLER_249_1216 ();
 b15zdnd11an1n64x5 FILLER_249_1280 ();
 b15zdnd11an1n64x5 FILLER_249_1344 ();
 b15zdnd11an1n64x5 FILLER_249_1408 ();
 b15zdnd11an1n64x5 FILLER_249_1472 ();
 b15zdnd11an1n64x5 FILLER_249_1536 ();
 b15zdnd11an1n64x5 FILLER_249_1600 ();
 b15zdnd11an1n64x5 FILLER_249_1664 ();
 b15zdnd11an1n64x5 FILLER_249_1728 ();
 b15zdnd11an1n64x5 FILLER_249_1792 ();
 b15zdnd11an1n64x5 FILLER_249_1856 ();
 b15zdnd11an1n64x5 FILLER_249_1920 ();
 b15zdnd11an1n64x5 FILLER_249_1984 ();
 b15zdnd11an1n64x5 FILLER_249_2048 ();
 b15zdnd11an1n64x5 FILLER_249_2112 ();
 b15zdnd11an1n64x5 FILLER_249_2176 ();
 b15zdnd11an1n32x5 FILLER_249_2240 ();
 b15zdnd11an1n08x5 FILLER_249_2272 ();
 b15zdnd11an1n04x5 FILLER_249_2280 ();
 b15zdnd11an1n64x5 FILLER_250_8 ();
 b15zdnd11an1n64x5 FILLER_250_72 ();
 b15zdnd11an1n64x5 FILLER_250_136 ();
 b15zdnd11an1n64x5 FILLER_250_200 ();
 b15zdnd11an1n64x5 FILLER_250_264 ();
 b15zdnd11an1n64x5 FILLER_250_328 ();
 b15zdnd11an1n64x5 FILLER_250_392 ();
 b15zdnd11an1n64x5 FILLER_250_456 ();
 b15zdnd11an1n64x5 FILLER_250_520 ();
 b15zdnd11an1n64x5 FILLER_250_584 ();
 b15zdnd11an1n64x5 FILLER_250_648 ();
 b15zdnd11an1n04x5 FILLER_250_712 ();
 b15zdnd00an1n02x5 FILLER_250_716 ();
 b15zdnd11an1n64x5 FILLER_250_726 ();
 b15zdnd11an1n64x5 FILLER_250_790 ();
 b15zdnd11an1n64x5 FILLER_250_854 ();
 b15zdnd11an1n64x5 FILLER_250_918 ();
 b15zdnd11an1n64x5 FILLER_250_982 ();
 b15zdnd11an1n64x5 FILLER_250_1046 ();
 b15zdnd11an1n64x5 FILLER_250_1110 ();
 b15zdnd11an1n64x5 FILLER_250_1174 ();
 b15zdnd11an1n64x5 FILLER_250_1238 ();
 b15zdnd11an1n64x5 FILLER_250_1302 ();
 b15zdnd11an1n64x5 FILLER_250_1366 ();
 b15zdnd11an1n64x5 FILLER_250_1430 ();
 b15zdnd11an1n64x5 FILLER_250_1494 ();
 b15zdnd11an1n64x5 FILLER_250_1558 ();
 b15zdnd11an1n64x5 FILLER_250_1622 ();
 b15zdnd11an1n64x5 FILLER_250_1686 ();
 b15zdnd11an1n64x5 FILLER_250_1750 ();
 b15zdnd11an1n64x5 FILLER_250_1814 ();
 b15zdnd11an1n64x5 FILLER_250_1878 ();
 b15zdnd11an1n64x5 FILLER_250_1942 ();
 b15zdnd11an1n64x5 FILLER_250_2006 ();
 b15zdnd11an1n64x5 FILLER_250_2070 ();
 b15zdnd11an1n16x5 FILLER_250_2134 ();
 b15zdnd11an1n04x5 FILLER_250_2150 ();
 b15zdnd11an1n64x5 FILLER_250_2162 ();
 b15zdnd11an1n32x5 FILLER_250_2226 ();
 b15zdnd11an1n16x5 FILLER_250_2258 ();
 b15zdnd00an1n02x5 FILLER_250_2274 ();
 b15zdnd11an1n64x5 FILLER_251_0 ();
 b15zdnd11an1n64x5 FILLER_251_64 ();
 b15zdnd11an1n64x5 FILLER_251_128 ();
 b15zdnd11an1n64x5 FILLER_251_192 ();
 b15zdnd11an1n64x5 FILLER_251_256 ();
 b15zdnd11an1n64x5 FILLER_251_320 ();
 b15zdnd11an1n64x5 FILLER_251_384 ();
 b15zdnd11an1n64x5 FILLER_251_448 ();
 b15zdnd11an1n64x5 FILLER_251_512 ();
 b15zdnd11an1n64x5 FILLER_251_576 ();
 b15zdnd11an1n64x5 FILLER_251_640 ();
 b15zdnd11an1n64x5 FILLER_251_704 ();
 b15zdnd11an1n64x5 FILLER_251_768 ();
 b15zdnd11an1n64x5 FILLER_251_832 ();
 b15zdnd11an1n64x5 FILLER_251_896 ();
 b15zdnd11an1n64x5 FILLER_251_960 ();
 b15zdnd11an1n64x5 FILLER_251_1024 ();
 b15zdnd11an1n64x5 FILLER_251_1088 ();
 b15zdnd11an1n64x5 FILLER_251_1152 ();
 b15zdnd11an1n64x5 FILLER_251_1216 ();
 b15zdnd11an1n64x5 FILLER_251_1280 ();
 b15zdnd11an1n64x5 FILLER_251_1344 ();
 b15zdnd11an1n64x5 FILLER_251_1408 ();
 b15zdnd11an1n64x5 FILLER_251_1472 ();
 b15zdnd11an1n64x5 FILLER_251_1536 ();
 b15zdnd11an1n64x5 FILLER_251_1600 ();
 b15zdnd11an1n64x5 FILLER_251_1664 ();
 b15zdnd11an1n64x5 FILLER_251_1728 ();
 b15zdnd11an1n64x5 FILLER_251_1792 ();
 b15zdnd11an1n64x5 FILLER_251_1856 ();
 b15zdnd11an1n64x5 FILLER_251_1920 ();
 b15zdnd11an1n64x5 FILLER_251_1984 ();
 b15zdnd11an1n32x5 FILLER_251_2048 ();
 b15zdnd11an1n16x5 FILLER_251_2080 ();
 b15zdnd11an1n08x5 FILLER_251_2096 ();
 b15zdnd11an1n04x5 FILLER_251_2104 ();
 b15zdnd11an1n64x5 FILLER_251_2124 ();
 b15zdnd11an1n64x5 FILLER_251_2188 ();
 b15zdnd11an1n32x5 FILLER_251_2252 ();
 b15zdnd11an1n64x5 FILLER_252_8 ();
 b15zdnd11an1n64x5 FILLER_252_72 ();
 b15zdnd11an1n64x5 FILLER_252_136 ();
 b15zdnd11an1n64x5 FILLER_252_200 ();
 b15zdnd11an1n64x5 FILLER_252_264 ();
 b15zdnd11an1n64x5 FILLER_252_328 ();
 b15zdnd11an1n64x5 FILLER_252_392 ();
 b15zdnd11an1n64x5 FILLER_252_456 ();
 b15zdnd11an1n64x5 FILLER_252_520 ();
 b15zdnd11an1n64x5 FILLER_252_584 ();
 b15zdnd11an1n64x5 FILLER_252_648 ();
 b15zdnd11an1n04x5 FILLER_252_712 ();
 b15zdnd00an1n02x5 FILLER_252_716 ();
 b15zdnd11an1n64x5 FILLER_252_726 ();
 b15zdnd11an1n64x5 FILLER_252_790 ();
 b15zdnd11an1n64x5 FILLER_252_854 ();
 b15zdnd11an1n64x5 FILLER_252_918 ();
 b15zdnd11an1n64x5 FILLER_252_982 ();
 b15zdnd11an1n64x5 FILLER_252_1046 ();
 b15zdnd11an1n64x5 FILLER_252_1110 ();
 b15zdnd11an1n64x5 FILLER_252_1174 ();
 b15zdnd11an1n64x5 FILLER_252_1238 ();
 b15zdnd11an1n64x5 FILLER_252_1302 ();
 b15zdnd11an1n64x5 FILLER_252_1366 ();
 b15zdnd11an1n64x5 FILLER_252_1430 ();
 b15zdnd11an1n64x5 FILLER_252_1494 ();
 b15zdnd11an1n64x5 FILLER_252_1558 ();
 b15zdnd11an1n64x5 FILLER_252_1622 ();
 b15zdnd11an1n64x5 FILLER_252_1686 ();
 b15zdnd11an1n64x5 FILLER_252_1750 ();
 b15zdnd11an1n64x5 FILLER_252_1814 ();
 b15zdnd11an1n64x5 FILLER_252_1878 ();
 b15zdnd11an1n64x5 FILLER_252_1942 ();
 b15zdnd11an1n64x5 FILLER_252_2006 ();
 b15zdnd11an1n32x5 FILLER_252_2070 ();
 b15zdnd11an1n08x5 FILLER_252_2102 ();
 b15zdnd00an1n01x5 FILLER_252_2110 ();
 b15zdnd11an1n16x5 FILLER_252_2127 ();
 b15zdnd11an1n08x5 FILLER_252_2143 ();
 b15zdnd00an1n02x5 FILLER_252_2151 ();
 b15zdnd00an1n01x5 FILLER_252_2153 ();
 b15zdnd11an1n64x5 FILLER_252_2162 ();
 b15zdnd11an1n32x5 FILLER_252_2226 ();
 b15zdnd11an1n16x5 FILLER_252_2258 ();
 b15zdnd00an1n02x5 FILLER_252_2274 ();
 b15zdnd11an1n64x5 FILLER_253_0 ();
 b15zdnd11an1n64x5 FILLER_253_64 ();
 b15zdnd11an1n64x5 FILLER_253_128 ();
 b15zdnd11an1n64x5 FILLER_253_192 ();
 b15zdnd11an1n64x5 FILLER_253_256 ();
 b15zdnd11an1n64x5 FILLER_253_320 ();
 b15zdnd11an1n64x5 FILLER_253_384 ();
 b15zdnd11an1n64x5 FILLER_253_448 ();
 b15zdnd11an1n64x5 FILLER_253_512 ();
 b15zdnd11an1n64x5 FILLER_253_576 ();
 b15zdnd11an1n64x5 FILLER_253_640 ();
 b15zdnd11an1n64x5 FILLER_253_704 ();
 b15zdnd11an1n64x5 FILLER_253_768 ();
 b15zdnd11an1n64x5 FILLER_253_832 ();
 b15zdnd11an1n64x5 FILLER_253_896 ();
 b15zdnd11an1n64x5 FILLER_253_960 ();
 b15zdnd11an1n64x5 FILLER_253_1024 ();
 b15zdnd11an1n64x5 FILLER_253_1088 ();
 b15zdnd11an1n64x5 FILLER_253_1152 ();
 b15zdnd11an1n64x5 FILLER_253_1216 ();
 b15zdnd11an1n64x5 FILLER_253_1280 ();
 b15zdnd11an1n64x5 FILLER_253_1344 ();
 b15zdnd11an1n64x5 FILLER_253_1408 ();
 b15zdnd11an1n64x5 FILLER_253_1472 ();
 b15zdnd11an1n64x5 FILLER_253_1536 ();
 b15zdnd11an1n64x5 FILLER_253_1600 ();
 b15zdnd11an1n64x5 FILLER_253_1664 ();
 b15zdnd11an1n64x5 FILLER_253_1728 ();
 b15zdnd11an1n64x5 FILLER_253_1792 ();
 b15zdnd11an1n64x5 FILLER_253_1856 ();
 b15zdnd11an1n64x5 FILLER_253_1920 ();
 b15zdnd11an1n64x5 FILLER_253_1984 ();
 b15zdnd11an1n64x5 FILLER_253_2048 ();
 b15zdnd11an1n64x5 FILLER_253_2112 ();
 b15zdnd11an1n64x5 FILLER_253_2176 ();
 b15zdnd11an1n32x5 FILLER_253_2240 ();
 b15zdnd11an1n08x5 FILLER_253_2272 ();
 b15zdnd11an1n04x5 FILLER_253_2280 ();
 b15zdnd11an1n64x5 FILLER_254_8 ();
 b15zdnd11an1n64x5 FILLER_254_72 ();
 b15zdnd11an1n64x5 FILLER_254_136 ();
 b15zdnd11an1n64x5 FILLER_254_200 ();
 b15zdnd11an1n64x5 FILLER_254_264 ();
 b15zdnd11an1n64x5 FILLER_254_328 ();
 b15zdnd11an1n64x5 FILLER_254_392 ();
 b15zdnd11an1n64x5 FILLER_254_456 ();
 b15zdnd11an1n64x5 FILLER_254_520 ();
 b15zdnd11an1n64x5 FILLER_254_584 ();
 b15zdnd11an1n64x5 FILLER_254_648 ();
 b15zdnd11an1n04x5 FILLER_254_712 ();
 b15zdnd00an1n02x5 FILLER_254_716 ();
 b15zdnd11an1n64x5 FILLER_254_726 ();
 b15zdnd11an1n64x5 FILLER_254_790 ();
 b15zdnd11an1n64x5 FILLER_254_854 ();
 b15zdnd11an1n64x5 FILLER_254_918 ();
 b15zdnd11an1n64x5 FILLER_254_982 ();
 b15zdnd11an1n64x5 FILLER_254_1046 ();
 b15zdnd11an1n64x5 FILLER_254_1110 ();
 b15zdnd11an1n64x5 FILLER_254_1174 ();
 b15zdnd11an1n64x5 FILLER_254_1238 ();
 b15zdnd11an1n64x5 FILLER_254_1302 ();
 b15zdnd11an1n64x5 FILLER_254_1366 ();
 b15zdnd11an1n64x5 FILLER_254_1430 ();
 b15zdnd11an1n64x5 FILLER_254_1494 ();
 b15zdnd11an1n64x5 FILLER_254_1558 ();
 b15zdnd11an1n64x5 FILLER_254_1622 ();
 b15zdnd11an1n64x5 FILLER_254_1686 ();
 b15zdnd11an1n64x5 FILLER_254_1750 ();
 b15zdnd11an1n64x5 FILLER_254_1814 ();
 b15zdnd11an1n64x5 FILLER_254_1878 ();
 b15zdnd11an1n64x5 FILLER_254_1942 ();
 b15zdnd11an1n64x5 FILLER_254_2006 ();
 b15zdnd11an1n64x5 FILLER_254_2070 ();
 b15zdnd11an1n16x5 FILLER_254_2134 ();
 b15zdnd11an1n04x5 FILLER_254_2150 ();
 b15zdnd11an1n64x5 FILLER_254_2162 ();
 b15zdnd11an1n32x5 FILLER_254_2226 ();
 b15zdnd11an1n16x5 FILLER_254_2258 ();
 b15zdnd00an1n02x5 FILLER_254_2274 ();
 b15zdnd11an1n64x5 FILLER_255_0 ();
 b15zdnd11an1n64x5 FILLER_255_64 ();
 b15zdnd11an1n64x5 FILLER_255_128 ();
 b15zdnd11an1n64x5 FILLER_255_192 ();
 b15zdnd11an1n64x5 FILLER_255_256 ();
 b15zdnd11an1n64x5 FILLER_255_320 ();
 b15zdnd11an1n64x5 FILLER_255_384 ();
 b15zdnd11an1n64x5 FILLER_255_448 ();
 b15zdnd11an1n64x5 FILLER_255_512 ();
 b15zdnd11an1n64x5 FILLER_255_576 ();
 b15zdnd11an1n64x5 FILLER_255_640 ();
 b15zdnd11an1n64x5 FILLER_255_704 ();
 b15zdnd11an1n64x5 FILLER_255_768 ();
 b15zdnd11an1n64x5 FILLER_255_832 ();
 b15zdnd11an1n64x5 FILLER_255_896 ();
 b15zdnd11an1n64x5 FILLER_255_960 ();
 b15zdnd11an1n64x5 FILLER_255_1024 ();
 b15zdnd11an1n64x5 FILLER_255_1088 ();
 b15zdnd11an1n64x5 FILLER_255_1152 ();
 b15zdnd11an1n64x5 FILLER_255_1216 ();
 b15zdnd11an1n64x5 FILLER_255_1280 ();
 b15zdnd11an1n64x5 FILLER_255_1344 ();
 b15zdnd11an1n64x5 FILLER_255_1408 ();
 b15zdnd11an1n64x5 FILLER_255_1472 ();
 b15zdnd11an1n64x5 FILLER_255_1536 ();
 b15zdnd11an1n64x5 FILLER_255_1600 ();
 b15zdnd11an1n64x5 FILLER_255_1664 ();
 b15zdnd11an1n64x5 FILLER_255_1728 ();
 b15zdnd11an1n64x5 FILLER_255_1792 ();
 b15zdnd11an1n64x5 FILLER_255_1856 ();
 b15zdnd11an1n64x5 FILLER_255_1920 ();
 b15zdnd11an1n64x5 FILLER_255_1984 ();
 b15zdnd11an1n64x5 FILLER_255_2048 ();
 b15zdnd11an1n64x5 FILLER_255_2112 ();
 b15zdnd11an1n64x5 FILLER_255_2176 ();
 b15zdnd11an1n32x5 FILLER_255_2240 ();
 b15zdnd11an1n08x5 FILLER_255_2272 ();
 b15zdnd11an1n04x5 FILLER_255_2280 ();
 b15zdnd11an1n64x5 FILLER_256_8 ();
 b15zdnd11an1n64x5 FILLER_256_72 ();
 b15zdnd11an1n64x5 FILLER_256_136 ();
 b15zdnd11an1n64x5 FILLER_256_200 ();
 b15zdnd11an1n64x5 FILLER_256_264 ();
 b15zdnd11an1n64x5 FILLER_256_328 ();
 b15zdnd11an1n64x5 FILLER_256_392 ();
 b15zdnd11an1n64x5 FILLER_256_456 ();
 b15zdnd11an1n64x5 FILLER_256_520 ();
 b15zdnd11an1n64x5 FILLER_256_584 ();
 b15zdnd11an1n64x5 FILLER_256_648 ();
 b15zdnd11an1n04x5 FILLER_256_712 ();
 b15zdnd00an1n02x5 FILLER_256_716 ();
 b15zdnd11an1n64x5 FILLER_256_726 ();
 b15zdnd11an1n64x5 FILLER_256_790 ();
 b15zdnd11an1n64x5 FILLER_256_854 ();
 b15zdnd11an1n64x5 FILLER_256_918 ();
 b15zdnd11an1n64x5 FILLER_256_982 ();
 b15zdnd11an1n64x5 FILLER_256_1046 ();
 b15zdnd11an1n64x5 FILLER_256_1110 ();
 b15zdnd11an1n64x5 FILLER_256_1174 ();
 b15zdnd11an1n64x5 FILLER_256_1238 ();
 b15zdnd11an1n64x5 FILLER_256_1302 ();
 b15zdnd11an1n64x5 FILLER_256_1366 ();
 b15zdnd11an1n64x5 FILLER_256_1430 ();
 b15zdnd11an1n64x5 FILLER_256_1494 ();
 b15zdnd11an1n64x5 FILLER_256_1558 ();
 b15zdnd11an1n64x5 FILLER_256_1622 ();
 b15zdnd11an1n64x5 FILLER_256_1686 ();
 b15zdnd11an1n64x5 FILLER_256_1750 ();
 b15zdnd11an1n64x5 FILLER_256_1814 ();
 b15zdnd11an1n64x5 FILLER_256_1878 ();
 b15zdnd11an1n64x5 FILLER_256_1942 ();
 b15zdnd11an1n64x5 FILLER_256_2006 ();
 b15zdnd11an1n64x5 FILLER_256_2070 ();
 b15zdnd11an1n16x5 FILLER_256_2134 ();
 b15zdnd11an1n04x5 FILLER_256_2150 ();
 b15zdnd11an1n64x5 FILLER_256_2162 ();
 b15zdnd11an1n32x5 FILLER_256_2226 ();
 b15zdnd11an1n16x5 FILLER_256_2258 ();
 b15zdnd00an1n02x5 FILLER_256_2274 ();
 b15zdnd11an1n64x5 FILLER_257_0 ();
 b15zdnd11an1n64x5 FILLER_257_64 ();
 b15zdnd11an1n64x5 FILLER_257_128 ();
 b15zdnd11an1n64x5 FILLER_257_192 ();
 b15zdnd11an1n64x5 FILLER_257_256 ();
 b15zdnd11an1n64x5 FILLER_257_320 ();
 b15zdnd11an1n64x5 FILLER_257_384 ();
 b15zdnd11an1n64x5 FILLER_257_448 ();
 b15zdnd11an1n64x5 FILLER_257_512 ();
 b15zdnd11an1n64x5 FILLER_257_576 ();
 b15zdnd11an1n64x5 FILLER_257_640 ();
 b15zdnd11an1n64x5 FILLER_257_704 ();
 b15zdnd11an1n64x5 FILLER_257_768 ();
 b15zdnd11an1n64x5 FILLER_257_832 ();
 b15zdnd11an1n64x5 FILLER_257_896 ();
 b15zdnd11an1n64x5 FILLER_257_960 ();
 b15zdnd11an1n64x5 FILLER_257_1024 ();
 b15zdnd11an1n64x5 FILLER_257_1088 ();
 b15zdnd11an1n64x5 FILLER_257_1152 ();
 b15zdnd11an1n64x5 FILLER_257_1216 ();
 b15zdnd11an1n64x5 FILLER_257_1280 ();
 b15zdnd11an1n64x5 FILLER_257_1344 ();
 b15zdnd11an1n64x5 FILLER_257_1408 ();
 b15zdnd11an1n64x5 FILLER_257_1472 ();
 b15zdnd11an1n64x5 FILLER_257_1536 ();
 b15zdnd11an1n64x5 FILLER_257_1600 ();
 b15zdnd11an1n64x5 FILLER_257_1664 ();
 b15zdnd11an1n64x5 FILLER_257_1728 ();
 b15zdnd11an1n64x5 FILLER_257_1792 ();
 b15zdnd11an1n64x5 FILLER_257_1856 ();
 b15zdnd11an1n64x5 FILLER_257_1920 ();
 b15zdnd11an1n64x5 FILLER_257_1984 ();
 b15zdnd11an1n64x5 FILLER_257_2048 ();
 b15zdnd11an1n64x5 FILLER_257_2112 ();
 b15zdnd11an1n64x5 FILLER_257_2176 ();
 b15zdnd11an1n32x5 FILLER_257_2240 ();
 b15zdnd11an1n08x5 FILLER_257_2272 ();
 b15zdnd11an1n04x5 FILLER_257_2280 ();
 b15zdnd11an1n64x5 FILLER_258_8 ();
 b15zdnd11an1n64x5 FILLER_258_72 ();
 b15zdnd11an1n64x5 FILLER_258_136 ();
 b15zdnd11an1n64x5 FILLER_258_200 ();
 b15zdnd11an1n64x5 FILLER_258_264 ();
 b15zdnd11an1n64x5 FILLER_258_328 ();
 b15zdnd11an1n64x5 FILLER_258_392 ();
 b15zdnd11an1n64x5 FILLER_258_456 ();
 b15zdnd11an1n64x5 FILLER_258_520 ();
 b15zdnd11an1n64x5 FILLER_258_584 ();
 b15zdnd11an1n64x5 FILLER_258_648 ();
 b15zdnd11an1n04x5 FILLER_258_712 ();
 b15zdnd00an1n02x5 FILLER_258_716 ();
 b15zdnd11an1n64x5 FILLER_258_726 ();
 b15zdnd11an1n64x5 FILLER_258_790 ();
 b15zdnd11an1n64x5 FILLER_258_854 ();
 b15zdnd11an1n64x5 FILLER_258_918 ();
 b15zdnd11an1n64x5 FILLER_258_982 ();
 b15zdnd11an1n64x5 FILLER_258_1046 ();
 b15zdnd11an1n64x5 FILLER_258_1110 ();
 b15zdnd11an1n64x5 FILLER_258_1174 ();
 b15zdnd11an1n64x5 FILLER_258_1238 ();
 b15zdnd11an1n64x5 FILLER_258_1302 ();
 b15zdnd11an1n64x5 FILLER_258_1366 ();
 b15zdnd11an1n64x5 FILLER_258_1430 ();
 b15zdnd11an1n64x5 FILLER_258_1494 ();
 b15zdnd11an1n64x5 FILLER_258_1558 ();
 b15zdnd11an1n64x5 FILLER_258_1622 ();
 b15zdnd11an1n64x5 FILLER_258_1686 ();
 b15zdnd11an1n64x5 FILLER_258_1750 ();
 b15zdnd11an1n64x5 FILLER_258_1814 ();
 b15zdnd11an1n64x5 FILLER_258_1878 ();
 b15zdnd11an1n64x5 FILLER_258_1942 ();
 b15zdnd11an1n64x5 FILLER_258_2006 ();
 b15zdnd11an1n64x5 FILLER_258_2070 ();
 b15zdnd11an1n16x5 FILLER_258_2134 ();
 b15zdnd11an1n04x5 FILLER_258_2150 ();
 b15zdnd11an1n64x5 FILLER_258_2162 ();
 b15zdnd11an1n32x5 FILLER_258_2226 ();
 b15zdnd11an1n16x5 FILLER_258_2258 ();
 b15zdnd00an1n02x5 FILLER_258_2274 ();
 b15zdnd11an1n64x5 FILLER_259_0 ();
 b15zdnd11an1n64x5 FILLER_259_64 ();
 b15zdnd11an1n64x5 FILLER_259_128 ();
 b15zdnd11an1n64x5 FILLER_259_192 ();
 b15zdnd11an1n64x5 FILLER_259_256 ();
 b15zdnd11an1n64x5 FILLER_259_320 ();
 b15zdnd11an1n64x5 FILLER_259_384 ();
 b15zdnd11an1n64x5 FILLER_259_448 ();
 b15zdnd11an1n64x5 FILLER_259_512 ();
 b15zdnd11an1n64x5 FILLER_259_576 ();
 b15zdnd11an1n64x5 FILLER_259_640 ();
 b15zdnd11an1n64x5 FILLER_259_704 ();
 b15zdnd11an1n64x5 FILLER_259_768 ();
 b15zdnd11an1n64x5 FILLER_259_832 ();
 b15zdnd11an1n64x5 FILLER_259_896 ();
 b15zdnd11an1n64x5 FILLER_259_960 ();
 b15zdnd11an1n64x5 FILLER_259_1024 ();
 b15zdnd11an1n64x5 FILLER_259_1088 ();
 b15zdnd11an1n64x5 FILLER_259_1152 ();
 b15zdnd11an1n64x5 FILLER_259_1216 ();
 b15zdnd11an1n64x5 FILLER_259_1280 ();
 b15zdnd11an1n64x5 FILLER_259_1344 ();
 b15zdnd11an1n64x5 FILLER_259_1408 ();
 b15zdnd11an1n64x5 FILLER_259_1472 ();
 b15zdnd11an1n64x5 FILLER_259_1536 ();
 b15zdnd11an1n64x5 FILLER_259_1600 ();
 b15zdnd11an1n64x5 FILLER_259_1664 ();
 b15zdnd11an1n64x5 FILLER_259_1728 ();
 b15zdnd11an1n64x5 FILLER_259_1792 ();
 b15zdnd11an1n64x5 FILLER_259_1856 ();
 b15zdnd11an1n64x5 FILLER_259_1920 ();
 b15zdnd11an1n64x5 FILLER_259_1984 ();
 b15zdnd11an1n64x5 FILLER_259_2048 ();
 b15zdnd11an1n64x5 FILLER_259_2112 ();
 b15zdnd11an1n64x5 FILLER_259_2176 ();
 b15zdnd11an1n32x5 FILLER_259_2240 ();
 b15zdnd11an1n08x5 FILLER_259_2272 ();
 b15zdnd11an1n04x5 FILLER_259_2280 ();
 b15zdnd11an1n64x5 FILLER_260_8 ();
 b15zdnd11an1n64x5 FILLER_260_72 ();
 b15zdnd11an1n64x5 FILLER_260_136 ();
 b15zdnd11an1n64x5 FILLER_260_200 ();
 b15zdnd11an1n64x5 FILLER_260_264 ();
 b15zdnd11an1n64x5 FILLER_260_328 ();
 b15zdnd11an1n64x5 FILLER_260_392 ();
 b15zdnd11an1n64x5 FILLER_260_456 ();
 b15zdnd11an1n64x5 FILLER_260_520 ();
 b15zdnd11an1n64x5 FILLER_260_584 ();
 b15zdnd11an1n64x5 FILLER_260_648 ();
 b15zdnd11an1n04x5 FILLER_260_712 ();
 b15zdnd00an1n02x5 FILLER_260_716 ();
 b15zdnd11an1n64x5 FILLER_260_726 ();
 b15zdnd11an1n64x5 FILLER_260_790 ();
 b15zdnd11an1n64x5 FILLER_260_854 ();
 b15zdnd11an1n64x5 FILLER_260_918 ();
 b15zdnd11an1n64x5 FILLER_260_982 ();
 b15zdnd11an1n64x5 FILLER_260_1046 ();
 b15zdnd11an1n64x5 FILLER_260_1110 ();
 b15zdnd11an1n64x5 FILLER_260_1174 ();
 b15zdnd11an1n64x5 FILLER_260_1238 ();
 b15zdnd11an1n64x5 FILLER_260_1302 ();
 b15zdnd11an1n64x5 FILLER_260_1366 ();
 b15zdnd11an1n64x5 FILLER_260_1430 ();
 b15zdnd11an1n64x5 FILLER_260_1494 ();
 b15zdnd11an1n64x5 FILLER_260_1558 ();
 b15zdnd11an1n64x5 FILLER_260_1622 ();
 b15zdnd11an1n64x5 FILLER_260_1686 ();
 b15zdnd11an1n64x5 FILLER_260_1750 ();
 b15zdnd11an1n64x5 FILLER_260_1814 ();
 b15zdnd11an1n64x5 FILLER_260_1878 ();
 b15zdnd11an1n64x5 FILLER_260_1942 ();
 b15zdnd11an1n64x5 FILLER_260_2006 ();
 b15zdnd11an1n64x5 FILLER_260_2070 ();
 b15zdnd11an1n16x5 FILLER_260_2134 ();
 b15zdnd11an1n04x5 FILLER_260_2150 ();
 b15zdnd11an1n64x5 FILLER_260_2162 ();
 b15zdnd11an1n32x5 FILLER_260_2226 ();
 b15zdnd11an1n16x5 FILLER_260_2258 ();
 b15zdnd00an1n02x5 FILLER_260_2274 ();
 b15zdnd11an1n64x5 FILLER_261_0 ();
 b15zdnd11an1n64x5 FILLER_261_64 ();
 b15zdnd11an1n64x5 FILLER_261_128 ();
 b15zdnd11an1n64x5 FILLER_261_192 ();
 b15zdnd11an1n64x5 FILLER_261_256 ();
 b15zdnd11an1n64x5 FILLER_261_320 ();
 b15zdnd11an1n64x5 FILLER_261_384 ();
 b15zdnd11an1n64x5 FILLER_261_448 ();
 b15zdnd11an1n64x5 FILLER_261_512 ();
 b15zdnd11an1n64x5 FILLER_261_576 ();
 b15zdnd11an1n64x5 FILLER_261_640 ();
 b15zdnd11an1n64x5 FILLER_261_704 ();
 b15zdnd11an1n64x5 FILLER_261_768 ();
 b15zdnd11an1n64x5 FILLER_261_832 ();
 b15zdnd11an1n64x5 FILLER_261_896 ();
 b15zdnd11an1n64x5 FILLER_261_960 ();
 b15zdnd11an1n64x5 FILLER_261_1024 ();
 b15zdnd11an1n64x5 FILLER_261_1088 ();
 b15zdnd11an1n64x5 FILLER_261_1152 ();
 b15zdnd11an1n64x5 FILLER_261_1216 ();
 b15zdnd11an1n64x5 FILLER_261_1280 ();
 b15zdnd11an1n64x5 FILLER_261_1344 ();
 b15zdnd11an1n64x5 FILLER_261_1408 ();
 b15zdnd11an1n64x5 FILLER_261_1472 ();
 b15zdnd11an1n64x5 FILLER_261_1536 ();
 b15zdnd11an1n64x5 FILLER_261_1600 ();
 b15zdnd11an1n64x5 FILLER_261_1664 ();
 b15zdnd11an1n64x5 FILLER_261_1728 ();
 b15zdnd11an1n64x5 FILLER_261_1792 ();
 b15zdnd11an1n64x5 FILLER_261_1856 ();
 b15zdnd11an1n64x5 FILLER_261_1920 ();
 b15zdnd11an1n64x5 FILLER_261_1984 ();
 b15zdnd11an1n64x5 FILLER_261_2048 ();
 b15zdnd11an1n64x5 FILLER_261_2112 ();
 b15zdnd11an1n64x5 FILLER_261_2176 ();
 b15zdnd11an1n32x5 FILLER_261_2240 ();
 b15zdnd11an1n08x5 FILLER_261_2272 ();
 b15zdnd11an1n04x5 FILLER_261_2280 ();
 b15zdnd11an1n64x5 FILLER_262_8 ();
 b15zdnd11an1n64x5 FILLER_262_72 ();
 b15zdnd11an1n64x5 FILLER_262_136 ();
 b15zdnd11an1n64x5 FILLER_262_200 ();
 b15zdnd11an1n64x5 FILLER_262_264 ();
 b15zdnd11an1n64x5 FILLER_262_328 ();
 b15zdnd11an1n64x5 FILLER_262_392 ();
 b15zdnd11an1n64x5 FILLER_262_456 ();
 b15zdnd11an1n64x5 FILLER_262_520 ();
 b15zdnd11an1n64x5 FILLER_262_584 ();
 b15zdnd11an1n64x5 FILLER_262_648 ();
 b15zdnd11an1n04x5 FILLER_262_712 ();
 b15zdnd00an1n02x5 FILLER_262_716 ();
 b15zdnd11an1n64x5 FILLER_262_726 ();
 b15zdnd11an1n64x5 FILLER_262_790 ();
 b15zdnd11an1n64x5 FILLER_262_854 ();
 b15zdnd11an1n64x5 FILLER_262_918 ();
 b15zdnd11an1n64x5 FILLER_262_982 ();
 b15zdnd11an1n64x5 FILLER_262_1046 ();
 b15zdnd11an1n64x5 FILLER_262_1110 ();
 b15zdnd11an1n64x5 FILLER_262_1174 ();
 b15zdnd11an1n64x5 FILLER_262_1238 ();
 b15zdnd11an1n64x5 FILLER_262_1302 ();
 b15zdnd11an1n64x5 FILLER_262_1366 ();
 b15zdnd11an1n64x5 FILLER_262_1430 ();
 b15zdnd11an1n64x5 FILLER_262_1494 ();
 b15zdnd11an1n64x5 FILLER_262_1558 ();
 b15zdnd11an1n64x5 FILLER_262_1622 ();
 b15zdnd11an1n64x5 FILLER_262_1686 ();
 b15zdnd11an1n64x5 FILLER_262_1750 ();
 b15zdnd11an1n64x5 FILLER_262_1814 ();
 b15zdnd11an1n64x5 FILLER_262_1878 ();
 b15zdnd11an1n64x5 FILLER_262_1942 ();
 b15zdnd11an1n64x5 FILLER_262_2006 ();
 b15zdnd11an1n64x5 FILLER_262_2070 ();
 b15zdnd11an1n16x5 FILLER_262_2134 ();
 b15zdnd11an1n04x5 FILLER_262_2150 ();
 b15zdnd11an1n64x5 FILLER_262_2162 ();
 b15zdnd11an1n32x5 FILLER_262_2226 ();
 b15zdnd11an1n16x5 FILLER_262_2258 ();
 b15zdnd00an1n02x5 FILLER_262_2274 ();
 b15zdnd11an1n64x5 FILLER_263_0 ();
 b15zdnd11an1n64x5 FILLER_263_64 ();
 b15zdnd11an1n64x5 FILLER_263_128 ();
 b15zdnd11an1n64x5 FILLER_263_192 ();
 b15zdnd11an1n64x5 FILLER_263_256 ();
 b15zdnd11an1n64x5 FILLER_263_320 ();
 b15zdnd11an1n64x5 FILLER_263_384 ();
 b15zdnd11an1n64x5 FILLER_263_448 ();
 b15zdnd11an1n64x5 FILLER_263_512 ();
 b15zdnd11an1n64x5 FILLER_263_576 ();
 b15zdnd11an1n64x5 FILLER_263_640 ();
 b15zdnd11an1n64x5 FILLER_263_704 ();
 b15zdnd11an1n64x5 FILLER_263_768 ();
 b15zdnd11an1n64x5 FILLER_263_832 ();
 b15zdnd11an1n64x5 FILLER_263_896 ();
 b15zdnd11an1n64x5 FILLER_263_960 ();
 b15zdnd11an1n64x5 FILLER_263_1024 ();
 b15zdnd11an1n64x5 FILLER_263_1088 ();
 b15zdnd11an1n64x5 FILLER_263_1152 ();
 b15zdnd11an1n64x5 FILLER_263_1216 ();
 b15zdnd11an1n64x5 FILLER_263_1280 ();
 b15zdnd11an1n64x5 FILLER_263_1344 ();
 b15zdnd11an1n64x5 FILLER_263_1408 ();
 b15zdnd11an1n64x5 FILLER_263_1472 ();
 b15zdnd11an1n64x5 FILLER_263_1536 ();
 b15zdnd11an1n64x5 FILLER_263_1600 ();
 b15zdnd11an1n64x5 FILLER_263_1664 ();
 b15zdnd11an1n64x5 FILLER_263_1728 ();
 b15zdnd11an1n64x5 FILLER_263_1792 ();
 b15zdnd11an1n64x5 FILLER_263_1856 ();
 b15zdnd11an1n64x5 FILLER_263_1920 ();
 b15zdnd11an1n64x5 FILLER_263_1984 ();
 b15zdnd11an1n64x5 FILLER_263_2048 ();
 b15zdnd11an1n64x5 FILLER_263_2112 ();
 b15zdnd11an1n64x5 FILLER_263_2176 ();
 b15zdnd11an1n32x5 FILLER_263_2240 ();
 b15zdnd11an1n08x5 FILLER_263_2272 ();
 b15zdnd11an1n04x5 FILLER_263_2280 ();
 b15zdnd11an1n64x5 FILLER_264_8 ();
 b15zdnd11an1n64x5 FILLER_264_72 ();
 b15zdnd11an1n64x5 FILLER_264_136 ();
 b15zdnd11an1n64x5 FILLER_264_200 ();
 b15zdnd11an1n64x5 FILLER_264_264 ();
 b15zdnd11an1n64x5 FILLER_264_328 ();
 b15zdnd11an1n64x5 FILLER_264_392 ();
 b15zdnd11an1n64x5 FILLER_264_456 ();
 b15zdnd11an1n64x5 FILLER_264_520 ();
 b15zdnd11an1n64x5 FILLER_264_584 ();
 b15zdnd11an1n64x5 FILLER_264_648 ();
 b15zdnd11an1n04x5 FILLER_264_712 ();
 b15zdnd00an1n02x5 FILLER_264_716 ();
 b15zdnd11an1n64x5 FILLER_264_726 ();
 b15zdnd11an1n64x5 FILLER_264_790 ();
 b15zdnd11an1n64x5 FILLER_264_854 ();
 b15zdnd11an1n64x5 FILLER_264_918 ();
 b15zdnd11an1n64x5 FILLER_264_982 ();
 b15zdnd11an1n64x5 FILLER_264_1046 ();
 b15zdnd11an1n64x5 FILLER_264_1110 ();
 b15zdnd11an1n64x5 FILLER_264_1174 ();
 b15zdnd11an1n64x5 FILLER_264_1238 ();
 b15zdnd11an1n64x5 FILLER_264_1302 ();
 b15zdnd11an1n64x5 FILLER_264_1366 ();
 b15zdnd11an1n64x5 FILLER_264_1430 ();
 b15zdnd11an1n64x5 FILLER_264_1494 ();
 b15zdnd11an1n64x5 FILLER_264_1558 ();
 b15zdnd11an1n64x5 FILLER_264_1622 ();
 b15zdnd11an1n64x5 FILLER_264_1686 ();
 b15zdnd11an1n64x5 FILLER_264_1750 ();
 b15zdnd11an1n64x5 FILLER_264_1814 ();
 b15zdnd11an1n64x5 FILLER_264_1878 ();
 b15zdnd11an1n64x5 FILLER_264_1942 ();
 b15zdnd11an1n64x5 FILLER_264_2006 ();
 b15zdnd11an1n64x5 FILLER_264_2070 ();
 b15zdnd11an1n16x5 FILLER_264_2134 ();
 b15zdnd11an1n04x5 FILLER_264_2150 ();
 b15zdnd11an1n64x5 FILLER_264_2162 ();
 b15zdnd11an1n32x5 FILLER_264_2226 ();
 b15zdnd11an1n16x5 FILLER_264_2258 ();
 b15zdnd00an1n02x5 FILLER_264_2274 ();
 b15zdnd11an1n64x5 FILLER_265_0 ();
 b15zdnd11an1n64x5 FILLER_265_64 ();
 b15zdnd11an1n64x5 FILLER_265_128 ();
 b15zdnd11an1n64x5 FILLER_265_192 ();
 b15zdnd11an1n64x5 FILLER_265_256 ();
 b15zdnd11an1n64x5 FILLER_265_320 ();
 b15zdnd11an1n64x5 FILLER_265_384 ();
 b15zdnd11an1n64x5 FILLER_265_448 ();
 b15zdnd11an1n64x5 FILLER_265_512 ();
 b15zdnd11an1n64x5 FILLER_265_576 ();
 b15zdnd11an1n64x5 FILLER_265_640 ();
 b15zdnd11an1n64x5 FILLER_265_704 ();
 b15zdnd11an1n64x5 FILLER_265_768 ();
 b15zdnd11an1n64x5 FILLER_265_832 ();
 b15zdnd11an1n64x5 FILLER_265_896 ();
 b15zdnd11an1n64x5 FILLER_265_960 ();
 b15zdnd11an1n64x5 FILLER_265_1024 ();
 b15zdnd11an1n64x5 FILLER_265_1088 ();
 b15zdnd11an1n64x5 FILLER_265_1152 ();
 b15zdnd11an1n64x5 FILLER_265_1216 ();
 b15zdnd11an1n64x5 FILLER_265_1280 ();
 b15zdnd11an1n64x5 FILLER_265_1344 ();
 b15zdnd11an1n64x5 FILLER_265_1408 ();
 b15zdnd11an1n64x5 FILLER_265_1472 ();
 b15zdnd11an1n64x5 FILLER_265_1536 ();
 b15zdnd11an1n64x5 FILLER_265_1600 ();
 b15zdnd11an1n64x5 FILLER_265_1664 ();
 b15zdnd11an1n64x5 FILLER_265_1728 ();
 b15zdnd11an1n64x5 FILLER_265_1792 ();
 b15zdnd11an1n64x5 FILLER_265_1856 ();
 b15zdnd11an1n64x5 FILLER_265_1920 ();
 b15zdnd11an1n64x5 FILLER_265_1984 ();
 b15zdnd11an1n64x5 FILLER_265_2048 ();
 b15zdnd11an1n64x5 FILLER_265_2112 ();
 b15zdnd11an1n64x5 FILLER_265_2176 ();
 b15zdnd11an1n32x5 FILLER_265_2240 ();
 b15zdnd11an1n08x5 FILLER_265_2272 ();
 b15zdnd11an1n04x5 FILLER_265_2280 ();
 b15zdnd11an1n64x5 FILLER_266_8 ();
 b15zdnd11an1n64x5 FILLER_266_72 ();
 b15zdnd11an1n64x5 FILLER_266_136 ();
 b15zdnd11an1n64x5 FILLER_266_200 ();
 b15zdnd11an1n64x5 FILLER_266_264 ();
 b15zdnd11an1n64x5 FILLER_266_328 ();
 b15zdnd11an1n64x5 FILLER_266_392 ();
 b15zdnd11an1n64x5 FILLER_266_456 ();
 b15zdnd11an1n64x5 FILLER_266_520 ();
 b15zdnd11an1n64x5 FILLER_266_584 ();
 b15zdnd11an1n64x5 FILLER_266_648 ();
 b15zdnd11an1n04x5 FILLER_266_712 ();
 b15zdnd00an1n02x5 FILLER_266_716 ();
 b15zdnd11an1n64x5 FILLER_266_726 ();
 b15zdnd11an1n64x5 FILLER_266_790 ();
 b15zdnd11an1n64x5 FILLER_266_854 ();
 b15zdnd11an1n64x5 FILLER_266_918 ();
 b15zdnd11an1n64x5 FILLER_266_982 ();
 b15zdnd11an1n64x5 FILLER_266_1046 ();
 b15zdnd11an1n64x5 FILLER_266_1110 ();
 b15zdnd11an1n64x5 FILLER_266_1174 ();
 b15zdnd11an1n64x5 FILLER_266_1238 ();
 b15zdnd11an1n64x5 FILLER_266_1302 ();
 b15zdnd11an1n64x5 FILLER_266_1366 ();
 b15zdnd11an1n64x5 FILLER_266_1430 ();
 b15zdnd11an1n64x5 FILLER_266_1494 ();
 b15zdnd11an1n64x5 FILLER_266_1558 ();
 b15zdnd11an1n64x5 FILLER_266_1622 ();
 b15zdnd11an1n64x5 FILLER_266_1686 ();
 b15zdnd11an1n64x5 FILLER_266_1750 ();
 b15zdnd11an1n64x5 FILLER_266_1814 ();
 b15zdnd11an1n64x5 FILLER_266_1878 ();
 b15zdnd11an1n64x5 FILLER_266_1942 ();
 b15zdnd11an1n64x5 FILLER_266_2006 ();
 b15zdnd11an1n64x5 FILLER_266_2070 ();
 b15zdnd11an1n16x5 FILLER_266_2134 ();
 b15zdnd11an1n04x5 FILLER_266_2150 ();
 b15zdnd11an1n64x5 FILLER_266_2162 ();
 b15zdnd11an1n32x5 FILLER_266_2226 ();
 b15zdnd11an1n16x5 FILLER_266_2258 ();
 b15zdnd00an1n02x5 FILLER_266_2274 ();
 b15zdnd11an1n64x5 FILLER_267_0 ();
 b15zdnd11an1n64x5 FILLER_267_64 ();
 b15zdnd11an1n64x5 FILLER_267_128 ();
 b15zdnd11an1n64x5 FILLER_267_192 ();
 b15zdnd11an1n64x5 FILLER_267_256 ();
 b15zdnd11an1n64x5 FILLER_267_320 ();
 b15zdnd11an1n64x5 FILLER_267_384 ();
 b15zdnd11an1n64x5 FILLER_267_448 ();
 b15zdnd11an1n64x5 FILLER_267_512 ();
 b15zdnd11an1n64x5 FILLER_267_576 ();
 b15zdnd11an1n64x5 FILLER_267_640 ();
 b15zdnd11an1n64x5 FILLER_267_704 ();
 b15zdnd11an1n64x5 FILLER_267_768 ();
 b15zdnd11an1n64x5 FILLER_267_832 ();
 b15zdnd11an1n64x5 FILLER_267_896 ();
 b15zdnd11an1n64x5 FILLER_267_960 ();
 b15zdnd11an1n64x5 FILLER_267_1024 ();
 b15zdnd11an1n64x5 FILLER_267_1088 ();
 b15zdnd11an1n64x5 FILLER_267_1152 ();
 b15zdnd11an1n64x5 FILLER_267_1216 ();
 b15zdnd11an1n64x5 FILLER_267_1280 ();
 b15zdnd11an1n64x5 FILLER_267_1344 ();
 b15zdnd11an1n64x5 FILLER_267_1408 ();
 b15zdnd11an1n64x5 FILLER_267_1472 ();
 b15zdnd11an1n64x5 FILLER_267_1536 ();
 b15zdnd11an1n64x5 FILLER_267_1600 ();
 b15zdnd11an1n64x5 FILLER_267_1664 ();
 b15zdnd11an1n64x5 FILLER_267_1728 ();
 b15zdnd11an1n64x5 FILLER_267_1792 ();
 b15zdnd11an1n64x5 FILLER_267_1856 ();
 b15zdnd11an1n64x5 FILLER_267_1920 ();
 b15zdnd11an1n64x5 FILLER_267_1984 ();
 b15zdnd11an1n64x5 FILLER_267_2048 ();
 b15zdnd11an1n64x5 FILLER_267_2112 ();
 b15zdnd11an1n64x5 FILLER_267_2176 ();
 b15zdnd11an1n32x5 FILLER_267_2240 ();
 b15zdnd11an1n08x5 FILLER_267_2272 ();
 b15zdnd11an1n04x5 FILLER_267_2280 ();
 b15zdnd11an1n64x5 FILLER_268_8 ();
 b15zdnd11an1n64x5 FILLER_268_72 ();
 b15zdnd11an1n64x5 FILLER_268_136 ();
 b15zdnd11an1n64x5 FILLER_268_200 ();
 b15zdnd11an1n64x5 FILLER_268_264 ();
 b15zdnd11an1n64x5 FILLER_268_328 ();
 b15zdnd11an1n64x5 FILLER_268_392 ();
 b15zdnd11an1n64x5 FILLER_268_456 ();
 b15zdnd11an1n64x5 FILLER_268_520 ();
 b15zdnd11an1n64x5 FILLER_268_584 ();
 b15zdnd11an1n64x5 FILLER_268_648 ();
 b15zdnd11an1n04x5 FILLER_268_712 ();
 b15zdnd00an1n02x5 FILLER_268_716 ();
 b15zdnd11an1n64x5 FILLER_268_726 ();
 b15zdnd11an1n64x5 FILLER_268_790 ();
 b15zdnd11an1n64x5 FILLER_268_854 ();
 b15zdnd11an1n64x5 FILLER_268_918 ();
 b15zdnd11an1n64x5 FILLER_268_982 ();
 b15zdnd11an1n64x5 FILLER_268_1046 ();
 b15zdnd11an1n64x5 FILLER_268_1110 ();
 b15zdnd11an1n64x5 FILLER_268_1174 ();
 b15zdnd11an1n64x5 FILLER_268_1238 ();
 b15zdnd11an1n64x5 FILLER_268_1302 ();
 b15zdnd11an1n64x5 FILLER_268_1366 ();
 b15zdnd11an1n64x5 FILLER_268_1430 ();
 b15zdnd11an1n64x5 FILLER_268_1494 ();
 b15zdnd11an1n64x5 FILLER_268_1558 ();
 b15zdnd11an1n64x5 FILLER_268_1622 ();
 b15zdnd11an1n64x5 FILLER_268_1686 ();
 b15zdnd11an1n64x5 FILLER_268_1750 ();
 b15zdnd11an1n64x5 FILLER_268_1814 ();
 b15zdnd11an1n64x5 FILLER_268_1878 ();
 b15zdnd11an1n64x5 FILLER_268_1942 ();
 b15zdnd11an1n64x5 FILLER_268_2006 ();
 b15zdnd11an1n64x5 FILLER_268_2070 ();
 b15zdnd11an1n16x5 FILLER_268_2134 ();
 b15zdnd11an1n04x5 FILLER_268_2150 ();
 b15zdnd11an1n64x5 FILLER_268_2162 ();
 b15zdnd11an1n32x5 FILLER_268_2226 ();
 b15zdnd11an1n16x5 FILLER_268_2258 ();
 b15zdnd00an1n02x5 FILLER_268_2274 ();
 b15zdnd11an1n64x5 FILLER_269_0 ();
 b15zdnd11an1n64x5 FILLER_269_64 ();
 b15zdnd11an1n64x5 FILLER_269_128 ();
 b15zdnd11an1n64x5 FILLER_269_192 ();
 b15zdnd11an1n64x5 FILLER_269_256 ();
 b15zdnd11an1n64x5 FILLER_269_320 ();
 b15zdnd11an1n64x5 FILLER_269_384 ();
 b15zdnd11an1n64x5 FILLER_269_448 ();
 b15zdnd11an1n64x5 FILLER_269_512 ();
 b15zdnd11an1n64x5 FILLER_269_576 ();
 b15zdnd11an1n64x5 FILLER_269_640 ();
 b15zdnd11an1n64x5 FILLER_269_704 ();
 b15zdnd11an1n64x5 FILLER_269_768 ();
 b15zdnd11an1n64x5 FILLER_269_832 ();
 b15zdnd11an1n64x5 FILLER_269_896 ();
 b15zdnd11an1n64x5 FILLER_269_960 ();
 b15zdnd11an1n64x5 FILLER_269_1024 ();
 b15zdnd11an1n64x5 FILLER_269_1088 ();
 b15zdnd11an1n64x5 FILLER_269_1152 ();
 b15zdnd11an1n64x5 FILLER_269_1216 ();
 b15zdnd11an1n64x5 FILLER_269_1280 ();
 b15zdnd11an1n64x5 FILLER_269_1344 ();
 b15zdnd11an1n64x5 FILLER_269_1408 ();
 b15zdnd11an1n64x5 FILLER_269_1472 ();
 b15zdnd11an1n64x5 FILLER_269_1536 ();
 b15zdnd11an1n64x5 FILLER_269_1600 ();
 b15zdnd11an1n64x5 FILLER_269_1664 ();
 b15zdnd11an1n64x5 FILLER_269_1728 ();
 b15zdnd11an1n64x5 FILLER_269_1792 ();
 b15zdnd11an1n64x5 FILLER_269_1856 ();
 b15zdnd11an1n64x5 FILLER_269_1920 ();
 b15zdnd11an1n64x5 FILLER_269_1984 ();
 b15zdnd11an1n64x5 FILLER_269_2048 ();
 b15zdnd11an1n64x5 FILLER_269_2112 ();
 b15zdnd11an1n64x5 FILLER_269_2176 ();
 b15zdnd11an1n32x5 FILLER_269_2240 ();
 b15zdnd11an1n08x5 FILLER_269_2272 ();
 b15zdnd11an1n04x5 FILLER_269_2280 ();
 b15zdnd11an1n64x5 FILLER_270_8 ();
 b15zdnd11an1n64x5 FILLER_270_72 ();
 b15zdnd11an1n64x5 FILLER_270_136 ();
 b15zdnd11an1n64x5 FILLER_270_200 ();
 b15zdnd11an1n64x5 FILLER_270_264 ();
 b15zdnd11an1n64x5 FILLER_270_328 ();
 b15zdnd11an1n64x5 FILLER_270_392 ();
 b15zdnd11an1n64x5 FILLER_270_456 ();
 b15zdnd11an1n64x5 FILLER_270_520 ();
 b15zdnd11an1n64x5 FILLER_270_584 ();
 b15zdnd11an1n64x5 FILLER_270_648 ();
 b15zdnd11an1n04x5 FILLER_270_712 ();
 b15zdnd00an1n02x5 FILLER_270_716 ();
 b15zdnd11an1n64x5 FILLER_270_726 ();
 b15zdnd11an1n64x5 FILLER_270_790 ();
 b15zdnd11an1n64x5 FILLER_270_854 ();
 b15zdnd11an1n64x5 FILLER_270_918 ();
 b15zdnd11an1n64x5 FILLER_270_982 ();
 b15zdnd11an1n64x5 FILLER_270_1046 ();
 b15zdnd11an1n64x5 FILLER_270_1110 ();
 b15zdnd11an1n64x5 FILLER_270_1174 ();
 b15zdnd11an1n64x5 FILLER_270_1238 ();
 b15zdnd11an1n64x5 FILLER_270_1302 ();
 b15zdnd11an1n64x5 FILLER_270_1366 ();
 b15zdnd11an1n64x5 FILLER_270_1430 ();
 b15zdnd11an1n64x5 FILLER_270_1494 ();
 b15zdnd11an1n64x5 FILLER_270_1558 ();
 b15zdnd11an1n64x5 FILLER_270_1622 ();
 b15zdnd11an1n64x5 FILLER_270_1686 ();
 b15zdnd11an1n64x5 FILLER_270_1750 ();
 b15zdnd11an1n64x5 FILLER_270_1814 ();
 b15zdnd11an1n64x5 FILLER_270_1878 ();
 b15zdnd11an1n64x5 FILLER_270_1942 ();
 b15zdnd11an1n64x5 FILLER_270_2006 ();
 b15zdnd11an1n64x5 FILLER_270_2070 ();
 b15zdnd11an1n16x5 FILLER_270_2134 ();
 b15zdnd11an1n04x5 FILLER_270_2150 ();
 b15zdnd11an1n64x5 FILLER_270_2162 ();
 b15zdnd11an1n32x5 FILLER_270_2226 ();
 b15zdnd11an1n16x5 FILLER_270_2258 ();
 b15zdnd00an1n02x5 FILLER_270_2274 ();
 b15zdnd11an1n64x5 FILLER_271_0 ();
 b15zdnd11an1n64x5 FILLER_271_64 ();
 b15zdnd11an1n64x5 FILLER_271_128 ();
 b15zdnd11an1n64x5 FILLER_271_192 ();
 b15zdnd11an1n64x5 FILLER_271_256 ();
 b15zdnd11an1n64x5 FILLER_271_320 ();
 b15zdnd11an1n64x5 FILLER_271_384 ();
 b15zdnd11an1n64x5 FILLER_271_448 ();
 b15zdnd11an1n64x5 FILLER_271_512 ();
 b15zdnd11an1n64x5 FILLER_271_576 ();
 b15zdnd11an1n64x5 FILLER_271_640 ();
 b15zdnd11an1n64x5 FILLER_271_704 ();
 b15zdnd11an1n64x5 FILLER_271_768 ();
 b15zdnd11an1n64x5 FILLER_271_832 ();
 b15zdnd11an1n64x5 FILLER_271_896 ();
 b15zdnd11an1n64x5 FILLER_271_960 ();
 b15zdnd11an1n64x5 FILLER_271_1024 ();
 b15zdnd11an1n64x5 FILLER_271_1088 ();
 b15zdnd11an1n64x5 FILLER_271_1152 ();
 b15zdnd11an1n64x5 FILLER_271_1216 ();
 b15zdnd11an1n64x5 FILLER_271_1280 ();
 b15zdnd11an1n64x5 FILLER_271_1344 ();
 b15zdnd11an1n64x5 FILLER_271_1408 ();
 b15zdnd11an1n64x5 FILLER_271_1472 ();
 b15zdnd11an1n64x5 FILLER_271_1536 ();
 b15zdnd11an1n64x5 FILLER_271_1600 ();
 b15zdnd11an1n64x5 FILLER_271_1664 ();
 b15zdnd11an1n64x5 FILLER_271_1728 ();
 b15zdnd11an1n64x5 FILLER_271_1792 ();
 b15zdnd11an1n64x5 FILLER_271_1856 ();
 b15zdnd11an1n64x5 FILLER_271_1920 ();
 b15zdnd11an1n64x5 FILLER_271_1984 ();
 b15zdnd11an1n64x5 FILLER_271_2048 ();
 b15zdnd11an1n64x5 FILLER_271_2112 ();
 b15zdnd11an1n64x5 FILLER_271_2176 ();
 b15zdnd11an1n32x5 FILLER_271_2240 ();
 b15zdnd11an1n08x5 FILLER_271_2272 ();
 b15zdnd11an1n04x5 FILLER_271_2280 ();
 b15zdnd11an1n64x5 FILLER_272_8 ();
 b15zdnd11an1n64x5 FILLER_272_72 ();
 b15zdnd11an1n64x5 FILLER_272_136 ();
 b15zdnd11an1n64x5 FILLER_272_200 ();
 b15zdnd11an1n64x5 FILLER_272_264 ();
 b15zdnd11an1n64x5 FILLER_272_328 ();
 b15zdnd11an1n64x5 FILLER_272_392 ();
 b15zdnd11an1n64x5 FILLER_272_456 ();
 b15zdnd11an1n64x5 FILLER_272_520 ();
 b15zdnd11an1n64x5 FILLER_272_584 ();
 b15zdnd11an1n64x5 FILLER_272_648 ();
 b15zdnd11an1n04x5 FILLER_272_712 ();
 b15zdnd00an1n02x5 FILLER_272_716 ();
 b15zdnd11an1n64x5 FILLER_272_726 ();
 b15zdnd11an1n64x5 FILLER_272_790 ();
 b15zdnd11an1n64x5 FILLER_272_854 ();
 b15zdnd11an1n64x5 FILLER_272_918 ();
 b15zdnd11an1n64x5 FILLER_272_982 ();
 b15zdnd11an1n64x5 FILLER_272_1046 ();
 b15zdnd11an1n64x5 FILLER_272_1110 ();
 b15zdnd11an1n64x5 FILLER_272_1174 ();
 b15zdnd11an1n64x5 FILLER_272_1238 ();
 b15zdnd11an1n64x5 FILLER_272_1302 ();
 b15zdnd11an1n64x5 FILLER_272_1366 ();
 b15zdnd11an1n64x5 FILLER_272_1430 ();
 b15zdnd11an1n64x5 FILLER_272_1494 ();
 b15zdnd11an1n64x5 FILLER_272_1558 ();
 b15zdnd11an1n64x5 FILLER_272_1622 ();
 b15zdnd11an1n64x5 FILLER_272_1686 ();
 b15zdnd11an1n64x5 FILLER_272_1750 ();
 b15zdnd11an1n64x5 FILLER_272_1814 ();
 b15zdnd11an1n64x5 FILLER_272_1878 ();
 b15zdnd11an1n64x5 FILLER_272_1942 ();
 b15zdnd11an1n64x5 FILLER_272_2006 ();
 b15zdnd11an1n64x5 FILLER_272_2070 ();
 b15zdnd11an1n16x5 FILLER_272_2134 ();
 b15zdnd11an1n04x5 FILLER_272_2150 ();
 b15zdnd11an1n64x5 FILLER_272_2162 ();
 b15zdnd11an1n32x5 FILLER_272_2226 ();
 b15zdnd11an1n16x5 FILLER_272_2258 ();
 b15zdnd00an1n02x5 FILLER_272_2274 ();
 b15zdnd11an1n64x5 FILLER_273_0 ();
 b15zdnd11an1n64x5 FILLER_273_64 ();
 b15zdnd11an1n64x5 FILLER_273_128 ();
 b15zdnd11an1n64x5 FILLER_273_192 ();
 b15zdnd11an1n64x5 FILLER_273_256 ();
 b15zdnd11an1n64x5 FILLER_273_320 ();
 b15zdnd11an1n64x5 FILLER_273_384 ();
 b15zdnd11an1n64x5 FILLER_273_448 ();
 b15zdnd11an1n64x5 FILLER_273_512 ();
 b15zdnd11an1n64x5 FILLER_273_576 ();
 b15zdnd11an1n64x5 FILLER_273_640 ();
 b15zdnd11an1n64x5 FILLER_273_704 ();
 b15zdnd11an1n64x5 FILLER_273_768 ();
 b15zdnd11an1n64x5 FILLER_273_832 ();
 b15zdnd11an1n64x5 FILLER_273_896 ();
 b15zdnd11an1n64x5 FILLER_273_960 ();
 b15zdnd11an1n64x5 FILLER_273_1024 ();
 b15zdnd11an1n64x5 FILLER_273_1088 ();
 b15zdnd11an1n64x5 FILLER_273_1152 ();
 b15zdnd11an1n64x5 FILLER_273_1216 ();
 b15zdnd11an1n64x5 FILLER_273_1280 ();
 b15zdnd11an1n64x5 FILLER_273_1344 ();
 b15zdnd11an1n64x5 FILLER_273_1408 ();
 b15zdnd11an1n64x5 FILLER_273_1472 ();
 b15zdnd11an1n64x5 FILLER_273_1536 ();
 b15zdnd11an1n64x5 FILLER_273_1600 ();
 b15zdnd11an1n64x5 FILLER_273_1664 ();
 b15zdnd11an1n64x5 FILLER_273_1728 ();
 b15zdnd11an1n64x5 FILLER_273_1792 ();
 b15zdnd11an1n64x5 FILLER_273_1856 ();
 b15zdnd11an1n64x5 FILLER_273_1920 ();
 b15zdnd11an1n64x5 FILLER_273_1984 ();
 b15zdnd11an1n64x5 FILLER_273_2048 ();
 b15zdnd11an1n64x5 FILLER_273_2112 ();
 b15zdnd11an1n64x5 FILLER_273_2176 ();
 b15zdnd11an1n32x5 FILLER_273_2240 ();
 b15zdnd11an1n08x5 FILLER_273_2272 ();
 b15zdnd11an1n04x5 FILLER_273_2280 ();
 b15zdnd11an1n64x5 FILLER_274_8 ();
 b15zdnd11an1n64x5 FILLER_274_72 ();
 b15zdnd11an1n64x5 FILLER_274_136 ();
 b15zdnd11an1n64x5 FILLER_274_200 ();
 b15zdnd11an1n64x5 FILLER_274_264 ();
 b15zdnd11an1n64x5 FILLER_274_328 ();
 b15zdnd11an1n64x5 FILLER_274_392 ();
 b15zdnd11an1n64x5 FILLER_274_456 ();
 b15zdnd11an1n64x5 FILLER_274_520 ();
 b15zdnd11an1n64x5 FILLER_274_584 ();
 b15zdnd11an1n64x5 FILLER_274_648 ();
 b15zdnd11an1n04x5 FILLER_274_712 ();
 b15zdnd00an1n02x5 FILLER_274_716 ();
 b15zdnd11an1n64x5 FILLER_274_726 ();
 b15zdnd11an1n64x5 FILLER_274_790 ();
 b15zdnd11an1n64x5 FILLER_274_854 ();
 b15zdnd11an1n64x5 FILLER_274_918 ();
 b15zdnd11an1n64x5 FILLER_274_982 ();
 b15zdnd11an1n64x5 FILLER_274_1046 ();
 b15zdnd11an1n64x5 FILLER_274_1110 ();
 b15zdnd11an1n64x5 FILLER_274_1174 ();
 b15zdnd11an1n64x5 FILLER_274_1238 ();
 b15zdnd11an1n64x5 FILLER_274_1302 ();
 b15zdnd11an1n64x5 FILLER_274_1366 ();
 b15zdnd11an1n64x5 FILLER_274_1430 ();
 b15zdnd11an1n64x5 FILLER_274_1494 ();
 b15zdnd11an1n64x5 FILLER_274_1558 ();
 b15zdnd11an1n64x5 FILLER_274_1622 ();
 b15zdnd11an1n64x5 FILLER_274_1686 ();
 b15zdnd11an1n64x5 FILLER_274_1750 ();
 b15zdnd11an1n64x5 FILLER_274_1814 ();
 b15zdnd11an1n64x5 FILLER_274_1878 ();
 b15zdnd11an1n64x5 FILLER_274_1942 ();
 b15zdnd11an1n64x5 FILLER_274_2006 ();
 b15zdnd11an1n64x5 FILLER_274_2070 ();
 b15zdnd11an1n16x5 FILLER_274_2134 ();
 b15zdnd11an1n04x5 FILLER_274_2150 ();
 b15zdnd11an1n64x5 FILLER_274_2162 ();
 b15zdnd11an1n32x5 FILLER_274_2226 ();
 b15zdnd11an1n16x5 FILLER_274_2258 ();
 b15zdnd00an1n02x5 FILLER_274_2274 ();
 b15zdnd11an1n64x5 FILLER_275_0 ();
 b15zdnd11an1n64x5 FILLER_275_64 ();
 b15zdnd11an1n64x5 FILLER_275_128 ();
 b15zdnd11an1n64x5 FILLER_275_192 ();
 b15zdnd11an1n64x5 FILLER_275_256 ();
 b15zdnd11an1n64x5 FILLER_275_320 ();
 b15zdnd11an1n64x5 FILLER_275_384 ();
 b15zdnd11an1n64x5 FILLER_275_448 ();
 b15zdnd11an1n64x5 FILLER_275_512 ();
 b15zdnd11an1n64x5 FILLER_275_576 ();
 b15zdnd11an1n64x5 FILLER_275_640 ();
 b15zdnd11an1n64x5 FILLER_275_704 ();
 b15zdnd11an1n64x5 FILLER_275_768 ();
 b15zdnd11an1n64x5 FILLER_275_832 ();
 b15zdnd11an1n64x5 FILLER_275_896 ();
 b15zdnd11an1n64x5 FILLER_275_960 ();
 b15zdnd11an1n64x5 FILLER_275_1024 ();
 b15zdnd11an1n64x5 FILLER_275_1088 ();
 b15zdnd11an1n64x5 FILLER_275_1152 ();
 b15zdnd11an1n64x5 FILLER_275_1216 ();
 b15zdnd11an1n64x5 FILLER_275_1280 ();
 b15zdnd11an1n64x5 FILLER_275_1344 ();
 b15zdnd11an1n64x5 FILLER_275_1408 ();
 b15zdnd11an1n64x5 FILLER_275_1472 ();
 b15zdnd11an1n64x5 FILLER_275_1536 ();
 b15zdnd11an1n64x5 FILLER_275_1600 ();
 b15zdnd11an1n64x5 FILLER_275_1664 ();
 b15zdnd11an1n64x5 FILLER_275_1728 ();
 b15zdnd11an1n64x5 FILLER_275_1792 ();
 b15zdnd11an1n64x5 FILLER_275_1856 ();
 b15zdnd11an1n64x5 FILLER_275_1920 ();
 b15zdnd11an1n64x5 FILLER_275_1984 ();
 b15zdnd11an1n64x5 FILLER_275_2048 ();
 b15zdnd11an1n64x5 FILLER_275_2112 ();
 b15zdnd11an1n64x5 FILLER_275_2176 ();
 b15zdnd11an1n32x5 FILLER_275_2240 ();
 b15zdnd11an1n08x5 FILLER_275_2272 ();
 b15zdnd11an1n04x5 FILLER_275_2280 ();
 b15zdnd11an1n64x5 FILLER_276_8 ();
 b15zdnd11an1n64x5 FILLER_276_72 ();
 b15zdnd11an1n64x5 FILLER_276_136 ();
 b15zdnd11an1n64x5 FILLER_276_200 ();
 b15zdnd11an1n64x5 FILLER_276_264 ();
 b15zdnd11an1n64x5 FILLER_276_328 ();
 b15zdnd11an1n64x5 FILLER_276_392 ();
 b15zdnd11an1n64x5 FILLER_276_456 ();
 b15zdnd11an1n64x5 FILLER_276_520 ();
 b15zdnd11an1n64x5 FILLER_276_584 ();
 b15zdnd11an1n64x5 FILLER_276_648 ();
 b15zdnd11an1n04x5 FILLER_276_712 ();
 b15zdnd00an1n02x5 FILLER_276_716 ();
 b15zdnd11an1n64x5 FILLER_276_726 ();
 b15zdnd11an1n64x5 FILLER_276_790 ();
 b15zdnd11an1n64x5 FILLER_276_854 ();
 b15zdnd11an1n64x5 FILLER_276_918 ();
 b15zdnd11an1n64x5 FILLER_276_982 ();
 b15zdnd11an1n64x5 FILLER_276_1046 ();
 b15zdnd11an1n64x5 FILLER_276_1110 ();
 b15zdnd11an1n64x5 FILLER_276_1174 ();
 b15zdnd11an1n64x5 FILLER_276_1238 ();
 b15zdnd11an1n64x5 FILLER_276_1302 ();
 b15zdnd11an1n64x5 FILLER_276_1366 ();
 b15zdnd11an1n64x5 FILLER_276_1430 ();
 b15zdnd11an1n64x5 FILLER_276_1494 ();
 b15zdnd11an1n64x5 FILLER_276_1558 ();
 b15zdnd11an1n64x5 FILLER_276_1622 ();
 b15zdnd11an1n64x5 FILLER_276_1686 ();
 b15zdnd11an1n64x5 FILLER_276_1750 ();
 b15zdnd11an1n64x5 FILLER_276_1814 ();
 b15zdnd11an1n64x5 FILLER_276_1878 ();
 b15zdnd11an1n64x5 FILLER_276_1942 ();
 b15zdnd11an1n64x5 FILLER_276_2006 ();
 b15zdnd11an1n64x5 FILLER_276_2070 ();
 b15zdnd11an1n16x5 FILLER_276_2134 ();
 b15zdnd11an1n04x5 FILLER_276_2150 ();
 b15zdnd11an1n64x5 FILLER_276_2162 ();
 b15zdnd11an1n32x5 FILLER_276_2226 ();
 b15zdnd11an1n16x5 FILLER_276_2258 ();
 b15zdnd00an1n02x5 FILLER_276_2274 ();
 b15zdnd11an1n64x5 FILLER_277_0 ();
 b15zdnd11an1n64x5 FILLER_277_64 ();
 b15zdnd11an1n64x5 FILLER_277_128 ();
 b15zdnd11an1n64x5 FILLER_277_192 ();
 b15zdnd11an1n64x5 FILLER_277_256 ();
 b15zdnd11an1n64x5 FILLER_277_320 ();
 b15zdnd11an1n64x5 FILLER_277_384 ();
 b15zdnd11an1n64x5 FILLER_277_448 ();
 b15zdnd11an1n64x5 FILLER_277_512 ();
 b15zdnd11an1n64x5 FILLER_277_576 ();
 b15zdnd11an1n64x5 FILLER_277_640 ();
 b15zdnd11an1n64x5 FILLER_277_704 ();
 b15zdnd11an1n64x5 FILLER_277_768 ();
 b15zdnd11an1n64x5 FILLER_277_832 ();
 b15zdnd11an1n64x5 FILLER_277_896 ();
 b15zdnd11an1n64x5 FILLER_277_960 ();
 b15zdnd11an1n64x5 FILLER_277_1024 ();
 b15zdnd11an1n64x5 FILLER_277_1088 ();
 b15zdnd11an1n64x5 FILLER_277_1152 ();
 b15zdnd11an1n64x5 FILLER_277_1216 ();
 b15zdnd11an1n64x5 FILLER_277_1280 ();
 b15zdnd11an1n64x5 FILLER_277_1344 ();
 b15zdnd11an1n64x5 FILLER_277_1408 ();
 b15zdnd11an1n64x5 FILLER_277_1472 ();
 b15zdnd11an1n64x5 FILLER_277_1536 ();
 b15zdnd11an1n64x5 FILLER_277_1600 ();
 b15zdnd11an1n64x5 FILLER_277_1664 ();
 b15zdnd11an1n64x5 FILLER_277_1728 ();
 b15zdnd11an1n64x5 FILLER_277_1792 ();
 b15zdnd11an1n64x5 FILLER_277_1856 ();
 b15zdnd11an1n64x5 FILLER_277_1920 ();
 b15zdnd11an1n64x5 FILLER_277_1984 ();
 b15zdnd11an1n64x5 FILLER_277_2048 ();
 b15zdnd11an1n64x5 FILLER_277_2112 ();
 b15zdnd11an1n64x5 FILLER_277_2176 ();
 b15zdnd11an1n32x5 FILLER_277_2240 ();
 b15zdnd11an1n08x5 FILLER_277_2272 ();
 b15zdnd11an1n04x5 FILLER_277_2280 ();
 b15zdnd11an1n64x5 FILLER_278_8 ();
 b15zdnd11an1n64x5 FILLER_278_72 ();
 b15zdnd11an1n64x5 FILLER_278_136 ();
 b15zdnd11an1n64x5 FILLER_278_200 ();
 b15zdnd11an1n64x5 FILLER_278_264 ();
 b15zdnd11an1n64x5 FILLER_278_328 ();
 b15zdnd11an1n64x5 FILLER_278_392 ();
 b15zdnd11an1n64x5 FILLER_278_456 ();
 b15zdnd11an1n64x5 FILLER_278_520 ();
 b15zdnd11an1n64x5 FILLER_278_584 ();
 b15zdnd11an1n64x5 FILLER_278_648 ();
 b15zdnd11an1n04x5 FILLER_278_712 ();
 b15zdnd00an1n02x5 FILLER_278_716 ();
 b15zdnd11an1n64x5 FILLER_278_726 ();
 b15zdnd11an1n64x5 FILLER_278_790 ();
 b15zdnd11an1n64x5 FILLER_278_854 ();
 b15zdnd11an1n64x5 FILLER_278_918 ();
 b15zdnd11an1n64x5 FILLER_278_982 ();
 b15zdnd11an1n64x5 FILLER_278_1046 ();
 b15zdnd11an1n64x5 FILLER_278_1110 ();
 b15zdnd11an1n64x5 FILLER_278_1174 ();
 b15zdnd11an1n64x5 FILLER_278_1238 ();
 b15zdnd11an1n64x5 FILLER_278_1302 ();
 b15zdnd11an1n64x5 FILLER_278_1366 ();
 b15zdnd11an1n64x5 FILLER_278_1430 ();
 b15zdnd11an1n64x5 FILLER_278_1494 ();
 b15zdnd11an1n64x5 FILLER_278_1558 ();
 b15zdnd11an1n64x5 FILLER_278_1622 ();
 b15zdnd11an1n64x5 FILLER_278_1686 ();
 b15zdnd11an1n64x5 FILLER_278_1750 ();
 b15zdnd11an1n64x5 FILLER_278_1814 ();
 b15zdnd11an1n64x5 FILLER_278_1878 ();
 b15zdnd11an1n64x5 FILLER_278_1942 ();
 b15zdnd11an1n64x5 FILLER_278_2006 ();
 b15zdnd11an1n64x5 FILLER_278_2070 ();
 b15zdnd11an1n16x5 FILLER_278_2134 ();
 b15zdnd11an1n04x5 FILLER_278_2150 ();
 b15zdnd11an1n64x5 FILLER_278_2162 ();
 b15zdnd11an1n32x5 FILLER_278_2226 ();
 b15zdnd11an1n16x5 FILLER_278_2258 ();
 b15zdnd00an1n02x5 FILLER_278_2274 ();
 b15zdnd11an1n64x5 FILLER_279_0 ();
 b15zdnd11an1n64x5 FILLER_279_64 ();
 b15zdnd11an1n64x5 FILLER_279_128 ();
 b15zdnd11an1n64x5 FILLER_279_192 ();
 b15zdnd11an1n64x5 FILLER_279_256 ();
 b15zdnd11an1n64x5 FILLER_279_320 ();
 b15zdnd11an1n64x5 FILLER_279_384 ();
 b15zdnd11an1n64x5 FILLER_279_448 ();
 b15zdnd11an1n64x5 FILLER_279_512 ();
 b15zdnd11an1n64x5 FILLER_279_576 ();
 b15zdnd11an1n64x5 FILLER_279_640 ();
 b15zdnd11an1n64x5 FILLER_279_704 ();
 b15zdnd11an1n64x5 FILLER_279_768 ();
 b15zdnd11an1n64x5 FILLER_279_832 ();
 b15zdnd11an1n64x5 FILLER_279_896 ();
 b15zdnd11an1n64x5 FILLER_279_960 ();
 b15zdnd11an1n64x5 FILLER_279_1024 ();
 b15zdnd11an1n64x5 FILLER_279_1088 ();
 b15zdnd11an1n64x5 FILLER_279_1152 ();
 b15zdnd11an1n64x5 FILLER_279_1216 ();
 b15zdnd11an1n64x5 FILLER_279_1280 ();
 b15zdnd11an1n64x5 FILLER_279_1344 ();
 b15zdnd11an1n64x5 FILLER_279_1408 ();
 b15zdnd11an1n64x5 FILLER_279_1472 ();
 b15zdnd11an1n64x5 FILLER_279_1536 ();
 b15zdnd11an1n64x5 FILLER_279_1600 ();
 b15zdnd11an1n64x5 FILLER_279_1664 ();
 b15zdnd11an1n64x5 FILLER_279_1728 ();
 b15zdnd11an1n64x5 FILLER_279_1792 ();
 b15zdnd11an1n64x5 FILLER_279_1856 ();
 b15zdnd11an1n64x5 FILLER_279_1920 ();
 b15zdnd11an1n64x5 FILLER_279_1984 ();
 b15zdnd11an1n64x5 FILLER_279_2048 ();
 b15zdnd11an1n64x5 FILLER_279_2112 ();
 b15zdnd11an1n64x5 FILLER_279_2176 ();
 b15zdnd11an1n32x5 FILLER_279_2240 ();
 b15zdnd11an1n08x5 FILLER_279_2272 ();
 b15zdnd11an1n04x5 FILLER_279_2280 ();
 b15zdnd11an1n64x5 FILLER_280_8 ();
 b15zdnd11an1n64x5 FILLER_280_72 ();
 b15zdnd11an1n64x5 FILLER_280_136 ();
 b15zdnd11an1n64x5 FILLER_280_200 ();
 b15zdnd11an1n64x5 FILLER_280_264 ();
 b15zdnd11an1n64x5 FILLER_280_328 ();
 b15zdnd11an1n64x5 FILLER_280_392 ();
 b15zdnd11an1n64x5 FILLER_280_456 ();
 b15zdnd11an1n64x5 FILLER_280_520 ();
 b15zdnd11an1n64x5 FILLER_280_584 ();
 b15zdnd11an1n64x5 FILLER_280_648 ();
 b15zdnd11an1n04x5 FILLER_280_712 ();
 b15zdnd00an1n02x5 FILLER_280_716 ();
 b15zdnd11an1n64x5 FILLER_280_726 ();
 b15zdnd11an1n64x5 FILLER_280_790 ();
 b15zdnd11an1n64x5 FILLER_280_854 ();
 b15zdnd11an1n64x5 FILLER_280_918 ();
 b15zdnd11an1n64x5 FILLER_280_982 ();
 b15zdnd11an1n64x5 FILLER_280_1046 ();
 b15zdnd11an1n64x5 FILLER_280_1110 ();
 b15zdnd11an1n64x5 FILLER_280_1174 ();
 b15zdnd11an1n64x5 FILLER_280_1238 ();
 b15zdnd11an1n64x5 FILLER_280_1302 ();
 b15zdnd11an1n64x5 FILLER_280_1366 ();
 b15zdnd11an1n64x5 FILLER_280_1430 ();
 b15zdnd11an1n64x5 FILLER_280_1494 ();
 b15zdnd11an1n64x5 FILLER_280_1558 ();
 b15zdnd11an1n64x5 FILLER_280_1622 ();
 b15zdnd11an1n64x5 FILLER_280_1686 ();
 b15zdnd11an1n64x5 FILLER_280_1750 ();
 b15zdnd11an1n64x5 FILLER_280_1814 ();
 b15zdnd11an1n64x5 FILLER_280_1878 ();
 b15zdnd11an1n64x5 FILLER_280_1942 ();
 b15zdnd11an1n64x5 FILLER_280_2006 ();
 b15zdnd11an1n64x5 FILLER_280_2070 ();
 b15zdnd11an1n16x5 FILLER_280_2134 ();
 b15zdnd11an1n04x5 FILLER_280_2150 ();
 b15zdnd11an1n64x5 FILLER_280_2162 ();
 b15zdnd11an1n32x5 FILLER_280_2226 ();
 b15zdnd11an1n16x5 FILLER_280_2258 ();
 b15zdnd00an1n02x5 FILLER_280_2274 ();
 b15zdnd11an1n64x5 FILLER_281_0 ();
 b15zdnd11an1n64x5 FILLER_281_64 ();
 b15zdnd11an1n64x5 FILLER_281_128 ();
 b15zdnd11an1n64x5 FILLER_281_192 ();
 b15zdnd11an1n64x5 FILLER_281_256 ();
 b15zdnd11an1n64x5 FILLER_281_320 ();
 b15zdnd11an1n64x5 FILLER_281_384 ();
 b15zdnd11an1n64x5 FILLER_281_448 ();
 b15zdnd11an1n64x5 FILLER_281_512 ();
 b15zdnd11an1n64x5 FILLER_281_576 ();
 b15zdnd11an1n64x5 FILLER_281_640 ();
 b15zdnd11an1n64x5 FILLER_281_704 ();
 b15zdnd11an1n64x5 FILLER_281_768 ();
 b15zdnd11an1n64x5 FILLER_281_832 ();
 b15zdnd11an1n64x5 FILLER_281_896 ();
 b15zdnd11an1n64x5 FILLER_281_960 ();
 b15zdnd11an1n64x5 FILLER_281_1024 ();
 b15zdnd11an1n64x5 FILLER_281_1088 ();
 b15zdnd11an1n64x5 FILLER_281_1152 ();
 b15zdnd11an1n64x5 FILLER_281_1216 ();
 b15zdnd11an1n64x5 FILLER_281_1280 ();
 b15zdnd11an1n64x5 FILLER_281_1344 ();
 b15zdnd11an1n64x5 FILLER_281_1408 ();
 b15zdnd11an1n64x5 FILLER_281_1472 ();
 b15zdnd11an1n64x5 FILLER_281_1536 ();
 b15zdnd11an1n64x5 FILLER_281_1600 ();
 b15zdnd11an1n32x5 FILLER_281_1664 ();
 b15zdnd11an1n16x5 FILLER_281_1696 ();
 b15zdnd00an1n02x5 FILLER_281_1712 ();
 b15zdnd11an1n64x5 FILLER_281_1730 ();
 b15zdnd11an1n64x5 FILLER_281_1794 ();
 b15zdnd11an1n64x5 FILLER_281_1858 ();
 b15zdnd11an1n64x5 FILLER_281_1922 ();
 b15zdnd11an1n64x5 FILLER_281_1986 ();
 b15zdnd11an1n64x5 FILLER_281_2050 ();
 b15zdnd11an1n64x5 FILLER_281_2114 ();
 b15zdnd11an1n64x5 FILLER_281_2178 ();
 b15zdnd11an1n32x5 FILLER_281_2242 ();
 b15zdnd11an1n08x5 FILLER_281_2274 ();
 b15zdnd00an1n02x5 FILLER_281_2282 ();
 b15zdnd11an1n64x5 FILLER_282_8 ();
 b15zdnd11an1n64x5 FILLER_282_72 ();
 b15zdnd11an1n64x5 FILLER_282_136 ();
 b15zdnd11an1n64x5 FILLER_282_200 ();
 b15zdnd11an1n64x5 FILLER_282_264 ();
 b15zdnd11an1n64x5 FILLER_282_328 ();
 b15zdnd11an1n64x5 FILLER_282_392 ();
 b15zdnd11an1n64x5 FILLER_282_456 ();
 b15zdnd11an1n64x5 FILLER_282_520 ();
 b15zdnd11an1n64x5 FILLER_282_584 ();
 b15zdnd11an1n64x5 FILLER_282_648 ();
 b15zdnd11an1n04x5 FILLER_282_712 ();
 b15zdnd00an1n02x5 FILLER_282_716 ();
 b15zdnd11an1n64x5 FILLER_282_726 ();
 b15zdnd11an1n64x5 FILLER_282_790 ();
 b15zdnd11an1n64x5 FILLER_282_854 ();
 b15zdnd11an1n64x5 FILLER_282_918 ();
 b15zdnd11an1n64x5 FILLER_282_982 ();
 b15zdnd11an1n64x5 FILLER_282_1046 ();
 b15zdnd11an1n64x5 FILLER_282_1110 ();
 b15zdnd11an1n64x5 FILLER_282_1174 ();
 b15zdnd11an1n64x5 FILLER_282_1238 ();
 b15zdnd11an1n64x5 FILLER_282_1302 ();
 b15zdnd11an1n64x5 FILLER_282_1366 ();
 b15zdnd11an1n64x5 FILLER_282_1430 ();
 b15zdnd11an1n64x5 FILLER_282_1494 ();
 b15zdnd11an1n64x5 FILLER_282_1558 ();
 b15zdnd11an1n64x5 FILLER_282_1622 ();
 b15zdnd11an1n64x5 FILLER_282_1686 ();
 b15zdnd11an1n64x5 FILLER_282_1750 ();
 b15zdnd11an1n64x5 FILLER_282_1814 ();
 b15zdnd11an1n64x5 FILLER_282_1878 ();
 b15zdnd11an1n64x5 FILLER_282_1942 ();
 b15zdnd11an1n64x5 FILLER_282_2006 ();
 b15zdnd11an1n64x5 FILLER_282_2070 ();
 b15zdnd11an1n16x5 FILLER_282_2134 ();
 b15zdnd11an1n04x5 FILLER_282_2150 ();
 b15zdnd11an1n64x5 FILLER_282_2162 ();
 b15zdnd11an1n32x5 FILLER_282_2226 ();
 b15zdnd11an1n16x5 FILLER_282_2258 ();
 b15zdnd00an1n02x5 FILLER_282_2274 ();
 b15zdnd11an1n64x5 FILLER_283_0 ();
 b15zdnd11an1n64x5 FILLER_283_64 ();
 b15zdnd11an1n64x5 FILLER_283_128 ();
 b15zdnd11an1n64x5 FILLER_283_192 ();
 b15zdnd11an1n64x5 FILLER_283_256 ();
 b15zdnd11an1n64x5 FILLER_283_320 ();
 b15zdnd11an1n64x5 FILLER_283_384 ();
 b15zdnd11an1n64x5 FILLER_283_448 ();
 b15zdnd11an1n64x5 FILLER_283_512 ();
 b15zdnd11an1n64x5 FILLER_283_576 ();
 b15zdnd11an1n64x5 FILLER_283_640 ();
 b15zdnd11an1n64x5 FILLER_283_704 ();
 b15zdnd11an1n64x5 FILLER_283_768 ();
 b15zdnd11an1n64x5 FILLER_283_832 ();
 b15zdnd11an1n64x5 FILLER_283_896 ();
 b15zdnd11an1n64x5 FILLER_283_960 ();
 b15zdnd11an1n64x5 FILLER_283_1024 ();
 b15zdnd11an1n64x5 FILLER_283_1088 ();
 b15zdnd11an1n64x5 FILLER_283_1152 ();
 b15zdnd11an1n64x5 FILLER_283_1216 ();
 b15zdnd11an1n64x5 FILLER_283_1280 ();
 b15zdnd11an1n64x5 FILLER_283_1344 ();
 b15zdnd11an1n64x5 FILLER_283_1408 ();
 b15zdnd11an1n64x5 FILLER_283_1472 ();
 b15zdnd11an1n64x5 FILLER_283_1536 ();
 b15zdnd11an1n64x5 FILLER_283_1600 ();
 b15zdnd11an1n64x5 FILLER_283_1664 ();
 b15zdnd11an1n64x5 FILLER_283_1728 ();
 b15zdnd11an1n64x5 FILLER_283_1792 ();
 b15zdnd11an1n64x5 FILLER_283_1856 ();
 b15zdnd11an1n64x5 FILLER_283_1920 ();
 b15zdnd11an1n64x5 FILLER_283_1984 ();
 b15zdnd11an1n64x5 FILLER_283_2048 ();
 b15zdnd11an1n64x5 FILLER_283_2112 ();
 b15zdnd11an1n64x5 FILLER_283_2176 ();
 b15zdnd11an1n32x5 FILLER_283_2240 ();
 b15zdnd11an1n08x5 FILLER_283_2272 ();
 b15zdnd11an1n04x5 FILLER_283_2280 ();
 b15zdnd11an1n64x5 FILLER_284_8 ();
 b15zdnd11an1n64x5 FILLER_284_72 ();
 b15zdnd11an1n64x5 FILLER_284_136 ();
 b15zdnd11an1n64x5 FILLER_284_200 ();
 b15zdnd11an1n64x5 FILLER_284_264 ();
 b15zdnd11an1n64x5 FILLER_284_328 ();
 b15zdnd11an1n64x5 FILLER_284_392 ();
 b15zdnd11an1n64x5 FILLER_284_456 ();
 b15zdnd11an1n64x5 FILLER_284_520 ();
 b15zdnd11an1n64x5 FILLER_284_584 ();
 b15zdnd11an1n64x5 FILLER_284_648 ();
 b15zdnd11an1n04x5 FILLER_284_712 ();
 b15zdnd00an1n02x5 FILLER_284_716 ();
 b15zdnd11an1n64x5 FILLER_284_726 ();
 b15zdnd11an1n64x5 FILLER_284_790 ();
 b15zdnd11an1n64x5 FILLER_284_854 ();
 b15zdnd11an1n64x5 FILLER_284_918 ();
 b15zdnd11an1n64x5 FILLER_284_982 ();
 b15zdnd11an1n64x5 FILLER_284_1046 ();
 b15zdnd11an1n64x5 FILLER_284_1110 ();
 b15zdnd11an1n64x5 FILLER_284_1174 ();
 b15zdnd11an1n64x5 FILLER_284_1238 ();
 b15zdnd11an1n64x5 FILLER_284_1302 ();
 b15zdnd11an1n64x5 FILLER_284_1366 ();
 b15zdnd11an1n64x5 FILLER_284_1430 ();
 b15zdnd11an1n64x5 FILLER_284_1494 ();
 b15zdnd11an1n64x5 FILLER_284_1558 ();
 b15zdnd11an1n64x5 FILLER_284_1622 ();
 b15zdnd11an1n64x5 FILLER_284_1686 ();
 b15zdnd11an1n64x5 FILLER_284_1750 ();
 b15zdnd11an1n64x5 FILLER_284_1814 ();
 b15zdnd11an1n64x5 FILLER_284_1878 ();
 b15zdnd11an1n64x5 FILLER_284_1942 ();
 b15zdnd11an1n64x5 FILLER_284_2006 ();
 b15zdnd11an1n64x5 FILLER_284_2070 ();
 b15zdnd11an1n16x5 FILLER_284_2134 ();
 b15zdnd11an1n04x5 FILLER_284_2150 ();
 b15zdnd11an1n64x5 FILLER_284_2162 ();
 b15zdnd11an1n32x5 FILLER_284_2226 ();
 b15zdnd11an1n16x5 FILLER_284_2258 ();
 b15zdnd00an1n02x5 FILLER_284_2274 ();
 b15zdnd11an1n64x5 FILLER_285_0 ();
 b15zdnd11an1n64x5 FILLER_285_64 ();
 b15zdnd11an1n64x5 FILLER_285_128 ();
 b15zdnd11an1n64x5 FILLER_285_192 ();
 b15zdnd11an1n64x5 FILLER_285_256 ();
 b15zdnd11an1n64x5 FILLER_285_320 ();
 b15zdnd11an1n64x5 FILLER_285_384 ();
 b15zdnd11an1n64x5 FILLER_285_448 ();
 b15zdnd11an1n64x5 FILLER_285_512 ();
 b15zdnd11an1n64x5 FILLER_285_576 ();
 b15zdnd11an1n64x5 FILLER_285_640 ();
 b15zdnd11an1n64x5 FILLER_285_704 ();
 b15zdnd11an1n64x5 FILLER_285_768 ();
 b15zdnd11an1n64x5 FILLER_285_832 ();
 b15zdnd11an1n64x5 FILLER_285_896 ();
 b15zdnd11an1n64x5 FILLER_285_960 ();
 b15zdnd11an1n64x5 FILLER_285_1024 ();
 b15zdnd11an1n64x5 FILLER_285_1088 ();
 b15zdnd11an1n64x5 FILLER_285_1152 ();
 b15zdnd11an1n64x5 FILLER_285_1216 ();
 b15zdnd11an1n64x5 FILLER_285_1280 ();
 b15zdnd11an1n32x5 FILLER_285_1344 ();
 b15zdnd11an1n04x5 FILLER_285_1376 ();
 b15zdnd00an1n02x5 FILLER_285_1380 ();
 b15zdnd11an1n64x5 FILLER_285_1398 ();
 b15zdnd11an1n64x5 FILLER_285_1462 ();
 b15zdnd11an1n64x5 FILLER_285_1526 ();
 b15zdnd11an1n64x5 FILLER_285_1590 ();
 b15zdnd11an1n64x5 FILLER_285_1654 ();
 b15zdnd11an1n64x5 FILLER_285_1718 ();
 b15zdnd11an1n64x5 FILLER_285_1782 ();
 b15zdnd11an1n64x5 FILLER_285_1846 ();
 b15zdnd11an1n64x5 FILLER_285_1910 ();
 b15zdnd11an1n64x5 FILLER_285_1974 ();
 b15zdnd11an1n64x5 FILLER_285_2038 ();
 b15zdnd11an1n64x5 FILLER_285_2102 ();
 b15zdnd11an1n64x5 FILLER_285_2166 ();
 b15zdnd11an1n32x5 FILLER_285_2230 ();
 b15zdnd11an1n16x5 FILLER_285_2262 ();
 b15zdnd11an1n04x5 FILLER_285_2278 ();
 b15zdnd00an1n02x5 FILLER_285_2282 ();
 b15zdnd11an1n64x5 FILLER_286_8 ();
 b15zdnd11an1n64x5 FILLER_286_72 ();
 b15zdnd11an1n64x5 FILLER_286_136 ();
 b15zdnd11an1n64x5 FILLER_286_200 ();
 b15zdnd11an1n64x5 FILLER_286_264 ();
 b15zdnd11an1n64x5 FILLER_286_328 ();
 b15zdnd11an1n64x5 FILLER_286_392 ();
 b15zdnd11an1n64x5 FILLER_286_456 ();
 b15zdnd11an1n64x5 FILLER_286_520 ();
 b15zdnd11an1n64x5 FILLER_286_584 ();
 b15zdnd11an1n64x5 FILLER_286_648 ();
 b15zdnd11an1n04x5 FILLER_286_712 ();
 b15zdnd00an1n02x5 FILLER_286_716 ();
 b15zdnd11an1n64x5 FILLER_286_726 ();
 b15zdnd11an1n64x5 FILLER_286_790 ();
 b15zdnd11an1n64x5 FILLER_286_854 ();
 b15zdnd11an1n64x5 FILLER_286_918 ();
 b15zdnd11an1n64x5 FILLER_286_982 ();
 b15zdnd11an1n64x5 FILLER_286_1046 ();
 b15zdnd11an1n64x5 FILLER_286_1110 ();
 b15zdnd11an1n64x5 FILLER_286_1174 ();
 b15zdnd11an1n64x5 FILLER_286_1238 ();
 b15zdnd11an1n64x5 FILLER_286_1302 ();
 b15zdnd11an1n64x5 FILLER_286_1366 ();
 b15zdnd11an1n64x5 FILLER_286_1430 ();
 b15zdnd11an1n64x5 FILLER_286_1494 ();
 b15zdnd11an1n64x5 FILLER_286_1558 ();
 b15zdnd11an1n64x5 FILLER_286_1622 ();
 b15zdnd11an1n64x5 FILLER_286_1686 ();
 b15zdnd11an1n64x5 FILLER_286_1750 ();
 b15zdnd11an1n64x5 FILLER_286_1814 ();
 b15zdnd11an1n64x5 FILLER_286_1878 ();
 b15zdnd11an1n64x5 FILLER_286_1942 ();
 b15zdnd11an1n64x5 FILLER_286_2006 ();
 b15zdnd11an1n64x5 FILLER_286_2070 ();
 b15zdnd11an1n16x5 FILLER_286_2134 ();
 b15zdnd11an1n04x5 FILLER_286_2150 ();
 b15zdnd11an1n64x5 FILLER_286_2162 ();
 b15zdnd11an1n32x5 FILLER_286_2226 ();
 b15zdnd11an1n16x5 FILLER_286_2258 ();
 b15zdnd00an1n02x5 FILLER_286_2274 ();
 b15zdnd11an1n64x5 FILLER_287_0 ();
 b15zdnd11an1n64x5 FILLER_287_64 ();
 b15zdnd11an1n64x5 FILLER_287_128 ();
 b15zdnd11an1n64x5 FILLER_287_192 ();
 b15zdnd11an1n64x5 FILLER_287_256 ();
 b15zdnd11an1n64x5 FILLER_287_320 ();
 b15zdnd11an1n64x5 FILLER_287_384 ();
 b15zdnd11an1n64x5 FILLER_287_448 ();
 b15zdnd11an1n64x5 FILLER_287_512 ();
 b15zdnd11an1n64x5 FILLER_287_576 ();
 b15zdnd11an1n64x5 FILLER_287_640 ();
 b15zdnd11an1n64x5 FILLER_287_704 ();
 b15zdnd11an1n64x5 FILLER_287_768 ();
 b15zdnd11an1n64x5 FILLER_287_832 ();
 b15zdnd11an1n64x5 FILLER_287_896 ();
 b15zdnd11an1n64x5 FILLER_287_960 ();
 b15zdnd11an1n64x5 FILLER_287_1024 ();
 b15zdnd11an1n64x5 FILLER_287_1088 ();
 b15zdnd11an1n64x5 FILLER_287_1152 ();
 b15zdnd11an1n64x5 FILLER_287_1216 ();
 b15zdnd11an1n64x5 FILLER_287_1280 ();
 b15zdnd11an1n64x5 FILLER_287_1344 ();
 b15zdnd11an1n64x5 FILLER_287_1408 ();
 b15zdnd11an1n64x5 FILLER_287_1472 ();
 b15zdnd11an1n64x5 FILLER_287_1536 ();
 b15zdnd11an1n64x5 FILLER_287_1600 ();
 b15zdnd11an1n64x5 FILLER_287_1664 ();
 b15zdnd11an1n64x5 FILLER_287_1728 ();
 b15zdnd11an1n64x5 FILLER_287_1792 ();
 b15zdnd11an1n64x5 FILLER_287_1856 ();
 b15zdnd11an1n64x5 FILLER_287_1920 ();
 b15zdnd11an1n64x5 FILLER_287_1984 ();
 b15zdnd11an1n64x5 FILLER_287_2048 ();
 b15zdnd11an1n64x5 FILLER_287_2112 ();
 b15zdnd11an1n64x5 FILLER_287_2176 ();
 b15zdnd11an1n32x5 FILLER_287_2240 ();
 b15zdnd11an1n08x5 FILLER_287_2272 ();
 b15zdnd11an1n04x5 FILLER_287_2280 ();
 b15zdnd11an1n64x5 FILLER_288_8 ();
 b15zdnd11an1n64x5 FILLER_288_72 ();
 b15zdnd11an1n64x5 FILLER_288_136 ();
 b15zdnd11an1n64x5 FILLER_288_200 ();
 b15zdnd11an1n64x5 FILLER_288_264 ();
 b15zdnd11an1n64x5 FILLER_288_328 ();
 b15zdnd11an1n64x5 FILLER_288_392 ();
 b15zdnd11an1n64x5 FILLER_288_456 ();
 b15zdnd11an1n64x5 FILLER_288_520 ();
 b15zdnd11an1n64x5 FILLER_288_584 ();
 b15zdnd11an1n64x5 FILLER_288_648 ();
 b15zdnd11an1n04x5 FILLER_288_712 ();
 b15zdnd00an1n02x5 FILLER_288_716 ();
 b15zdnd11an1n64x5 FILLER_288_726 ();
 b15zdnd11an1n64x5 FILLER_288_790 ();
 b15zdnd11an1n64x5 FILLER_288_854 ();
 b15zdnd11an1n64x5 FILLER_288_918 ();
 b15zdnd11an1n64x5 FILLER_288_982 ();
 b15zdnd11an1n64x5 FILLER_288_1046 ();
 b15zdnd11an1n64x5 FILLER_288_1110 ();
 b15zdnd11an1n64x5 FILLER_288_1174 ();
 b15zdnd11an1n64x5 FILLER_288_1238 ();
 b15zdnd11an1n64x5 FILLER_288_1302 ();
 b15zdnd11an1n64x5 FILLER_288_1366 ();
 b15zdnd11an1n64x5 FILLER_288_1430 ();
 b15zdnd11an1n64x5 FILLER_288_1494 ();
 b15zdnd11an1n64x5 FILLER_288_1558 ();
 b15zdnd11an1n64x5 FILLER_288_1622 ();
 b15zdnd11an1n64x5 FILLER_288_1686 ();
 b15zdnd11an1n64x5 FILLER_288_1750 ();
 b15zdnd11an1n64x5 FILLER_288_1814 ();
 b15zdnd11an1n64x5 FILLER_288_1878 ();
 b15zdnd11an1n64x5 FILLER_288_1942 ();
 b15zdnd11an1n64x5 FILLER_288_2006 ();
 b15zdnd11an1n64x5 FILLER_288_2070 ();
 b15zdnd11an1n16x5 FILLER_288_2134 ();
 b15zdnd11an1n04x5 FILLER_288_2150 ();
 b15zdnd11an1n64x5 FILLER_288_2162 ();
 b15zdnd11an1n32x5 FILLER_288_2226 ();
 b15zdnd11an1n16x5 FILLER_288_2258 ();
 b15zdnd00an1n02x5 FILLER_288_2274 ();
 b15zdnd11an1n64x5 FILLER_289_0 ();
 b15zdnd11an1n64x5 FILLER_289_64 ();
 b15zdnd11an1n64x5 FILLER_289_128 ();
 b15zdnd11an1n64x5 FILLER_289_192 ();
 b15zdnd11an1n64x5 FILLER_289_256 ();
 b15zdnd11an1n64x5 FILLER_289_320 ();
 b15zdnd11an1n64x5 FILLER_289_384 ();
 b15zdnd11an1n64x5 FILLER_289_448 ();
 b15zdnd11an1n64x5 FILLER_289_512 ();
 b15zdnd11an1n64x5 FILLER_289_576 ();
 b15zdnd11an1n64x5 FILLER_289_640 ();
 b15zdnd11an1n64x5 FILLER_289_704 ();
 b15zdnd11an1n64x5 FILLER_289_768 ();
 b15zdnd11an1n64x5 FILLER_289_832 ();
 b15zdnd11an1n64x5 FILLER_289_896 ();
 b15zdnd11an1n64x5 FILLER_289_960 ();
 b15zdnd11an1n64x5 FILLER_289_1024 ();
 b15zdnd11an1n64x5 FILLER_289_1088 ();
 b15zdnd11an1n64x5 FILLER_289_1152 ();
 b15zdnd11an1n64x5 FILLER_289_1216 ();
 b15zdnd11an1n64x5 FILLER_289_1280 ();
 b15zdnd11an1n64x5 FILLER_289_1344 ();
 b15zdnd11an1n64x5 FILLER_289_1408 ();
 b15zdnd11an1n64x5 FILLER_289_1472 ();
 b15zdnd11an1n64x5 FILLER_289_1536 ();
 b15zdnd11an1n64x5 FILLER_289_1600 ();
 b15zdnd11an1n64x5 FILLER_289_1664 ();
 b15zdnd11an1n64x5 FILLER_289_1728 ();
 b15zdnd11an1n64x5 FILLER_289_1792 ();
 b15zdnd11an1n64x5 FILLER_289_1856 ();
 b15zdnd11an1n64x5 FILLER_289_1920 ();
 b15zdnd11an1n64x5 FILLER_289_1984 ();
 b15zdnd11an1n64x5 FILLER_289_2048 ();
 b15zdnd11an1n64x5 FILLER_289_2112 ();
 b15zdnd11an1n64x5 FILLER_289_2176 ();
 b15zdnd11an1n32x5 FILLER_289_2240 ();
 b15zdnd11an1n08x5 FILLER_289_2272 ();
 b15zdnd11an1n04x5 FILLER_289_2280 ();
 b15zdnd11an1n64x5 FILLER_290_8 ();
 b15zdnd11an1n64x5 FILLER_290_72 ();
 b15zdnd11an1n64x5 FILLER_290_136 ();
 b15zdnd11an1n64x5 FILLER_290_200 ();
 b15zdnd11an1n64x5 FILLER_290_264 ();
 b15zdnd11an1n64x5 FILLER_290_328 ();
 b15zdnd11an1n64x5 FILLER_290_392 ();
 b15zdnd11an1n64x5 FILLER_290_456 ();
 b15zdnd11an1n64x5 FILLER_290_520 ();
 b15zdnd11an1n64x5 FILLER_290_584 ();
 b15zdnd11an1n64x5 FILLER_290_648 ();
 b15zdnd11an1n04x5 FILLER_290_712 ();
 b15zdnd00an1n02x5 FILLER_290_716 ();
 b15zdnd11an1n64x5 FILLER_290_726 ();
 b15zdnd11an1n64x5 FILLER_290_790 ();
 b15zdnd11an1n64x5 FILLER_290_854 ();
 b15zdnd11an1n64x5 FILLER_290_918 ();
 b15zdnd11an1n64x5 FILLER_290_982 ();
 b15zdnd11an1n64x5 FILLER_290_1046 ();
 b15zdnd11an1n64x5 FILLER_290_1110 ();
 b15zdnd11an1n64x5 FILLER_290_1174 ();
 b15zdnd11an1n64x5 FILLER_290_1238 ();
 b15zdnd11an1n64x5 FILLER_290_1302 ();
 b15zdnd11an1n64x5 FILLER_290_1366 ();
 b15zdnd11an1n64x5 FILLER_290_1430 ();
 b15zdnd11an1n64x5 FILLER_290_1494 ();
 b15zdnd11an1n64x5 FILLER_290_1558 ();
 b15zdnd11an1n64x5 FILLER_290_1622 ();
 b15zdnd11an1n32x5 FILLER_290_1686 ();
 b15zdnd11an1n16x5 FILLER_290_1718 ();
 b15zdnd11an1n04x5 FILLER_290_1734 ();
 b15zdnd11an1n64x5 FILLER_290_1754 ();
 b15zdnd11an1n64x5 FILLER_290_1818 ();
 b15zdnd11an1n64x5 FILLER_290_1882 ();
 b15zdnd11an1n64x5 FILLER_290_1946 ();
 b15zdnd11an1n64x5 FILLER_290_2010 ();
 b15zdnd11an1n64x5 FILLER_290_2074 ();
 b15zdnd11an1n16x5 FILLER_290_2138 ();
 b15zdnd11an1n64x5 FILLER_290_2162 ();
 b15zdnd11an1n32x5 FILLER_290_2226 ();
 b15zdnd11an1n16x5 FILLER_290_2258 ();
 b15zdnd00an1n02x5 FILLER_290_2274 ();
 b15zdnd11an1n64x5 FILLER_291_0 ();
 b15zdnd11an1n64x5 FILLER_291_64 ();
 b15zdnd11an1n64x5 FILLER_291_128 ();
 b15zdnd11an1n64x5 FILLER_291_192 ();
 b15zdnd11an1n64x5 FILLER_291_256 ();
 b15zdnd11an1n64x5 FILLER_291_320 ();
 b15zdnd11an1n64x5 FILLER_291_384 ();
 b15zdnd11an1n64x5 FILLER_291_448 ();
 b15zdnd11an1n64x5 FILLER_291_512 ();
 b15zdnd11an1n64x5 FILLER_291_576 ();
 b15zdnd11an1n64x5 FILLER_291_640 ();
 b15zdnd11an1n64x5 FILLER_291_704 ();
 b15zdnd11an1n64x5 FILLER_291_768 ();
 b15zdnd11an1n64x5 FILLER_291_832 ();
 b15zdnd11an1n64x5 FILLER_291_896 ();
 b15zdnd11an1n64x5 FILLER_291_960 ();
 b15zdnd11an1n64x5 FILLER_291_1024 ();
 b15zdnd11an1n64x5 FILLER_291_1088 ();
 b15zdnd11an1n64x5 FILLER_291_1152 ();
 b15zdnd11an1n64x5 FILLER_291_1216 ();
 b15zdnd11an1n64x5 FILLER_291_1280 ();
 b15zdnd11an1n64x5 FILLER_291_1344 ();
 b15zdnd11an1n64x5 FILLER_291_1408 ();
 b15zdnd11an1n64x5 FILLER_291_1472 ();
 b15zdnd11an1n64x5 FILLER_291_1536 ();
 b15zdnd11an1n64x5 FILLER_291_1600 ();
 b15zdnd11an1n64x5 FILLER_291_1664 ();
 b15zdnd11an1n64x5 FILLER_291_1728 ();
 b15zdnd11an1n64x5 FILLER_291_1792 ();
 b15zdnd11an1n64x5 FILLER_291_1856 ();
 b15zdnd11an1n64x5 FILLER_291_1920 ();
 b15zdnd11an1n64x5 FILLER_291_1984 ();
 b15zdnd11an1n64x5 FILLER_291_2048 ();
 b15zdnd11an1n64x5 FILLER_291_2112 ();
 b15zdnd11an1n64x5 FILLER_291_2176 ();
 b15zdnd11an1n32x5 FILLER_291_2240 ();
 b15zdnd11an1n08x5 FILLER_291_2272 ();
 b15zdnd11an1n04x5 FILLER_291_2280 ();
 b15zdnd11an1n64x5 FILLER_292_8 ();
 b15zdnd11an1n64x5 FILLER_292_72 ();
 b15zdnd11an1n64x5 FILLER_292_136 ();
 b15zdnd11an1n64x5 FILLER_292_200 ();
 b15zdnd11an1n64x5 FILLER_292_264 ();
 b15zdnd11an1n64x5 FILLER_292_328 ();
 b15zdnd11an1n64x5 FILLER_292_392 ();
 b15zdnd11an1n64x5 FILLER_292_456 ();
 b15zdnd11an1n64x5 FILLER_292_520 ();
 b15zdnd11an1n64x5 FILLER_292_584 ();
 b15zdnd11an1n64x5 FILLER_292_648 ();
 b15zdnd11an1n04x5 FILLER_292_712 ();
 b15zdnd00an1n02x5 FILLER_292_716 ();
 b15zdnd11an1n64x5 FILLER_292_726 ();
 b15zdnd11an1n64x5 FILLER_292_790 ();
 b15zdnd11an1n64x5 FILLER_292_854 ();
 b15zdnd11an1n64x5 FILLER_292_918 ();
 b15zdnd11an1n64x5 FILLER_292_982 ();
 b15zdnd11an1n64x5 FILLER_292_1046 ();
 b15zdnd11an1n64x5 FILLER_292_1110 ();
 b15zdnd11an1n64x5 FILLER_292_1174 ();
 b15zdnd11an1n64x5 FILLER_292_1238 ();
 b15zdnd11an1n64x5 FILLER_292_1302 ();
 b15zdnd11an1n64x5 FILLER_292_1366 ();
 b15zdnd11an1n64x5 FILLER_292_1430 ();
 b15zdnd11an1n64x5 FILLER_292_1494 ();
 b15zdnd11an1n64x5 FILLER_292_1558 ();
 b15zdnd11an1n64x5 FILLER_292_1622 ();
 b15zdnd11an1n64x5 FILLER_292_1686 ();
 b15zdnd11an1n64x5 FILLER_292_1750 ();
 b15zdnd11an1n64x5 FILLER_292_1814 ();
 b15zdnd11an1n64x5 FILLER_292_1878 ();
 b15zdnd11an1n64x5 FILLER_292_1942 ();
 b15zdnd11an1n64x5 FILLER_292_2006 ();
 b15zdnd11an1n64x5 FILLER_292_2070 ();
 b15zdnd11an1n16x5 FILLER_292_2134 ();
 b15zdnd11an1n04x5 FILLER_292_2150 ();
 b15zdnd11an1n64x5 FILLER_292_2162 ();
 b15zdnd11an1n32x5 FILLER_292_2226 ();
 b15zdnd11an1n16x5 FILLER_292_2258 ();
 b15zdnd00an1n02x5 FILLER_292_2274 ();
 b15zdnd11an1n64x5 FILLER_293_0 ();
 b15zdnd11an1n64x5 FILLER_293_64 ();
 b15zdnd11an1n64x5 FILLER_293_128 ();
 b15zdnd11an1n64x5 FILLER_293_192 ();
 b15zdnd11an1n64x5 FILLER_293_256 ();
 b15zdnd11an1n64x5 FILLER_293_320 ();
 b15zdnd11an1n64x5 FILLER_293_384 ();
 b15zdnd11an1n64x5 FILLER_293_448 ();
 b15zdnd11an1n64x5 FILLER_293_512 ();
 b15zdnd11an1n64x5 FILLER_293_576 ();
 b15zdnd11an1n64x5 FILLER_293_640 ();
 b15zdnd11an1n64x5 FILLER_293_704 ();
 b15zdnd11an1n64x5 FILLER_293_768 ();
 b15zdnd11an1n64x5 FILLER_293_832 ();
 b15zdnd11an1n64x5 FILLER_293_896 ();
 b15zdnd11an1n64x5 FILLER_293_960 ();
 b15zdnd11an1n64x5 FILLER_293_1024 ();
 b15zdnd11an1n64x5 FILLER_293_1088 ();
 b15zdnd11an1n64x5 FILLER_293_1152 ();
 b15zdnd11an1n64x5 FILLER_293_1216 ();
 b15zdnd11an1n64x5 FILLER_293_1280 ();
 b15zdnd11an1n64x5 FILLER_293_1344 ();
 b15zdnd11an1n64x5 FILLER_293_1408 ();
 b15zdnd11an1n64x5 FILLER_293_1472 ();
 b15zdnd11an1n64x5 FILLER_293_1536 ();
 b15zdnd11an1n64x5 FILLER_293_1600 ();
 b15zdnd11an1n64x5 FILLER_293_1664 ();
 b15zdnd11an1n64x5 FILLER_293_1728 ();
 b15zdnd11an1n64x5 FILLER_293_1792 ();
 b15zdnd11an1n64x5 FILLER_293_1856 ();
 b15zdnd11an1n64x5 FILLER_293_1920 ();
 b15zdnd11an1n64x5 FILLER_293_1984 ();
 b15zdnd11an1n64x5 FILLER_293_2048 ();
 b15zdnd11an1n64x5 FILLER_293_2112 ();
 b15zdnd11an1n64x5 FILLER_293_2176 ();
 b15zdnd11an1n32x5 FILLER_293_2240 ();
 b15zdnd11an1n08x5 FILLER_293_2272 ();
 b15zdnd11an1n04x5 FILLER_293_2280 ();
 b15zdnd11an1n64x5 FILLER_294_8 ();
 b15zdnd11an1n64x5 FILLER_294_72 ();
 b15zdnd11an1n64x5 FILLER_294_136 ();
 b15zdnd11an1n64x5 FILLER_294_200 ();
 b15zdnd11an1n64x5 FILLER_294_264 ();
 b15zdnd11an1n64x5 FILLER_294_328 ();
 b15zdnd11an1n64x5 FILLER_294_392 ();
 b15zdnd11an1n64x5 FILLER_294_456 ();
 b15zdnd11an1n64x5 FILLER_294_520 ();
 b15zdnd11an1n64x5 FILLER_294_584 ();
 b15zdnd11an1n64x5 FILLER_294_648 ();
 b15zdnd11an1n04x5 FILLER_294_712 ();
 b15zdnd00an1n02x5 FILLER_294_716 ();
 b15zdnd11an1n64x5 FILLER_294_726 ();
 b15zdnd11an1n64x5 FILLER_294_790 ();
 b15zdnd11an1n64x5 FILLER_294_854 ();
 b15zdnd11an1n64x5 FILLER_294_918 ();
 b15zdnd11an1n64x5 FILLER_294_982 ();
 b15zdnd11an1n64x5 FILLER_294_1046 ();
 b15zdnd11an1n64x5 FILLER_294_1110 ();
 b15zdnd11an1n64x5 FILLER_294_1174 ();
 b15zdnd11an1n64x5 FILLER_294_1238 ();
 b15zdnd11an1n64x5 FILLER_294_1302 ();
 b15zdnd11an1n64x5 FILLER_294_1366 ();
 b15zdnd11an1n64x5 FILLER_294_1430 ();
 b15zdnd11an1n64x5 FILLER_294_1494 ();
 b15zdnd11an1n64x5 FILLER_294_1558 ();
 b15zdnd11an1n64x5 FILLER_294_1622 ();
 b15zdnd11an1n64x5 FILLER_294_1686 ();
 b15zdnd11an1n64x5 FILLER_294_1750 ();
 b15zdnd11an1n64x5 FILLER_294_1814 ();
 b15zdnd11an1n64x5 FILLER_294_1878 ();
 b15zdnd11an1n64x5 FILLER_294_1942 ();
 b15zdnd11an1n64x5 FILLER_294_2006 ();
 b15zdnd11an1n64x5 FILLER_294_2070 ();
 b15zdnd11an1n16x5 FILLER_294_2134 ();
 b15zdnd11an1n04x5 FILLER_294_2150 ();
 b15zdnd11an1n64x5 FILLER_294_2162 ();
 b15zdnd11an1n32x5 FILLER_294_2226 ();
 b15zdnd11an1n16x5 FILLER_294_2258 ();
 b15zdnd00an1n02x5 FILLER_294_2274 ();
 b15zdnd11an1n64x5 FILLER_295_0 ();
 b15zdnd11an1n64x5 FILLER_295_64 ();
 b15zdnd11an1n64x5 FILLER_295_128 ();
 b15zdnd11an1n64x5 FILLER_295_192 ();
 b15zdnd11an1n64x5 FILLER_295_256 ();
 b15zdnd11an1n64x5 FILLER_295_320 ();
 b15zdnd11an1n64x5 FILLER_295_384 ();
 b15zdnd11an1n64x5 FILLER_295_448 ();
 b15zdnd11an1n64x5 FILLER_295_512 ();
 b15zdnd11an1n64x5 FILLER_295_576 ();
 b15zdnd11an1n64x5 FILLER_295_640 ();
 b15zdnd11an1n64x5 FILLER_295_704 ();
 b15zdnd11an1n64x5 FILLER_295_768 ();
 b15zdnd11an1n64x5 FILLER_295_832 ();
 b15zdnd11an1n64x5 FILLER_295_896 ();
 b15zdnd11an1n64x5 FILLER_295_960 ();
 b15zdnd11an1n64x5 FILLER_295_1024 ();
 b15zdnd11an1n64x5 FILLER_295_1088 ();
 b15zdnd11an1n64x5 FILLER_295_1152 ();
 b15zdnd11an1n64x5 FILLER_295_1216 ();
 b15zdnd11an1n64x5 FILLER_295_1280 ();
 b15zdnd11an1n64x5 FILLER_295_1344 ();
 b15zdnd11an1n64x5 FILLER_295_1408 ();
 b15zdnd11an1n64x5 FILLER_295_1472 ();
 b15zdnd11an1n64x5 FILLER_295_1536 ();
 b15zdnd11an1n64x5 FILLER_295_1600 ();
 b15zdnd11an1n64x5 FILLER_295_1664 ();
 b15zdnd11an1n64x5 FILLER_295_1728 ();
 b15zdnd11an1n64x5 FILLER_295_1792 ();
 b15zdnd11an1n64x5 FILLER_295_1856 ();
 b15zdnd11an1n64x5 FILLER_295_1920 ();
 b15zdnd11an1n64x5 FILLER_295_1984 ();
 b15zdnd11an1n64x5 FILLER_295_2048 ();
 b15zdnd11an1n64x5 FILLER_295_2112 ();
 b15zdnd11an1n64x5 FILLER_295_2176 ();
 b15zdnd11an1n32x5 FILLER_295_2240 ();
 b15zdnd11an1n08x5 FILLER_295_2272 ();
 b15zdnd11an1n04x5 FILLER_295_2280 ();
 b15zdnd11an1n64x5 FILLER_296_8 ();
 b15zdnd11an1n64x5 FILLER_296_72 ();
 b15zdnd11an1n64x5 FILLER_296_136 ();
 b15zdnd11an1n64x5 FILLER_296_200 ();
 b15zdnd11an1n64x5 FILLER_296_264 ();
 b15zdnd11an1n64x5 FILLER_296_328 ();
 b15zdnd11an1n64x5 FILLER_296_392 ();
 b15zdnd11an1n64x5 FILLER_296_456 ();
 b15zdnd11an1n64x5 FILLER_296_520 ();
 b15zdnd11an1n64x5 FILLER_296_584 ();
 b15zdnd11an1n64x5 FILLER_296_648 ();
 b15zdnd11an1n04x5 FILLER_296_712 ();
 b15zdnd00an1n02x5 FILLER_296_716 ();
 b15zdnd11an1n64x5 FILLER_296_726 ();
 b15zdnd11an1n64x5 FILLER_296_790 ();
 b15zdnd11an1n64x5 FILLER_296_854 ();
 b15zdnd11an1n64x5 FILLER_296_918 ();
 b15zdnd11an1n64x5 FILLER_296_982 ();
 b15zdnd11an1n64x5 FILLER_296_1046 ();
 b15zdnd11an1n64x5 FILLER_296_1110 ();
 b15zdnd11an1n64x5 FILLER_296_1174 ();
 b15zdnd11an1n64x5 FILLER_296_1238 ();
 b15zdnd11an1n64x5 FILLER_296_1302 ();
 b15zdnd11an1n64x5 FILLER_296_1366 ();
 b15zdnd11an1n64x5 FILLER_296_1430 ();
 b15zdnd11an1n64x5 FILLER_296_1494 ();
 b15zdnd11an1n64x5 FILLER_296_1558 ();
 b15zdnd11an1n64x5 FILLER_296_1622 ();
 b15zdnd11an1n64x5 FILLER_296_1686 ();
 b15zdnd11an1n64x5 FILLER_296_1750 ();
 b15zdnd11an1n64x5 FILLER_296_1814 ();
 b15zdnd11an1n64x5 FILLER_296_1878 ();
 b15zdnd11an1n64x5 FILLER_296_1942 ();
 b15zdnd11an1n64x5 FILLER_296_2006 ();
 b15zdnd11an1n64x5 FILLER_296_2070 ();
 b15zdnd11an1n16x5 FILLER_296_2134 ();
 b15zdnd11an1n04x5 FILLER_296_2150 ();
 b15zdnd11an1n64x5 FILLER_296_2162 ();
 b15zdnd11an1n32x5 FILLER_296_2226 ();
 b15zdnd11an1n16x5 FILLER_296_2258 ();
 b15zdnd00an1n02x5 FILLER_296_2274 ();
 b15zdnd11an1n64x5 FILLER_297_0 ();
 b15zdnd11an1n64x5 FILLER_297_64 ();
 b15zdnd11an1n64x5 FILLER_297_128 ();
 b15zdnd11an1n64x5 FILLER_297_192 ();
 b15zdnd11an1n64x5 FILLER_297_256 ();
 b15zdnd11an1n64x5 FILLER_297_320 ();
 b15zdnd11an1n64x5 FILLER_297_384 ();
 b15zdnd11an1n64x5 FILLER_297_448 ();
 b15zdnd11an1n64x5 FILLER_297_512 ();
 b15zdnd11an1n64x5 FILLER_297_576 ();
 b15zdnd11an1n64x5 FILLER_297_640 ();
 b15zdnd11an1n64x5 FILLER_297_704 ();
 b15zdnd11an1n64x5 FILLER_297_768 ();
 b15zdnd11an1n64x5 FILLER_297_832 ();
 b15zdnd11an1n64x5 FILLER_297_896 ();
 b15zdnd11an1n64x5 FILLER_297_960 ();
 b15zdnd11an1n64x5 FILLER_297_1024 ();
 b15zdnd11an1n64x5 FILLER_297_1088 ();
 b15zdnd11an1n64x5 FILLER_297_1152 ();
 b15zdnd11an1n64x5 FILLER_297_1216 ();
 b15zdnd11an1n64x5 FILLER_297_1280 ();
 b15zdnd11an1n64x5 FILLER_297_1344 ();
 b15zdnd11an1n64x5 FILLER_297_1408 ();
 b15zdnd11an1n64x5 FILLER_297_1472 ();
 b15zdnd11an1n64x5 FILLER_297_1536 ();
 b15zdnd11an1n64x5 FILLER_297_1600 ();
 b15zdnd11an1n64x5 FILLER_297_1664 ();
 b15zdnd11an1n64x5 FILLER_297_1728 ();
 b15zdnd11an1n64x5 FILLER_297_1792 ();
 b15zdnd11an1n64x5 FILLER_297_1856 ();
 b15zdnd11an1n64x5 FILLER_297_1920 ();
 b15zdnd11an1n64x5 FILLER_297_1984 ();
 b15zdnd11an1n64x5 FILLER_297_2048 ();
 b15zdnd11an1n64x5 FILLER_297_2112 ();
 b15zdnd11an1n64x5 FILLER_297_2176 ();
 b15zdnd11an1n32x5 FILLER_297_2240 ();
 b15zdnd11an1n08x5 FILLER_297_2272 ();
 b15zdnd11an1n04x5 FILLER_297_2280 ();
 b15zdnd11an1n64x5 FILLER_298_8 ();
 b15zdnd11an1n64x5 FILLER_298_72 ();
 b15zdnd11an1n64x5 FILLER_298_136 ();
 b15zdnd11an1n64x5 FILLER_298_200 ();
 b15zdnd11an1n64x5 FILLER_298_264 ();
 b15zdnd11an1n64x5 FILLER_298_328 ();
 b15zdnd11an1n64x5 FILLER_298_392 ();
 b15zdnd11an1n64x5 FILLER_298_456 ();
 b15zdnd11an1n64x5 FILLER_298_520 ();
 b15zdnd11an1n64x5 FILLER_298_584 ();
 b15zdnd11an1n64x5 FILLER_298_648 ();
 b15zdnd11an1n04x5 FILLER_298_712 ();
 b15zdnd00an1n02x5 FILLER_298_716 ();
 b15zdnd11an1n64x5 FILLER_298_726 ();
 b15zdnd11an1n64x5 FILLER_298_790 ();
 b15zdnd11an1n64x5 FILLER_298_854 ();
 b15zdnd11an1n64x5 FILLER_298_918 ();
 b15zdnd11an1n64x5 FILLER_298_982 ();
 b15zdnd11an1n64x5 FILLER_298_1046 ();
 b15zdnd11an1n64x5 FILLER_298_1110 ();
 b15zdnd11an1n64x5 FILLER_298_1174 ();
 b15zdnd11an1n64x5 FILLER_298_1238 ();
 b15zdnd11an1n64x5 FILLER_298_1302 ();
 b15zdnd11an1n64x5 FILLER_298_1366 ();
 b15zdnd11an1n64x5 FILLER_298_1430 ();
 b15zdnd11an1n64x5 FILLER_298_1494 ();
 b15zdnd11an1n64x5 FILLER_298_1558 ();
 b15zdnd11an1n64x5 FILLER_298_1622 ();
 b15zdnd11an1n64x5 FILLER_298_1686 ();
 b15zdnd11an1n64x5 FILLER_298_1750 ();
 b15zdnd11an1n64x5 FILLER_298_1814 ();
 b15zdnd11an1n64x5 FILLER_298_1878 ();
 b15zdnd11an1n64x5 FILLER_298_1942 ();
 b15zdnd11an1n64x5 FILLER_298_2006 ();
 b15zdnd11an1n64x5 FILLER_298_2070 ();
 b15zdnd11an1n16x5 FILLER_298_2134 ();
 b15zdnd11an1n04x5 FILLER_298_2150 ();
 b15zdnd11an1n64x5 FILLER_298_2162 ();
 b15zdnd11an1n32x5 FILLER_298_2226 ();
 b15zdnd11an1n16x5 FILLER_298_2258 ();
 b15zdnd00an1n02x5 FILLER_298_2274 ();
 b15zdnd11an1n64x5 FILLER_299_0 ();
 b15zdnd11an1n64x5 FILLER_299_64 ();
 b15zdnd11an1n64x5 FILLER_299_128 ();
 b15zdnd11an1n64x5 FILLER_299_192 ();
 b15zdnd11an1n64x5 FILLER_299_256 ();
 b15zdnd11an1n64x5 FILLER_299_320 ();
 b15zdnd11an1n64x5 FILLER_299_384 ();
 b15zdnd11an1n64x5 FILLER_299_448 ();
 b15zdnd11an1n64x5 FILLER_299_512 ();
 b15zdnd11an1n64x5 FILLER_299_576 ();
 b15zdnd11an1n64x5 FILLER_299_640 ();
 b15zdnd11an1n64x5 FILLER_299_704 ();
 b15zdnd11an1n64x5 FILLER_299_768 ();
 b15zdnd11an1n64x5 FILLER_299_832 ();
 b15zdnd11an1n64x5 FILLER_299_896 ();
 b15zdnd11an1n64x5 FILLER_299_960 ();
 b15zdnd11an1n64x5 FILLER_299_1024 ();
 b15zdnd11an1n64x5 FILLER_299_1088 ();
 b15zdnd11an1n64x5 FILLER_299_1152 ();
 b15zdnd11an1n64x5 FILLER_299_1216 ();
 b15zdnd11an1n64x5 FILLER_299_1280 ();
 b15zdnd11an1n64x5 FILLER_299_1344 ();
 b15zdnd11an1n32x5 FILLER_299_1408 ();
 b15zdnd11an1n16x5 FILLER_299_1440 ();
 b15zdnd11an1n08x5 FILLER_299_1456 ();
 b15zdnd00an1n02x5 FILLER_299_1464 ();
 b15zdnd00an1n01x5 FILLER_299_1466 ();
 b15zdnd11an1n64x5 FILLER_299_1483 ();
 b15zdnd11an1n64x5 FILLER_299_1547 ();
 b15zdnd11an1n64x5 FILLER_299_1611 ();
 b15zdnd11an1n64x5 FILLER_299_1675 ();
 b15zdnd11an1n64x5 FILLER_299_1739 ();
 b15zdnd11an1n64x5 FILLER_299_1803 ();
 b15zdnd11an1n64x5 FILLER_299_1867 ();
 b15zdnd11an1n64x5 FILLER_299_1931 ();
 b15zdnd11an1n64x5 FILLER_299_1995 ();
 b15zdnd11an1n64x5 FILLER_299_2059 ();
 b15zdnd11an1n64x5 FILLER_299_2123 ();
 b15zdnd11an1n64x5 FILLER_299_2187 ();
 b15zdnd11an1n32x5 FILLER_299_2251 ();
 b15zdnd00an1n01x5 FILLER_299_2283 ();
 b15zdnd11an1n64x5 FILLER_300_8 ();
 b15zdnd11an1n64x5 FILLER_300_72 ();
 b15zdnd11an1n64x5 FILLER_300_136 ();
 b15zdnd11an1n64x5 FILLER_300_200 ();
 b15zdnd11an1n64x5 FILLER_300_264 ();
 b15zdnd11an1n64x5 FILLER_300_328 ();
 b15zdnd11an1n64x5 FILLER_300_392 ();
 b15zdnd11an1n64x5 FILLER_300_456 ();
 b15zdnd11an1n64x5 FILLER_300_520 ();
 b15zdnd11an1n64x5 FILLER_300_584 ();
 b15zdnd11an1n64x5 FILLER_300_648 ();
 b15zdnd11an1n04x5 FILLER_300_712 ();
 b15zdnd00an1n02x5 FILLER_300_716 ();
 b15zdnd11an1n64x5 FILLER_300_726 ();
 b15zdnd11an1n64x5 FILLER_300_790 ();
 b15zdnd11an1n64x5 FILLER_300_854 ();
 b15zdnd11an1n64x5 FILLER_300_918 ();
 b15zdnd11an1n64x5 FILLER_300_982 ();
 b15zdnd11an1n64x5 FILLER_300_1046 ();
 b15zdnd11an1n64x5 FILLER_300_1110 ();
 b15zdnd11an1n64x5 FILLER_300_1174 ();
 b15zdnd11an1n64x5 FILLER_300_1238 ();
 b15zdnd11an1n64x5 FILLER_300_1302 ();
 b15zdnd11an1n64x5 FILLER_300_1366 ();
 b15zdnd11an1n64x5 FILLER_300_1430 ();
 b15zdnd11an1n64x5 FILLER_300_1494 ();
 b15zdnd11an1n64x5 FILLER_300_1558 ();
 b15zdnd11an1n64x5 FILLER_300_1622 ();
 b15zdnd11an1n64x5 FILLER_300_1686 ();
 b15zdnd11an1n64x5 FILLER_300_1750 ();
 b15zdnd11an1n64x5 FILLER_300_1814 ();
 b15zdnd11an1n64x5 FILLER_300_1878 ();
 b15zdnd11an1n64x5 FILLER_300_1942 ();
 b15zdnd11an1n64x5 FILLER_300_2006 ();
 b15zdnd11an1n64x5 FILLER_300_2070 ();
 b15zdnd11an1n16x5 FILLER_300_2134 ();
 b15zdnd11an1n04x5 FILLER_300_2150 ();
 b15zdnd11an1n64x5 FILLER_300_2162 ();
 b15zdnd11an1n32x5 FILLER_300_2226 ();
 b15zdnd11an1n16x5 FILLER_300_2258 ();
 b15zdnd00an1n02x5 FILLER_300_2274 ();
 b15zdnd11an1n64x5 FILLER_301_0 ();
 b15zdnd11an1n64x5 FILLER_301_64 ();
 b15zdnd11an1n64x5 FILLER_301_128 ();
 b15zdnd11an1n64x5 FILLER_301_192 ();
 b15zdnd11an1n64x5 FILLER_301_256 ();
 b15zdnd11an1n64x5 FILLER_301_320 ();
 b15zdnd11an1n64x5 FILLER_301_384 ();
 b15zdnd11an1n64x5 FILLER_301_448 ();
 b15zdnd11an1n64x5 FILLER_301_512 ();
 b15zdnd11an1n64x5 FILLER_301_576 ();
 b15zdnd11an1n64x5 FILLER_301_640 ();
 b15zdnd11an1n64x5 FILLER_301_704 ();
 b15zdnd11an1n64x5 FILLER_301_768 ();
 b15zdnd11an1n64x5 FILLER_301_832 ();
 b15zdnd11an1n64x5 FILLER_301_896 ();
 b15zdnd11an1n64x5 FILLER_301_960 ();
 b15zdnd11an1n64x5 FILLER_301_1024 ();
 b15zdnd11an1n64x5 FILLER_301_1088 ();
 b15zdnd11an1n64x5 FILLER_301_1152 ();
 b15zdnd11an1n64x5 FILLER_301_1216 ();
 b15zdnd11an1n64x5 FILLER_301_1280 ();
 b15zdnd11an1n64x5 FILLER_301_1344 ();
 b15zdnd11an1n64x5 FILLER_301_1408 ();
 b15zdnd11an1n64x5 FILLER_301_1472 ();
 b15zdnd11an1n64x5 FILLER_301_1536 ();
 b15zdnd11an1n64x5 FILLER_301_1600 ();
 b15zdnd11an1n64x5 FILLER_301_1664 ();
 b15zdnd11an1n64x5 FILLER_301_1728 ();
 b15zdnd11an1n64x5 FILLER_301_1792 ();
 b15zdnd11an1n64x5 FILLER_301_1856 ();
 b15zdnd11an1n64x5 FILLER_301_1920 ();
 b15zdnd11an1n64x5 FILLER_301_1984 ();
 b15zdnd11an1n64x5 FILLER_301_2048 ();
 b15zdnd11an1n64x5 FILLER_301_2112 ();
 b15zdnd11an1n64x5 FILLER_301_2176 ();
 b15zdnd11an1n32x5 FILLER_301_2240 ();
 b15zdnd11an1n08x5 FILLER_301_2272 ();
 b15zdnd11an1n04x5 FILLER_301_2280 ();
 b15zdnd11an1n64x5 FILLER_302_8 ();
 b15zdnd11an1n64x5 FILLER_302_72 ();
 b15zdnd11an1n64x5 FILLER_302_136 ();
 b15zdnd11an1n64x5 FILLER_302_200 ();
 b15zdnd11an1n64x5 FILLER_302_264 ();
 b15zdnd11an1n64x5 FILLER_302_328 ();
 b15zdnd11an1n64x5 FILLER_302_392 ();
 b15zdnd11an1n64x5 FILLER_302_456 ();
 b15zdnd11an1n64x5 FILLER_302_520 ();
 b15zdnd11an1n64x5 FILLER_302_584 ();
 b15zdnd11an1n64x5 FILLER_302_648 ();
 b15zdnd11an1n04x5 FILLER_302_712 ();
 b15zdnd00an1n02x5 FILLER_302_716 ();
 b15zdnd11an1n64x5 FILLER_302_726 ();
 b15zdnd11an1n64x5 FILLER_302_790 ();
 b15zdnd11an1n64x5 FILLER_302_854 ();
 b15zdnd11an1n32x5 FILLER_302_918 ();
 b15zdnd11an1n08x5 FILLER_302_950 ();
 b15zdnd00an1n02x5 FILLER_302_958 ();
 b15zdnd00an1n01x5 FILLER_302_960 ();
 b15zdnd11an1n64x5 FILLER_302_1003 ();
 b15zdnd11an1n64x5 FILLER_302_1067 ();
 b15zdnd11an1n64x5 FILLER_302_1131 ();
 b15zdnd11an1n64x5 FILLER_302_1195 ();
 b15zdnd11an1n64x5 FILLER_302_1259 ();
 b15zdnd11an1n64x5 FILLER_302_1323 ();
 b15zdnd11an1n64x5 FILLER_302_1387 ();
 b15zdnd11an1n64x5 FILLER_302_1451 ();
 b15zdnd11an1n64x5 FILLER_302_1515 ();
 b15zdnd11an1n64x5 FILLER_302_1579 ();
 b15zdnd11an1n64x5 FILLER_302_1643 ();
 b15zdnd11an1n64x5 FILLER_302_1707 ();
 b15zdnd11an1n64x5 FILLER_302_1771 ();
 b15zdnd11an1n64x5 FILLER_302_1835 ();
 b15zdnd11an1n64x5 FILLER_302_1899 ();
 b15zdnd11an1n64x5 FILLER_302_1963 ();
 b15zdnd11an1n64x5 FILLER_302_2027 ();
 b15zdnd11an1n32x5 FILLER_302_2091 ();
 b15zdnd11an1n16x5 FILLER_302_2123 ();
 b15zdnd11an1n08x5 FILLER_302_2139 ();
 b15zdnd11an1n04x5 FILLER_302_2147 ();
 b15zdnd00an1n02x5 FILLER_302_2151 ();
 b15zdnd00an1n01x5 FILLER_302_2153 ();
 b15zdnd11an1n64x5 FILLER_302_2162 ();
 b15zdnd11an1n32x5 FILLER_302_2226 ();
 b15zdnd11an1n16x5 FILLER_302_2258 ();
 b15zdnd00an1n02x5 FILLER_302_2274 ();
 b15zdnd11an1n64x5 FILLER_303_0 ();
 b15zdnd11an1n64x5 FILLER_303_64 ();
 b15zdnd11an1n64x5 FILLER_303_128 ();
 b15zdnd11an1n64x5 FILLER_303_192 ();
 b15zdnd11an1n64x5 FILLER_303_256 ();
 b15zdnd11an1n64x5 FILLER_303_320 ();
 b15zdnd11an1n64x5 FILLER_303_384 ();
 b15zdnd11an1n64x5 FILLER_303_448 ();
 b15zdnd11an1n64x5 FILLER_303_512 ();
 b15zdnd11an1n64x5 FILLER_303_576 ();
 b15zdnd11an1n64x5 FILLER_303_640 ();
 b15zdnd11an1n64x5 FILLER_303_704 ();
 b15zdnd11an1n64x5 FILLER_303_768 ();
 b15zdnd11an1n64x5 FILLER_303_832 ();
 b15zdnd11an1n64x5 FILLER_303_896 ();
 b15zdnd11an1n04x5 FILLER_303_960 ();
 b15zdnd00an1n02x5 FILLER_303_964 ();
 b15zdnd11an1n64x5 FILLER_303_1008 ();
 b15zdnd11an1n64x5 FILLER_303_1072 ();
 b15zdnd11an1n64x5 FILLER_303_1136 ();
 b15zdnd11an1n64x5 FILLER_303_1200 ();
 b15zdnd11an1n64x5 FILLER_303_1264 ();
 b15zdnd11an1n64x5 FILLER_303_1328 ();
 b15zdnd11an1n64x5 FILLER_303_1392 ();
 b15zdnd11an1n64x5 FILLER_303_1456 ();
 b15zdnd11an1n64x5 FILLER_303_1520 ();
 b15zdnd11an1n64x5 FILLER_303_1584 ();
 b15zdnd11an1n64x5 FILLER_303_1648 ();
 b15zdnd11an1n64x5 FILLER_303_1712 ();
 b15zdnd11an1n64x5 FILLER_303_1776 ();
 b15zdnd11an1n64x5 FILLER_303_1840 ();
 b15zdnd11an1n64x5 FILLER_303_1904 ();
 b15zdnd11an1n64x5 FILLER_303_1968 ();
 b15zdnd11an1n64x5 FILLER_303_2032 ();
 b15zdnd11an1n64x5 FILLER_303_2096 ();
 b15zdnd11an1n64x5 FILLER_303_2160 ();
 b15zdnd11an1n32x5 FILLER_303_2224 ();
 b15zdnd11an1n16x5 FILLER_303_2256 ();
 b15zdnd11an1n08x5 FILLER_303_2272 ();
 b15zdnd11an1n04x5 FILLER_303_2280 ();
 b15zdnd11an1n64x5 FILLER_304_8 ();
 b15zdnd11an1n64x5 FILLER_304_72 ();
 b15zdnd11an1n64x5 FILLER_304_136 ();
 b15zdnd11an1n64x5 FILLER_304_200 ();
 b15zdnd11an1n64x5 FILLER_304_264 ();
 b15zdnd11an1n64x5 FILLER_304_328 ();
 b15zdnd11an1n64x5 FILLER_304_392 ();
 b15zdnd11an1n64x5 FILLER_304_456 ();
 b15zdnd11an1n64x5 FILLER_304_520 ();
 b15zdnd11an1n64x5 FILLER_304_584 ();
 b15zdnd11an1n64x5 FILLER_304_648 ();
 b15zdnd11an1n04x5 FILLER_304_712 ();
 b15zdnd00an1n02x5 FILLER_304_716 ();
 b15zdnd11an1n64x5 FILLER_304_726 ();
 b15zdnd11an1n64x5 FILLER_304_790 ();
 b15zdnd11an1n64x5 FILLER_304_854 ();
 b15zdnd11an1n32x5 FILLER_304_918 ();
 b15zdnd11an1n16x5 FILLER_304_950 ();
 b15zdnd11an1n04x5 FILLER_304_966 ();
 b15zdnd00an1n01x5 FILLER_304_970 ();
 b15zdnd11an1n64x5 FILLER_304_1013 ();
 b15zdnd11an1n64x5 FILLER_304_1077 ();
 b15zdnd11an1n64x5 FILLER_304_1141 ();
 b15zdnd11an1n64x5 FILLER_304_1205 ();
 b15zdnd11an1n64x5 FILLER_304_1269 ();
 b15zdnd11an1n64x5 FILLER_304_1333 ();
 b15zdnd11an1n64x5 FILLER_304_1397 ();
 b15zdnd11an1n64x5 FILLER_304_1461 ();
 b15zdnd11an1n64x5 FILLER_304_1525 ();
 b15zdnd11an1n64x5 FILLER_304_1589 ();
 b15zdnd11an1n64x5 FILLER_304_1653 ();
 b15zdnd11an1n64x5 FILLER_304_1717 ();
 b15zdnd11an1n08x5 FILLER_304_1781 ();
 b15zdnd11an1n04x5 FILLER_304_1789 ();
 b15zdnd00an1n02x5 FILLER_304_1793 ();
 b15zdnd11an1n64x5 FILLER_304_1811 ();
 b15zdnd11an1n64x5 FILLER_304_1875 ();
 b15zdnd11an1n64x5 FILLER_304_1939 ();
 b15zdnd11an1n64x5 FILLER_304_2003 ();
 b15zdnd11an1n64x5 FILLER_304_2067 ();
 b15zdnd11an1n16x5 FILLER_304_2131 ();
 b15zdnd11an1n04x5 FILLER_304_2147 ();
 b15zdnd00an1n02x5 FILLER_304_2151 ();
 b15zdnd00an1n01x5 FILLER_304_2153 ();
 b15zdnd11an1n64x5 FILLER_304_2162 ();
 b15zdnd11an1n32x5 FILLER_304_2226 ();
 b15zdnd11an1n16x5 FILLER_304_2258 ();
 b15zdnd00an1n02x5 FILLER_304_2274 ();
 b15zdnd11an1n64x5 FILLER_305_0 ();
 b15zdnd11an1n64x5 FILLER_305_64 ();
 b15zdnd11an1n64x5 FILLER_305_128 ();
 b15zdnd11an1n64x5 FILLER_305_192 ();
 b15zdnd11an1n64x5 FILLER_305_256 ();
 b15zdnd11an1n64x5 FILLER_305_320 ();
 b15zdnd11an1n64x5 FILLER_305_384 ();
 b15zdnd11an1n64x5 FILLER_305_448 ();
 b15zdnd11an1n64x5 FILLER_305_512 ();
 b15zdnd11an1n64x5 FILLER_305_576 ();
 b15zdnd11an1n64x5 FILLER_305_640 ();
 b15zdnd11an1n64x5 FILLER_305_704 ();
 b15zdnd11an1n64x5 FILLER_305_768 ();
 b15zdnd11an1n64x5 FILLER_305_832 ();
 b15zdnd11an1n64x5 FILLER_305_896 ();
 b15zdnd11an1n64x5 FILLER_305_960 ();
 b15zdnd11an1n64x5 FILLER_305_1024 ();
 b15zdnd11an1n64x5 FILLER_305_1088 ();
 b15zdnd11an1n64x5 FILLER_305_1152 ();
 b15zdnd11an1n64x5 FILLER_305_1216 ();
 b15zdnd11an1n64x5 FILLER_305_1280 ();
 b15zdnd11an1n64x5 FILLER_305_1344 ();
 b15zdnd11an1n64x5 FILLER_305_1408 ();
 b15zdnd11an1n32x5 FILLER_305_1472 ();
 b15zdnd11an1n04x5 FILLER_305_1504 ();
 b15zdnd00an1n02x5 FILLER_305_1508 ();
 b15zdnd00an1n01x5 FILLER_305_1510 ();
 b15zdnd11an1n64x5 FILLER_305_1527 ();
 b15zdnd11an1n64x5 FILLER_305_1591 ();
 b15zdnd11an1n64x5 FILLER_305_1655 ();
 b15zdnd11an1n64x5 FILLER_305_1719 ();
 b15zdnd11an1n64x5 FILLER_305_1783 ();
 b15zdnd11an1n64x5 FILLER_305_1847 ();
 b15zdnd11an1n64x5 FILLER_305_1911 ();
 b15zdnd11an1n64x5 FILLER_305_1975 ();
 b15zdnd11an1n64x5 FILLER_305_2039 ();
 b15zdnd11an1n64x5 FILLER_305_2103 ();
 b15zdnd11an1n64x5 FILLER_305_2167 ();
 b15zdnd11an1n32x5 FILLER_305_2231 ();
 b15zdnd11an1n16x5 FILLER_305_2263 ();
 b15zdnd11an1n04x5 FILLER_305_2279 ();
 b15zdnd00an1n01x5 FILLER_305_2283 ();
 b15zdnd11an1n64x5 FILLER_306_8 ();
 b15zdnd11an1n64x5 FILLER_306_72 ();
 b15zdnd11an1n64x5 FILLER_306_136 ();
 b15zdnd11an1n64x5 FILLER_306_200 ();
 b15zdnd11an1n64x5 FILLER_306_264 ();
 b15zdnd11an1n64x5 FILLER_306_328 ();
 b15zdnd11an1n64x5 FILLER_306_392 ();
 b15zdnd11an1n64x5 FILLER_306_456 ();
 b15zdnd11an1n64x5 FILLER_306_520 ();
 b15zdnd11an1n64x5 FILLER_306_584 ();
 b15zdnd11an1n64x5 FILLER_306_648 ();
 b15zdnd11an1n04x5 FILLER_306_712 ();
 b15zdnd00an1n02x5 FILLER_306_716 ();
 b15zdnd11an1n64x5 FILLER_306_726 ();
 b15zdnd11an1n64x5 FILLER_306_790 ();
 b15zdnd11an1n64x5 FILLER_306_854 ();
 b15zdnd11an1n64x5 FILLER_306_918 ();
 b15zdnd11an1n64x5 FILLER_306_982 ();
 b15zdnd11an1n64x5 FILLER_306_1046 ();
 b15zdnd11an1n64x5 FILLER_306_1110 ();
 b15zdnd11an1n64x5 FILLER_306_1174 ();
 b15zdnd11an1n64x5 FILLER_306_1238 ();
 b15zdnd11an1n64x5 FILLER_306_1302 ();
 b15zdnd11an1n64x5 FILLER_306_1366 ();
 b15zdnd11an1n64x5 FILLER_306_1430 ();
 b15zdnd11an1n64x5 FILLER_306_1494 ();
 b15zdnd11an1n64x5 FILLER_306_1558 ();
 b15zdnd11an1n64x5 FILLER_306_1622 ();
 b15zdnd11an1n64x5 FILLER_306_1686 ();
 b15zdnd11an1n64x5 FILLER_306_1750 ();
 b15zdnd11an1n64x5 FILLER_306_1814 ();
 b15zdnd11an1n64x5 FILLER_306_1878 ();
 b15zdnd11an1n64x5 FILLER_306_1942 ();
 b15zdnd11an1n64x5 FILLER_306_2006 ();
 b15zdnd11an1n64x5 FILLER_306_2070 ();
 b15zdnd11an1n16x5 FILLER_306_2134 ();
 b15zdnd11an1n04x5 FILLER_306_2150 ();
 b15zdnd11an1n64x5 FILLER_306_2162 ();
 b15zdnd11an1n32x5 FILLER_306_2226 ();
 b15zdnd11an1n16x5 FILLER_306_2258 ();
 b15zdnd00an1n02x5 FILLER_306_2274 ();
 b15zdnd11an1n64x5 FILLER_307_0 ();
 b15zdnd11an1n64x5 FILLER_307_64 ();
 b15zdnd11an1n64x5 FILLER_307_128 ();
 b15zdnd11an1n64x5 FILLER_307_192 ();
 b15zdnd11an1n64x5 FILLER_307_256 ();
 b15zdnd11an1n64x5 FILLER_307_320 ();
 b15zdnd11an1n64x5 FILLER_307_384 ();
 b15zdnd11an1n64x5 FILLER_307_448 ();
 b15zdnd11an1n64x5 FILLER_307_512 ();
 b15zdnd11an1n64x5 FILLER_307_576 ();
 b15zdnd11an1n64x5 FILLER_307_640 ();
 b15zdnd11an1n64x5 FILLER_307_704 ();
 b15zdnd11an1n64x5 FILLER_307_768 ();
 b15zdnd11an1n64x5 FILLER_307_832 ();
 b15zdnd11an1n64x5 FILLER_307_896 ();
 b15zdnd11an1n64x5 FILLER_307_960 ();
 b15zdnd11an1n64x5 FILLER_307_1024 ();
 b15zdnd11an1n64x5 FILLER_307_1088 ();
 b15zdnd11an1n64x5 FILLER_307_1152 ();
 b15zdnd11an1n64x5 FILLER_307_1216 ();
 b15zdnd11an1n64x5 FILLER_307_1280 ();
 b15zdnd11an1n64x5 FILLER_307_1344 ();
 b15zdnd11an1n64x5 FILLER_307_1408 ();
 b15zdnd11an1n64x5 FILLER_307_1472 ();
 b15zdnd11an1n64x5 FILLER_307_1536 ();
 b15zdnd11an1n64x5 FILLER_307_1600 ();
 b15zdnd11an1n64x5 FILLER_307_1664 ();
 b15zdnd11an1n64x5 FILLER_307_1728 ();
 b15zdnd11an1n64x5 FILLER_307_1792 ();
 b15zdnd11an1n64x5 FILLER_307_1856 ();
 b15zdnd11an1n64x5 FILLER_307_1920 ();
 b15zdnd11an1n64x5 FILLER_307_1984 ();
 b15zdnd11an1n64x5 FILLER_307_2048 ();
 b15zdnd11an1n64x5 FILLER_307_2112 ();
 b15zdnd11an1n64x5 FILLER_307_2176 ();
 b15zdnd11an1n32x5 FILLER_307_2240 ();
 b15zdnd11an1n08x5 FILLER_307_2272 ();
 b15zdnd11an1n04x5 FILLER_307_2280 ();
 b15zdnd11an1n64x5 FILLER_308_8 ();
 b15zdnd11an1n64x5 FILLER_308_72 ();
 b15zdnd11an1n64x5 FILLER_308_136 ();
 b15zdnd11an1n64x5 FILLER_308_200 ();
 b15zdnd11an1n64x5 FILLER_308_264 ();
 b15zdnd11an1n64x5 FILLER_308_328 ();
 b15zdnd11an1n64x5 FILLER_308_392 ();
 b15zdnd11an1n64x5 FILLER_308_456 ();
 b15zdnd11an1n64x5 FILLER_308_520 ();
 b15zdnd11an1n64x5 FILLER_308_584 ();
 b15zdnd11an1n64x5 FILLER_308_648 ();
 b15zdnd11an1n04x5 FILLER_308_712 ();
 b15zdnd00an1n02x5 FILLER_308_716 ();
 b15zdnd11an1n64x5 FILLER_308_726 ();
 b15zdnd11an1n64x5 FILLER_308_790 ();
 b15zdnd11an1n64x5 FILLER_308_854 ();
 b15zdnd11an1n64x5 FILLER_308_918 ();
 b15zdnd11an1n64x5 FILLER_308_982 ();
 b15zdnd11an1n64x5 FILLER_308_1046 ();
 b15zdnd11an1n64x5 FILLER_308_1110 ();
 b15zdnd11an1n64x5 FILLER_308_1174 ();
 b15zdnd11an1n64x5 FILLER_308_1238 ();
 b15zdnd11an1n64x5 FILLER_308_1302 ();
 b15zdnd11an1n64x5 FILLER_308_1366 ();
 b15zdnd11an1n64x5 FILLER_308_1430 ();
 b15zdnd11an1n32x5 FILLER_308_1494 ();
 b15zdnd11an1n16x5 FILLER_308_1526 ();
 b15zdnd11an1n04x5 FILLER_308_1542 ();
 b15zdnd00an1n02x5 FILLER_308_1546 ();
 b15zdnd00an1n01x5 FILLER_308_1548 ();
 b15zdnd11an1n64x5 FILLER_308_1565 ();
 b15zdnd11an1n64x5 FILLER_308_1629 ();
 b15zdnd11an1n64x5 FILLER_308_1693 ();
 b15zdnd11an1n64x5 FILLER_308_1757 ();
 b15zdnd11an1n64x5 FILLER_308_1821 ();
 b15zdnd11an1n64x5 FILLER_308_1885 ();
 b15zdnd11an1n64x5 FILLER_308_1949 ();
 b15zdnd11an1n64x5 FILLER_308_2013 ();
 b15zdnd11an1n64x5 FILLER_308_2077 ();
 b15zdnd11an1n08x5 FILLER_308_2141 ();
 b15zdnd11an1n04x5 FILLER_308_2149 ();
 b15zdnd00an1n01x5 FILLER_308_2153 ();
 b15zdnd11an1n64x5 FILLER_308_2162 ();
 b15zdnd11an1n32x5 FILLER_308_2226 ();
 b15zdnd11an1n16x5 FILLER_308_2258 ();
 b15zdnd00an1n02x5 FILLER_308_2274 ();
 b15zdnd11an1n64x5 FILLER_309_0 ();
 b15zdnd11an1n64x5 FILLER_309_64 ();
 b15zdnd11an1n64x5 FILLER_309_128 ();
 b15zdnd11an1n64x5 FILLER_309_192 ();
 b15zdnd11an1n64x5 FILLER_309_256 ();
 b15zdnd11an1n64x5 FILLER_309_320 ();
 b15zdnd11an1n64x5 FILLER_309_384 ();
 b15zdnd11an1n64x5 FILLER_309_448 ();
 b15zdnd11an1n64x5 FILLER_309_512 ();
 b15zdnd11an1n64x5 FILLER_309_576 ();
 b15zdnd11an1n64x5 FILLER_309_640 ();
 b15zdnd11an1n64x5 FILLER_309_704 ();
 b15zdnd11an1n64x5 FILLER_309_768 ();
 b15zdnd11an1n64x5 FILLER_309_832 ();
 b15zdnd11an1n64x5 FILLER_309_896 ();
 b15zdnd11an1n16x5 FILLER_309_960 ();
 b15zdnd11an1n04x5 FILLER_309_976 ();
 b15zdnd00an1n02x5 FILLER_309_980 ();
 b15zdnd11an1n32x5 FILLER_309_1024 ();
 b15zdnd11an1n16x5 FILLER_309_1056 ();
 b15zdnd11an1n08x5 FILLER_309_1072 ();
 b15zdnd11an1n04x5 FILLER_309_1080 ();
 b15zdnd00an1n01x5 FILLER_309_1084 ();
 b15zdnd11an1n64x5 FILLER_309_1127 ();
 b15zdnd11an1n64x5 FILLER_309_1191 ();
 b15zdnd11an1n64x5 FILLER_309_1255 ();
 b15zdnd11an1n64x5 FILLER_309_1319 ();
 b15zdnd11an1n64x5 FILLER_309_1383 ();
 b15zdnd11an1n64x5 FILLER_309_1447 ();
 b15zdnd11an1n64x5 FILLER_309_1511 ();
 b15zdnd11an1n64x5 FILLER_309_1575 ();
 b15zdnd11an1n64x5 FILLER_309_1639 ();
 b15zdnd11an1n64x5 FILLER_309_1703 ();
 b15zdnd11an1n64x5 FILLER_309_1767 ();
 b15zdnd11an1n64x5 FILLER_309_1831 ();
 b15zdnd11an1n64x5 FILLER_309_1895 ();
 b15zdnd11an1n64x5 FILLER_309_1959 ();
 b15zdnd11an1n64x5 FILLER_309_2023 ();
 b15zdnd11an1n64x5 FILLER_309_2087 ();
 b15zdnd11an1n64x5 FILLER_309_2151 ();
 b15zdnd11an1n64x5 FILLER_309_2215 ();
 b15zdnd11an1n04x5 FILLER_309_2279 ();
 b15zdnd00an1n01x5 FILLER_309_2283 ();
 b15zdnd11an1n64x5 FILLER_310_8 ();
 b15zdnd11an1n64x5 FILLER_310_72 ();
 b15zdnd11an1n64x5 FILLER_310_136 ();
 b15zdnd11an1n64x5 FILLER_310_200 ();
 b15zdnd11an1n64x5 FILLER_310_264 ();
 b15zdnd11an1n64x5 FILLER_310_328 ();
 b15zdnd11an1n64x5 FILLER_310_392 ();
 b15zdnd11an1n64x5 FILLER_310_456 ();
 b15zdnd11an1n64x5 FILLER_310_520 ();
 b15zdnd11an1n64x5 FILLER_310_584 ();
 b15zdnd11an1n64x5 FILLER_310_648 ();
 b15zdnd11an1n04x5 FILLER_310_712 ();
 b15zdnd00an1n02x5 FILLER_310_716 ();
 b15zdnd11an1n64x5 FILLER_310_726 ();
 b15zdnd11an1n64x5 FILLER_310_790 ();
 b15zdnd11an1n64x5 FILLER_310_854 ();
 b15zdnd11an1n64x5 FILLER_310_918 ();
 b15zdnd11an1n64x5 FILLER_310_982 ();
 b15zdnd11an1n64x5 FILLER_310_1046 ();
 b15zdnd11an1n64x5 FILLER_310_1110 ();
 b15zdnd11an1n64x5 FILLER_310_1174 ();
 b15zdnd11an1n32x5 FILLER_310_1238 ();
 b15zdnd11an1n04x5 FILLER_310_1270 ();
 b15zdnd00an1n02x5 FILLER_310_1274 ();
 b15zdnd00an1n01x5 FILLER_310_1276 ();
 b15zdnd11an1n16x5 FILLER_310_1319 ();
 b15zdnd11an1n08x5 FILLER_310_1335 ();
 b15zdnd11an1n04x5 FILLER_310_1343 ();
 b15zdnd00an1n01x5 FILLER_310_1347 ();
 b15zdnd11an1n64x5 FILLER_310_1390 ();
 b15zdnd11an1n64x5 FILLER_310_1454 ();
 b15zdnd11an1n64x5 FILLER_310_1518 ();
 b15zdnd11an1n64x5 FILLER_310_1582 ();
 b15zdnd11an1n64x5 FILLER_310_1646 ();
 b15zdnd11an1n64x5 FILLER_310_1710 ();
 b15zdnd11an1n64x5 FILLER_310_1774 ();
 b15zdnd11an1n64x5 FILLER_310_1838 ();
 b15zdnd11an1n64x5 FILLER_310_1902 ();
 b15zdnd11an1n64x5 FILLER_310_1966 ();
 b15zdnd11an1n64x5 FILLER_310_2030 ();
 b15zdnd11an1n32x5 FILLER_310_2094 ();
 b15zdnd11an1n16x5 FILLER_310_2126 ();
 b15zdnd11an1n08x5 FILLER_310_2142 ();
 b15zdnd11an1n04x5 FILLER_310_2150 ();
 b15zdnd11an1n64x5 FILLER_310_2162 ();
 b15zdnd11an1n32x5 FILLER_310_2226 ();
 b15zdnd11an1n16x5 FILLER_310_2258 ();
 b15zdnd00an1n02x5 FILLER_310_2274 ();
 b15zdnd11an1n64x5 FILLER_311_0 ();
 b15zdnd11an1n64x5 FILLER_311_64 ();
 b15zdnd11an1n64x5 FILLER_311_128 ();
 b15zdnd11an1n64x5 FILLER_311_192 ();
 b15zdnd11an1n64x5 FILLER_311_256 ();
 b15zdnd11an1n64x5 FILLER_311_320 ();
 b15zdnd11an1n64x5 FILLER_311_384 ();
 b15zdnd11an1n64x5 FILLER_311_448 ();
 b15zdnd11an1n64x5 FILLER_311_512 ();
 b15zdnd11an1n64x5 FILLER_311_576 ();
 b15zdnd11an1n64x5 FILLER_311_640 ();
 b15zdnd11an1n64x5 FILLER_311_704 ();
 b15zdnd11an1n64x5 FILLER_311_768 ();
 b15zdnd11an1n64x5 FILLER_311_832 ();
 b15zdnd11an1n64x5 FILLER_311_896 ();
 b15zdnd11an1n64x5 FILLER_311_960 ();
 b15zdnd11an1n64x5 FILLER_311_1024 ();
 b15zdnd11an1n08x5 FILLER_311_1088 ();
 b15zdnd11an1n04x5 FILLER_311_1096 ();
 b15zdnd00an1n01x5 FILLER_311_1100 ();
 b15zdnd11an1n64x5 FILLER_311_1143 ();
 b15zdnd11an1n64x5 FILLER_311_1207 ();
 b15zdnd11an1n64x5 FILLER_311_1271 ();
 b15zdnd11an1n64x5 FILLER_311_1335 ();
 b15zdnd11an1n64x5 FILLER_311_1399 ();
 b15zdnd11an1n64x5 FILLER_311_1463 ();
 b15zdnd11an1n64x5 FILLER_311_1527 ();
 b15zdnd11an1n64x5 FILLER_311_1591 ();
 b15zdnd11an1n64x5 FILLER_311_1655 ();
 b15zdnd11an1n64x5 FILLER_311_1719 ();
 b15zdnd11an1n64x5 FILLER_311_1783 ();
 b15zdnd11an1n64x5 FILLER_311_1847 ();
 b15zdnd11an1n64x5 FILLER_311_1911 ();
 b15zdnd11an1n64x5 FILLER_311_1975 ();
 b15zdnd11an1n64x5 FILLER_311_2039 ();
 b15zdnd11an1n64x5 FILLER_311_2103 ();
 b15zdnd11an1n64x5 FILLER_311_2167 ();
 b15zdnd11an1n32x5 FILLER_311_2231 ();
 b15zdnd11an1n16x5 FILLER_311_2263 ();
 b15zdnd11an1n04x5 FILLER_311_2279 ();
 b15zdnd00an1n01x5 FILLER_311_2283 ();
 b15zdnd11an1n64x5 FILLER_312_8 ();
 b15zdnd11an1n64x5 FILLER_312_72 ();
 b15zdnd11an1n64x5 FILLER_312_136 ();
 b15zdnd11an1n64x5 FILLER_312_200 ();
 b15zdnd11an1n64x5 FILLER_312_264 ();
 b15zdnd11an1n64x5 FILLER_312_328 ();
 b15zdnd11an1n64x5 FILLER_312_392 ();
 b15zdnd11an1n64x5 FILLER_312_456 ();
 b15zdnd11an1n64x5 FILLER_312_520 ();
 b15zdnd11an1n64x5 FILLER_312_584 ();
 b15zdnd11an1n64x5 FILLER_312_648 ();
 b15zdnd11an1n04x5 FILLER_312_712 ();
 b15zdnd00an1n02x5 FILLER_312_716 ();
 b15zdnd11an1n64x5 FILLER_312_726 ();
 b15zdnd11an1n64x5 FILLER_312_790 ();
 b15zdnd11an1n64x5 FILLER_312_854 ();
 b15zdnd11an1n64x5 FILLER_312_918 ();
 b15zdnd11an1n64x5 FILLER_312_982 ();
 b15zdnd11an1n32x5 FILLER_312_1046 ();
 b15zdnd11an1n16x5 FILLER_312_1078 ();
 b15zdnd00an1n02x5 FILLER_312_1094 ();
 b15zdnd00an1n01x5 FILLER_312_1096 ();
 b15zdnd11an1n64x5 FILLER_312_1139 ();
 b15zdnd11an1n64x5 FILLER_312_1203 ();
 b15zdnd11an1n64x5 FILLER_312_1267 ();
 b15zdnd11an1n64x5 FILLER_312_1331 ();
 b15zdnd11an1n64x5 FILLER_312_1395 ();
 b15zdnd11an1n64x5 FILLER_312_1459 ();
 b15zdnd11an1n64x5 FILLER_312_1523 ();
 b15zdnd11an1n64x5 FILLER_312_1587 ();
 b15zdnd11an1n64x5 FILLER_312_1651 ();
 b15zdnd11an1n64x5 FILLER_312_1715 ();
 b15zdnd11an1n64x5 FILLER_312_1779 ();
 b15zdnd11an1n64x5 FILLER_312_1843 ();
 b15zdnd11an1n64x5 FILLER_312_1907 ();
 b15zdnd11an1n64x5 FILLER_312_1971 ();
 b15zdnd11an1n64x5 FILLER_312_2035 ();
 b15zdnd11an1n32x5 FILLER_312_2099 ();
 b15zdnd11an1n16x5 FILLER_312_2131 ();
 b15zdnd11an1n04x5 FILLER_312_2147 ();
 b15zdnd00an1n02x5 FILLER_312_2151 ();
 b15zdnd00an1n01x5 FILLER_312_2153 ();
 b15zdnd11an1n64x5 FILLER_312_2162 ();
 b15zdnd11an1n32x5 FILLER_312_2226 ();
 b15zdnd11an1n16x5 FILLER_312_2258 ();
 b15zdnd00an1n02x5 FILLER_312_2274 ();
 b15zdnd11an1n64x5 FILLER_313_0 ();
 b15zdnd11an1n64x5 FILLER_313_64 ();
 b15zdnd11an1n64x5 FILLER_313_128 ();
 b15zdnd11an1n64x5 FILLER_313_192 ();
 b15zdnd11an1n64x5 FILLER_313_256 ();
 b15zdnd11an1n64x5 FILLER_313_320 ();
 b15zdnd11an1n64x5 FILLER_313_384 ();
 b15zdnd11an1n64x5 FILLER_313_448 ();
 b15zdnd11an1n64x5 FILLER_313_512 ();
 b15zdnd11an1n64x5 FILLER_313_576 ();
 b15zdnd11an1n64x5 FILLER_313_640 ();
 b15zdnd11an1n64x5 FILLER_313_704 ();
 b15zdnd11an1n64x5 FILLER_313_768 ();
 b15zdnd11an1n64x5 FILLER_313_832 ();
 b15zdnd11an1n64x5 FILLER_313_896 ();
 b15zdnd11an1n64x5 FILLER_313_960 ();
 b15zdnd11an1n64x5 FILLER_313_1024 ();
 b15zdnd11an1n64x5 FILLER_313_1088 ();
 b15zdnd11an1n64x5 FILLER_313_1152 ();
 b15zdnd11an1n64x5 FILLER_313_1216 ();
 b15zdnd11an1n64x5 FILLER_313_1280 ();
 b15zdnd11an1n64x5 FILLER_313_1344 ();
 b15zdnd11an1n64x5 FILLER_313_1408 ();
 b15zdnd11an1n64x5 FILLER_313_1472 ();
 b15zdnd11an1n64x5 FILLER_313_1536 ();
 b15zdnd11an1n64x5 FILLER_313_1600 ();
 b15zdnd11an1n64x5 FILLER_313_1664 ();
 b15zdnd11an1n64x5 FILLER_313_1728 ();
 b15zdnd11an1n64x5 FILLER_313_1792 ();
 b15zdnd11an1n64x5 FILLER_313_1856 ();
 b15zdnd11an1n64x5 FILLER_313_1920 ();
 b15zdnd11an1n64x5 FILLER_313_1984 ();
 b15zdnd11an1n64x5 FILLER_313_2048 ();
 b15zdnd11an1n64x5 FILLER_313_2112 ();
 b15zdnd11an1n64x5 FILLER_313_2176 ();
 b15zdnd11an1n32x5 FILLER_313_2240 ();
 b15zdnd11an1n08x5 FILLER_313_2272 ();
 b15zdnd11an1n04x5 FILLER_313_2280 ();
 b15zdnd11an1n64x5 FILLER_314_8 ();
 b15zdnd11an1n64x5 FILLER_314_72 ();
 b15zdnd11an1n64x5 FILLER_314_136 ();
 b15zdnd11an1n64x5 FILLER_314_200 ();
 b15zdnd11an1n64x5 FILLER_314_264 ();
 b15zdnd11an1n64x5 FILLER_314_328 ();
 b15zdnd11an1n64x5 FILLER_314_392 ();
 b15zdnd11an1n64x5 FILLER_314_456 ();
 b15zdnd11an1n64x5 FILLER_314_520 ();
 b15zdnd11an1n64x5 FILLER_314_584 ();
 b15zdnd11an1n64x5 FILLER_314_648 ();
 b15zdnd11an1n04x5 FILLER_314_712 ();
 b15zdnd00an1n02x5 FILLER_314_716 ();
 b15zdnd11an1n64x5 FILLER_314_726 ();
 b15zdnd11an1n64x5 FILLER_314_790 ();
 b15zdnd11an1n64x5 FILLER_314_854 ();
 b15zdnd11an1n64x5 FILLER_314_918 ();
 b15zdnd11an1n64x5 FILLER_314_982 ();
 b15zdnd11an1n64x5 FILLER_314_1046 ();
 b15zdnd11an1n64x5 FILLER_314_1110 ();
 b15zdnd11an1n64x5 FILLER_314_1174 ();
 b15zdnd11an1n64x5 FILLER_314_1238 ();
 b15zdnd11an1n64x5 FILLER_314_1302 ();
 b15zdnd11an1n64x5 FILLER_314_1366 ();
 b15zdnd11an1n64x5 FILLER_314_1430 ();
 b15zdnd11an1n64x5 FILLER_314_1494 ();
 b15zdnd11an1n64x5 FILLER_314_1558 ();
 b15zdnd11an1n64x5 FILLER_314_1622 ();
 b15zdnd11an1n64x5 FILLER_314_1686 ();
 b15zdnd11an1n64x5 FILLER_314_1750 ();
 b15zdnd11an1n64x5 FILLER_314_1814 ();
 b15zdnd11an1n64x5 FILLER_314_1878 ();
 b15zdnd11an1n64x5 FILLER_314_1942 ();
 b15zdnd11an1n64x5 FILLER_314_2006 ();
 b15zdnd11an1n64x5 FILLER_314_2070 ();
 b15zdnd11an1n16x5 FILLER_314_2134 ();
 b15zdnd11an1n04x5 FILLER_314_2150 ();
 b15zdnd11an1n64x5 FILLER_314_2162 ();
 b15zdnd11an1n32x5 FILLER_314_2226 ();
 b15zdnd11an1n16x5 FILLER_314_2258 ();
 b15zdnd00an1n02x5 FILLER_314_2274 ();
 b15zdnd11an1n64x5 FILLER_315_0 ();
 b15zdnd11an1n64x5 FILLER_315_64 ();
 b15zdnd11an1n64x5 FILLER_315_128 ();
 b15zdnd11an1n64x5 FILLER_315_192 ();
 b15zdnd11an1n64x5 FILLER_315_256 ();
 b15zdnd11an1n64x5 FILLER_315_320 ();
 b15zdnd11an1n64x5 FILLER_315_384 ();
 b15zdnd11an1n64x5 FILLER_315_448 ();
 b15zdnd11an1n64x5 FILLER_315_512 ();
 b15zdnd11an1n64x5 FILLER_315_576 ();
 b15zdnd11an1n64x5 FILLER_315_640 ();
 b15zdnd11an1n64x5 FILLER_315_704 ();
 b15zdnd11an1n64x5 FILLER_315_768 ();
 b15zdnd11an1n64x5 FILLER_315_832 ();
 b15zdnd11an1n64x5 FILLER_315_896 ();
 b15zdnd11an1n64x5 FILLER_315_960 ();
 b15zdnd11an1n64x5 FILLER_315_1024 ();
 b15zdnd11an1n64x5 FILLER_315_1088 ();
 b15zdnd11an1n64x5 FILLER_315_1152 ();
 b15zdnd11an1n64x5 FILLER_315_1216 ();
 b15zdnd11an1n64x5 FILLER_315_1280 ();
 b15zdnd11an1n64x5 FILLER_315_1344 ();
 b15zdnd11an1n64x5 FILLER_315_1408 ();
 b15zdnd11an1n64x5 FILLER_315_1472 ();
 b15zdnd11an1n64x5 FILLER_315_1536 ();
 b15zdnd11an1n64x5 FILLER_315_1600 ();
 b15zdnd11an1n64x5 FILLER_315_1664 ();
 b15zdnd11an1n64x5 FILLER_315_1728 ();
 b15zdnd11an1n64x5 FILLER_315_1792 ();
 b15zdnd11an1n64x5 FILLER_315_1856 ();
 b15zdnd11an1n64x5 FILLER_315_1920 ();
 b15zdnd11an1n64x5 FILLER_315_1984 ();
 b15zdnd11an1n64x5 FILLER_315_2048 ();
 b15zdnd11an1n64x5 FILLER_315_2112 ();
 b15zdnd11an1n64x5 FILLER_315_2176 ();
 b15zdnd11an1n32x5 FILLER_315_2240 ();
 b15zdnd11an1n08x5 FILLER_315_2272 ();
 b15zdnd11an1n04x5 FILLER_315_2280 ();
 b15zdnd11an1n64x5 FILLER_316_8 ();
 b15zdnd11an1n64x5 FILLER_316_72 ();
 b15zdnd11an1n64x5 FILLER_316_136 ();
 b15zdnd11an1n64x5 FILLER_316_200 ();
 b15zdnd11an1n64x5 FILLER_316_264 ();
 b15zdnd11an1n64x5 FILLER_316_328 ();
 b15zdnd11an1n64x5 FILLER_316_392 ();
 b15zdnd11an1n64x5 FILLER_316_456 ();
 b15zdnd11an1n64x5 FILLER_316_520 ();
 b15zdnd11an1n64x5 FILLER_316_584 ();
 b15zdnd11an1n64x5 FILLER_316_648 ();
 b15zdnd11an1n04x5 FILLER_316_712 ();
 b15zdnd00an1n02x5 FILLER_316_716 ();
 b15zdnd11an1n64x5 FILLER_316_726 ();
 b15zdnd11an1n64x5 FILLER_316_790 ();
 b15zdnd11an1n64x5 FILLER_316_854 ();
 b15zdnd11an1n64x5 FILLER_316_918 ();
 b15zdnd11an1n64x5 FILLER_316_982 ();
 b15zdnd11an1n64x5 FILLER_316_1046 ();
 b15zdnd11an1n64x5 FILLER_316_1110 ();
 b15zdnd11an1n64x5 FILLER_316_1174 ();
 b15zdnd11an1n64x5 FILLER_316_1238 ();
 b15zdnd11an1n64x5 FILLER_316_1302 ();
 b15zdnd11an1n64x5 FILLER_316_1366 ();
 b15zdnd11an1n64x5 FILLER_316_1430 ();
 b15zdnd11an1n64x5 FILLER_316_1494 ();
 b15zdnd11an1n64x5 FILLER_316_1558 ();
 b15zdnd11an1n64x5 FILLER_316_1622 ();
 b15zdnd11an1n64x5 FILLER_316_1686 ();
 b15zdnd11an1n64x5 FILLER_316_1750 ();
 b15zdnd11an1n64x5 FILLER_316_1814 ();
 b15zdnd11an1n64x5 FILLER_316_1878 ();
 b15zdnd11an1n64x5 FILLER_316_1942 ();
 b15zdnd11an1n64x5 FILLER_316_2006 ();
 b15zdnd11an1n64x5 FILLER_316_2070 ();
 b15zdnd11an1n16x5 FILLER_316_2134 ();
 b15zdnd11an1n04x5 FILLER_316_2150 ();
 b15zdnd11an1n64x5 FILLER_316_2162 ();
 b15zdnd11an1n32x5 FILLER_316_2226 ();
 b15zdnd11an1n16x5 FILLER_316_2258 ();
 b15zdnd00an1n02x5 FILLER_316_2274 ();
 b15zdnd11an1n64x5 FILLER_317_0 ();
 b15zdnd11an1n64x5 FILLER_317_64 ();
 b15zdnd11an1n64x5 FILLER_317_128 ();
 b15zdnd11an1n64x5 FILLER_317_192 ();
 b15zdnd11an1n64x5 FILLER_317_256 ();
 b15zdnd11an1n64x5 FILLER_317_320 ();
 b15zdnd11an1n64x5 FILLER_317_384 ();
 b15zdnd11an1n64x5 FILLER_317_448 ();
 b15zdnd11an1n64x5 FILLER_317_512 ();
 b15zdnd11an1n64x5 FILLER_317_576 ();
 b15zdnd11an1n64x5 FILLER_317_640 ();
 b15zdnd11an1n64x5 FILLER_317_704 ();
 b15zdnd11an1n64x5 FILLER_317_768 ();
 b15zdnd11an1n64x5 FILLER_317_832 ();
 b15zdnd11an1n64x5 FILLER_317_896 ();
 b15zdnd11an1n64x5 FILLER_317_960 ();
 b15zdnd11an1n64x5 FILLER_317_1024 ();
 b15zdnd11an1n64x5 FILLER_317_1088 ();
 b15zdnd11an1n64x5 FILLER_317_1152 ();
 b15zdnd11an1n64x5 FILLER_317_1216 ();
 b15zdnd11an1n64x5 FILLER_317_1280 ();
 b15zdnd11an1n64x5 FILLER_317_1344 ();
 b15zdnd11an1n64x5 FILLER_317_1408 ();
 b15zdnd11an1n64x5 FILLER_317_1472 ();
 b15zdnd11an1n64x5 FILLER_317_1536 ();
 b15zdnd11an1n64x5 FILLER_317_1600 ();
 b15zdnd11an1n64x5 FILLER_317_1664 ();
 b15zdnd11an1n64x5 FILLER_317_1728 ();
 b15zdnd11an1n64x5 FILLER_317_1792 ();
 b15zdnd11an1n64x5 FILLER_317_1856 ();
 b15zdnd11an1n64x5 FILLER_317_1920 ();
 b15zdnd11an1n64x5 FILLER_317_1984 ();
 b15zdnd11an1n64x5 FILLER_317_2048 ();
 b15zdnd11an1n64x5 FILLER_317_2112 ();
 b15zdnd11an1n64x5 FILLER_317_2176 ();
 b15zdnd11an1n32x5 FILLER_317_2240 ();
 b15zdnd11an1n08x5 FILLER_317_2272 ();
 b15zdnd11an1n04x5 FILLER_317_2280 ();
 b15zdnd11an1n64x5 FILLER_318_8 ();
 b15zdnd11an1n64x5 FILLER_318_72 ();
 b15zdnd11an1n64x5 FILLER_318_136 ();
 b15zdnd11an1n64x5 FILLER_318_200 ();
 b15zdnd11an1n64x5 FILLER_318_264 ();
 b15zdnd11an1n64x5 FILLER_318_328 ();
 b15zdnd11an1n64x5 FILLER_318_392 ();
 b15zdnd11an1n64x5 FILLER_318_456 ();
 b15zdnd11an1n64x5 FILLER_318_520 ();
 b15zdnd11an1n64x5 FILLER_318_584 ();
 b15zdnd11an1n64x5 FILLER_318_648 ();
 b15zdnd11an1n04x5 FILLER_318_712 ();
 b15zdnd00an1n02x5 FILLER_318_716 ();
 b15zdnd11an1n64x5 FILLER_318_726 ();
 b15zdnd11an1n64x5 FILLER_318_790 ();
 b15zdnd11an1n64x5 FILLER_318_854 ();
 b15zdnd11an1n64x5 FILLER_318_918 ();
 b15zdnd11an1n64x5 FILLER_318_982 ();
 b15zdnd11an1n64x5 FILLER_318_1046 ();
 b15zdnd11an1n64x5 FILLER_318_1110 ();
 b15zdnd11an1n64x5 FILLER_318_1174 ();
 b15zdnd11an1n64x5 FILLER_318_1238 ();
 b15zdnd11an1n64x5 FILLER_318_1302 ();
 b15zdnd11an1n64x5 FILLER_318_1366 ();
 b15zdnd11an1n64x5 FILLER_318_1430 ();
 b15zdnd11an1n64x5 FILLER_318_1494 ();
 b15zdnd11an1n64x5 FILLER_318_1558 ();
 b15zdnd11an1n64x5 FILLER_318_1622 ();
 b15zdnd11an1n64x5 FILLER_318_1686 ();
 b15zdnd11an1n64x5 FILLER_318_1750 ();
 b15zdnd11an1n64x5 FILLER_318_1814 ();
 b15zdnd11an1n32x5 FILLER_318_1878 ();
 b15zdnd11an1n08x5 FILLER_318_1910 ();
 b15zdnd00an1n02x5 FILLER_318_1918 ();
 b15zdnd00an1n01x5 FILLER_318_1920 ();
 b15zdnd11an1n64x5 FILLER_318_1929 ();
 b15zdnd11an1n64x5 FILLER_318_1993 ();
 b15zdnd11an1n64x5 FILLER_318_2057 ();
 b15zdnd11an1n32x5 FILLER_318_2121 ();
 b15zdnd00an1n01x5 FILLER_318_2153 ();
 b15zdnd11an1n64x5 FILLER_318_2162 ();
 b15zdnd11an1n32x5 FILLER_318_2226 ();
 b15zdnd11an1n16x5 FILLER_318_2258 ();
 b15zdnd00an1n02x5 FILLER_318_2274 ();
 b15zdnd11an1n64x5 FILLER_319_0 ();
 b15zdnd11an1n64x5 FILLER_319_64 ();
 b15zdnd11an1n64x5 FILLER_319_128 ();
 b15zdnd11an1n64x5 FILLER_319_192 ();
 b15zdnd11an1n64x5 FILLER_319_256 ();
 b15zdnd11an1n64x5 FILLER_319_320 ();
 b15zdnd11an1n64x5 FILLER_319_384 ();
 b15zdnd11an1n64x5 FILLER_319_448 ();
 b15zdnd11an1n64x5 FILLER_319_512 ();
 b15zdnd11an1n64x5 FILLER_319_576 ();
 b15zdnd11an1n64x5 FILLER_319_640 ();
 b15zdnd11an1n64x5 FILLER_319_704 ();
 b15zdnd11an1n64x5 FILLER_319_768 ();
 b15zdnd11an1n64x5 FILLER_319_832 ();
 b15zdnd11an1n64x5 FILLER_319_896 ();
 b15zdnd11an1n64x5 FILLER_319_960 ();
 b15zdnd11an1n64x5 FILLER_319_1024 ();
 b15zdnd11an1n64x5 FILLER_319_1088 ();
 b15zdnd11an1n64x5 FILLER_319_1152 ();
 b15zdnd11an1n64x5 FILLER_319_1216 ();
 b15zdnd11an1n64x5 FILLER_319_1280 ();
 b15zdnd11an1n64x5 FILLER_319_1344 ();
 b15zdnd11an1n64x5 FILLER_319_1408 ();
 b15zdnd11an1n64x5 FILLER_319_1472 ();
 b15zdnd11an1n64x5 FILLER_319_1536 ();
 b15zdnd11an1n64x5 FILLER_319_1600 ();
 b15zdnd11an1n64x5 FILLER_319_1664 ();
 b15zdnd11an1n64x5 FILLER_319_1728 ();
 b15zdnd11an1n64x5 FILLER_319_1792 ();
 b15zdnd11an1n64x5 FILLER_319_1856 ();
 b15zdnd11an1n64x5 FILLER_319_1920 ();
 b15zdnd11an1n64x5 FILLER_319_1984 ();
 b15zdnd11an1n64x5 FILLER_319_2048 ();
 b15zdnd11an1n64x5 FILLER_319_2112 ();
 b15zdnd11an1n64x5 FILLER_319_2176 ();
 b15zdnd11an1n32x5 FILLER_319_2240 ();
 b15zdnd11an1n08x5 FILLER_319_2272 ();
 b15zdnd11an1n04x5 FILLER_319_2280 ();
 b15zdnd11an1n64x5 FILLER_320_8 ();
 b15zdnd11an1n64x5 FILLER_320_72 ();
 b15zdnd11an1n64x5 FILLER_320_136 ();
 b15zdnd11an1n64x5 FILLER_320_200 ();
 b15zdnd11an1n64x5 FILLER_320_264 ();
 b15zdnd11an1n64x5 FILLER_320_328 ();
 b15zdnd11an1n64x5 FILLER_320_392 ();
 b15zdnd11an1n64x5 FILLER_320_456 ();
 b15zdnd11an1n64x5 FILLER_320_520 ();
 b15zdnd11an1n64x5 FILLER_320_584 ();
 b15zdnd11an1n64x5 FILLER_320_648 ();
 b15zdnd11an1n04x5 FILLER_320_712 ();
 b15zdnd00an1n02x5 FILLER_320_716 ();
 b15zdnd11an1n64x5 FILLER_320_726 ();
 b15zdnd11an1n64x5 FILLER_320_790 ();
 b15zdnd11an1n64x5 FILLER_320_854 ();
 b15zdnd11an1n64x5 FILLER_320_918 ();
 b15zdnd11an1n64x5 FILLER_320_982 ();
 b15zdnd11an1n64x5 FILLER_320_1046 ();
 b15zdnd11an1n64x5 FILLER_320_1110 ();
 b15zdnd11an1n64x5 FILLER_320_1174 ();
 b15zdnd11an1n64x5 FILLER_320_1238 ();
 b15zdnd11an1n64x5 FILLER_320_1302 ();
 b15zdnd11an1n64x5 FILLER_320_1366 ();
 b15zdnd11an1n64x5 FILLER_320_1430 ();
 b15zdnd11an1n64x5 FILLER_320_1494 ();
 b15zdnd11an1n64x5 FILLER_320_1558 ();
 b15zdnd11an1n64x5 FILLER_320_1622 ();
 b15zdnd11an1n64x5 FILLER_320_1686 ();
 b15zdnd11an1n64x5 FILLER_320_1750 ();
 b15zdnd11an1n64x5 FILLER_320_1814 ();
 b15zdnd11an1n64x5 FILLER_320_1878 ();
 b15zdnd11an1n64x5 FILLER_320_1942 ();
 b15zdnd11an1n64x5 FILLER_320_2006 ();
 b15zdnd11an1n64x5 FILLER_320_2070 ();
 b15zdnd11an1n16x5 FILLER_320_2134 ();
 b15zdnd11an1n04x5 FILLER_320_2150 ();
 b15zdnd11an1n64x5 FILLER_320_2162 ();
 b15zdnd11an1n32x5 FILLER_320_2226 ();
 b15zdnd11an1n16x5 FILLER_320_2258 ();
 b15zdnd00an1n02x5 FILLER_320_2274 ();
 b15zdnd11an1n64x5 FILLER_321_0 ();
 b15zdnd11an1n64x5 FILLER_321_64 ();
 b15zdnd11an1n64x5 FILLER_321_128 ();
 b15zdnd11an1n64x5 FILLER_321_192 ();
 b15zdnd11an1n64x5 FILLER_321_256 ();
 b15zdnd11an1n64x5 FILLER_321_320 ();
 b15zdnd11an1n64x5 FILLER_321_384 ();
 b15zdnd11an1n64x5 FILLER_321_448 ();
 b15zdnd11an1n64x5 FILLER_321_512 ();
 b15zdnd11an1n64x5 FILLER_321_576 ();
 b15zdnd11an1n64x5 FILLER_321_640 ();
 b15zdnd11an1n64x5 FILLER_321_704 ();
 b15zdnd11an1n64x5 FILLER_321_768 ();
 b15zdnd11an1n64x5 FILLER_321_832 ();
 b15zdnd11an1n64x5 FILLER_321_896 ();
 b15zdnd11an1n64x5 FILLER_321_960 ();
 b15zdnd11an1n64x5 FILLER_321_1024 ();
 b15zdnd11an1n64x5 FILLER_321_1088 ();
 b15zdnd11an1n64x5 FILLER_321_1152 ();
 b15zdnd11an1n64x5 FILLER_321_1216 ();
 b15zdnd11an1n64x5 FILLER_321_1280 ();
 b15zdnd11an1n64x5 FILLER_321_1344 ();
 b15zdnd11an1n64x5 FILLER_321_1408 ();
 b15zdnd11an1n64x5 FILLER_321_1472 ();
 b15zdnd11an1n64x5 FILLER_321_1536 ();
 b15zdnd11an1n64x5 FILLER_321_1600 ();
 b15zdnd11an1n64x5 FILLER_321_1664 ();
 b15zdnd11an1n64x5 FILLER_321_1728 ();
 b15zdnd11an1n64x5 FILLER_321_1792 ();
 b15zdnd11an1n64x5 FILLER_321_1856 ();
 b15zdnd11an1n64x5 FILLER_321_1920 ();
 b15zdnd11an1n64x5 FILLER_321_1984 ();
 b15zdnd11an1n64x5 FILLER_321_2048 ();
 b15zdnd11an1n64x5 FILLER_321_2112 ();
 b15zdnd11an1n64x5 FILLER_321_2176 ();
 b15zdnd11an1n32x5 FILLER_321_2240 ();
 b15zdnd11an1n08x5 FILLER_321_2272 ();
 b15zdnd11an1n04x5 FILLER_321_2280 ();
 b15zdnd11an1n64x5 FILLER_322_8 ();
 b15zdnd11an1n64x5 FILLER_322_72 ();
 b15zdnd11an1n64x5 FILLER_322_136 ();
 b15zdnd11an1n64x5 FILLER_322_200 ();
 b15zdnd11an1n64x5 FILLER_322_264 ();
 b15zdnd11an1n64x5 FILLER_322_328 ();
 b15zdnd11an1n64x5 FILLER_322_392 ();
 b15zdnd11an1n64x5 FILLER_322_456 ();
 b15zdnd11an1n64x5 FILLER_322_520 ();
 b15zdnd11an1n64x5 FILLER_322_584 ();
 b15zdnd11an1n64x5 FILLER_322_648 ();
 b15zdnd11an1n04x5 FILLER_322_712 ();
 b15zdnd00an1n02x5 FILLER_322_716 ();
 b15zdnd11an1n64x5 FILLER_322_726 ();
 b15zdnd11an1n64x5 FILLER_322_790 ();
 b15zdnd11an1n64x5 FILLER_322_854 ();
 b15zdnd11an1n64x5 FILLER_322_918 ();
 b15zdnd11an1n64x5 FILLER_322_982 ();
 b15zdnd11an1n64x5 FILLER_322_1046 ();
 b15zdnd11an1n64x5 FILLER_322_1110 ();
 b15zdnd11an1n64x5 FILLER_322_1174 ();
 b15zdnd11an1n64x5 FILLER_322_1238 ();
 b15zdnd11an1n64x5 FILLER_322_1302 ();
 b15zdnd11an1n64x5 FILLER_322_1366 ();
 b15zdnd11an1n64x5 FILLER_322_1430 ();
 b15zdnd11an1n64x5 FILLER_322_1494 ();
 b15zdnd11an1n64x5 FILLER_322_1558 ();
 b15zdnd11an1n64x5 FILLER_322_1622 ();
 b15zdnd11an1n64x5 FILLER_322_1686 ();
 b15zdnd11an1n64x5 FILLER_322_1750 ();
 b15zdnd11an1n64x5 FILLER_322_1814 ();
 b15zdnd11an1n64x5 FILLER_322_1878 ();
 b15zdnd11an1n64x5 FILLER_322_1942 ();
 b15zdnd11an1n64x5 FILLER_322_2006 ();
 b15zdnd11an1n64x5 FILLER_322_2070 ();
 b15zdnd11an1n16x5 FILLER_322_2134 ();
 b15zdnd11an1n04x5 FILLER_322_2150 ();
 b15zdnd11an1n64x5 FILLER_322_2162 ();
 b15zdnd11an1n32x5 FILLER_322_2226 ();
 b15zdnd11an1n16x5 FILLER_322_2258 ();
 b15zdnd00an1n02x5 FILLER_322_2274 ();
 b15zdnd11an1n64x5 FILLER_323_0 ();
 b15zdnd11an1n64x5 FILLER_323_64 ();
 b15zdnd11an1n64x5 FILLER_323_128 ();
 b15zdnd11an1n64x5 FILLER_323_192 ();
 b15zdnd11an1n64x5 FILLER_323_256 ();
 b15zdnd11an1n64x5 FILLER_323_320 ();
 b15zdnd11an1n64x5 FILLER_323_384 ();
 b15zdnd11an1n64x5 FILLER_323_448 ();
 b15zdnd11an1n64x5 FILLER_323_512 ();
 b15zdnd11an1n64x5 FILLER_323_576 ();
 b15zdnd11an1n64x5 FILLER_323_640 ();
 b15zdnd11an1n64x5 FILLER_323_704 ();
 b15zdnd11an1n64x5 FILLER_323_768 ();
 b15zdnd11an1n64x5 FILLER_323_832 ();
 b15zdnd11an1n64x5 FILLER_323_896 ();
 b15zdnd11an1n64x5 FILLER_323_960 ();
 b15zdnd11an1n64x5 FILLER_323_1024 ();
 b15zdnd11an1n64x5 FILLER_323_1088 ();
 b15zdnd11an1n64x5 FILLER_323_1152 ();
 b15zdnd11an1n64x5 FILLER_323_1216 ();
 b15zdnd11an1n64x5 FILLER_323_1280 ();
 b15zdnd11an1n64x5 FILLER_323_1344 ();
 b15zdnd11an1n64x5 FILLER_323_1408 ();
 b15zdnd11an1n64x5 FILLER_323_1472 ();
 b15zdnd11an1n64x5 FILLER_323_1536 ();
 b15zdnd11an1n64x5 FILLER_323_1600 ();
 b15zdnd11an1n64x5 FILLER_323_1664 ();
 b15zdnd11an1n64x5 FILLER_323_1728 ();
 b15zdnd11an1n64x5 FILLER_323_1792 ();
 b15zdnd11an1n64x5 FILLER_323_1856 ();
 b15zdnd11an1n64x5 FILLER_323_1920 ();
 b15zdnd11an1n64x5 FILLER_323_1984 ();
 b15zdnd11an1n64x5 FILLER_323_2048 ();
 b15zdnd11an1n64x5 FILLER_323_2112 ();
 b15zdnd11an1n64x5 FILLER_323_2176 ();
 b15zdnd11an1n32x5 FILLER_323_2240 ();
 b15zdnd11an1n08x5 FILLER_323_2272 ();
 b15zdnd11an1n04x5 FILLER_323_2280 ();
 b15zdnd11an1n64x5 FILLER_324_8 ();
 b15zdnd11an1n64x5 FILLER_324_72 ();
 b15zdnd11an1n64x5 FILLER_324_136 ();
 b15zdnd11an1n64x5 FILLER_324_200 ();
 b15zdnd11an1n64x5 FILLER_324_264 ();
 b15zdnd11an1n64x5 FILLER_324_328 ();
 b15zdnd11an1n64x5 FILLER_324_392 ();
 b15zdnd11an1n64x5 FILLER_324_456 ();
 b15zdnd11an1n64x5 FILLER_324_520 ();
 b15zdnd11an1n64x5 FILLER_324_584 ();
 b15zdnd11an1n64x5 FILLER_324_648 ();
 b15zdnd11an1n04x5 FILLER_324_712 ();
 b15zdnd00an1n02x5 FILLER_324_716 ();
 b15zdnd11an1n64x5 FILLER_324_726 ();
 b15zdnd11an1n64x5 FILLER_324_790 ();
 b15zdnd11an1n64x5 FILLER_324_854 ();
 b15zdnd11an1n64x5 FILLER_324_918 ();
 b15zdnd11an1n64x5 FILLER_324_982 ();
 b15zdnd11an1n64x5 FILLER_324_1046 ();
 b15zdnd11an1n64x5 FILLER_324_1110 ();
 b15zdnd11an1n64x5 FILLER_324_1174 ();
 b15zdnd11an1n64x5 FILLER_324_1238 ();
 b15zdnd11an1n64x5 FILLER_324_1302 ();
 b15zdnd11an1n64x5 FILLER_324_1366 ();
 b15zdnd11an1n64x5 FILLER_324_1430 ();
 b15zdnd11an1n64x5 FILLER_324_1494 ();
 b15zdnd11an1n64x5 FILLER_324_1558 ();
 b15zdnd11an1n64x5 FILLER_324_1622 ();
 b15zdnd11an1n64x5 FILLER_324_1686 ();
 b15zdnd11an1n64x5 FILLER_324_1750 ();
 b15zdnd11an1n64x5 FILLER_324_1814 ();
 b15zdnd11an1n64x5 FILLER_324_1878 ();
 b15zdnd11an1n64x5 FILLER_324_1942 ();
 b15zdnd11an1n64x5 FILLER_324_2006 ();
 b15zdnd11an1n64x5 FILLER_324_2070 ();
 b15zdnd11an1n16x5 FILLER_324_2134 ();
 b15zdnd11an1n04x5 FILLER_324_2150 ();
 b15zdnd11an1n64x5 FILLER_324_2162 ();
 b15zdnd11an1n32x5 FILLER_324_2226 ();
 b15zdnd11an1n16x5 FILLER_324_2258 ();
 b15zdnd00an1n02x5 FILLER_324_2274 ();
 b15zdnd11an1n64x5 FILLER_325_0 ();
 b15zdnd11an1n64x5 FILLER_325_64 ();
 b15zdnd11an1n64x5 FILLER_325_128 ();
 b15zdnd11an1n64x5 FILLER_325_192 ();
 b15zdnd11an1n64x5 FILLER_325_256 ();
 b15zdnd11an1n64x5 FILLER_325_320 ();
 b15zdnd11an1n64x5 FILLER_325_384 ();
 b15zdnd11an1n64x5 FILLER_325_448 ();
 b15zdnd11an1n64x5 FILLER_325_512 ();
 b15zdnd11an1n64x5 FILLER_325_576 ();
 b15zdnd11an1n64x5 FILLER_325_640 ();
 b15zdnd11an1n64x5 FILLER_325_704 ();
 b15zdnd11an1n64x5 FILLER_325_768 ();
 b15zdnd11an1n64x5 FILLER_325_832 ();
 b15zdnd11an1n64x5 FILLER_325_896 ();
 b15zdnd11an1n64x5 FILLER_325_960 ();
 b15zdnd11an1n64x5 FILLER_325_1024 ();
 b15zdnd11an1n64x5 FILLER_325_1088 ();
 b15zdnd11an1n64x5 FILLER_325_1152 ();
 b15zdnd11an1n64x5 FILLER_325_1216 ();
 b15zdnd11an1n64x5 FILLER_325_1280 ();
 b15zdnd11an1n64x5 FILLER_325_1344 ();
 b15zdnd11an1n64x5 FILLER_325_1408 ();
 b15zdnd11an1n64x5 FILLER_325_1472 ();
 b15zdnd11an1n64x5 FILLER_325_1536 ();
 b15zdnd11an1n64x5 FILLER_325_1600 ();
 b15zdnd11an1n64x5 FILLER_325_1664 ();
 b15zdnd11an1n64x5 FILLER_325_1728 ();
 b15zdnd11an1n64x5 FILLER_325_1792 ();
 b15zdnd11an1n64x5 FILLER_325_1856 ();
 b15zdnd11an1n64x5 FILLER_325_1920 ();
 b15zdnd11an1n64x5 FILLER_325_1984 ();
 b15zdnd11an1n64x5 FILLER_325_2048 ();
 b15zdnd11an1n64x5 FILLER_325_2112 ();
 b15zdnd11an1n64x5 FILLER_325_2176 ();
 b15zdnd11an1n32x5 FILLER_325_2240 ();
 b15zdnd11an1n08x5 FILLER_325_2272 ();
 b15zdnd11an1n04x5 FILLER_325_2280 ();
 b15zdnd11an1n64x5 FILLER_326_8 ();
 b15zdnd11an1n64x5 FILLER_326_72 ();
 b15zdnd11an1n64x5 FILLER_326_136 ();
 b15zdnd11an1n64x5 FILLER_326_200 ();
 b15zdnd11an1n64x5 FILLER_326_264 ();
 b15zdnd11an1n64x5 FILLER_326_328 ();
 b15zdnd11an1n64x5 FILLER_326_392 ();
 b15zdnd11an1n64x5 FILLER_326_456 ();
 b15zdnd11an1n64x5 FILLER_326_520 ();
 b15zdnd11an1n64x5 FILLER_326_584 ();
 b15zdnd11an1n64x5 FILLER_326_648 ();
 b15zdnd11an1n04x5 FILLER_326_712 ();
 b15zdnd00an1n02x5 FILLER_326_716 ();
 b15zdnd11an1n64x5 FILLER_326_726 ();
 b15zdnd11an1n64x5 FILLER_326_790 ();
 b15zdnd11an1n64x5 FILLER_326_854 ();
 b15zdnd11an1n64x5 FILLER_326_918 ();
 b15zdnd11an1n64x5 FILLER_326_982 ();
 b15zdnd11an1n64x5 FILLER_326_1046 ();
 b15zdnd11an1n64x5 FILLER_326_1110 ();
 b15zdnd11an1n64x5 FILLER_326_1174 ();
 b15zdnd11an1n64x5 FILLER_326_1238 ();
 b15zdnd11an1n64x5 FILLER_326_1302 ();
 b15zdnd11an1n64x5 FILLER_326_1366 ();
 b15zdnd11an1n64x5 FILLER_326_1430 ();
 b15zdnd11an1n64x5 FILLER_326_1494 ();
 b15zdnd11an1n64x5 FILLER_326_1558 ();
 b15zdnd11an1n64x5 FILLER_326_1622 ();
 b15zdnd11an1n64x5 FILLER_326_1686 ();
 b15zdnd11an1n64x5 FILLER_326_1750 ();
 b15zdnd11an1n64x5 FILLER_326_1814 ();
 b15zdnd11an1n64x5 FILLER_326_1878 ();
 b15zdnd11an1n64x5 FILLER_326_1942 ();
 b15zdnd11an1n64x5 FILLER_326_2006 ();
 b15zdnd11an1n64x5 FILLER_326_2070 ();
 b15zdnd11an1n16x5 FILLER_326_2134 ();
 b15zdnd11an1n04x5 FILLER_326_2150 ();
 b15zdnd11an1n64x5 FILLER_326_2162 ();
 b15zdnd11an1n32x5 FILLER_326_2226 ();
 b15zdnd11an1n16x5 FILLER_326_2258 ();
 b15zdnd00an1n02x5 FILLER_326_2274 ();
 b15zdnd11an1n64x5 FILLER_327_0 ();
 b15zdnd11an1n64x5 FILLER_327_64 ();
 b15zdnd11an1n64x5 FILLER_327_128 ();
 b15zdnd11an1n64x5 FILLER_327_192 ();
 b15zdnd11an1n64x5 FILLER_327_256 ();
 b15zdnd11an1n64x5 FILLER_327_320 ();
 b15zdnd11an1n64x5 FILLER_327_384 ();
 b15zdnd11an1n64x5 FILLER_327_448 ();
 b15zdnd11an1n64x5 FILLER_327_512 ();
 b15zdnd11an1n64x5 FILLER_327_576 ();
 b15zdnd11an1n64x5 FILLER_327_640 ();
 b15zdnd11an1n64x5 FILLER_327_704 ();
 b15zdnd11an1n64x5 FILLER_327_768 ();
 b15zdnd11an1n64x5 FILLER_327_832 ();
 b15zdnd11an1n64x5 FILLER_327_896 ();
 b15zdnd11an1n64x5 FILLER_327_960 ();
 b15zdnd11an1n64x5 FILLER_327_1024 ();
 b15zdnd11an1n64x5 FILLER_327_1088 ();
 b15zdnd11an1n64x5 FILLER_327_1152 ();
 b15zdnd11an1n64x5 FILLER_327_1216 ();
 b15zdnd11an1n64x5 FILLER_327_1280 ();
 b15zdnd11an1n64x5 FILLER_327_1344 ();
 b15zdnd11an1n64x5 FILLER_327_1408 ();
 b15zdnd11an1n64x5 FILLER_327_1472 ();
 b15zdnd11an1n64x5 FILLER_327_1536 ();
 b15zdnd11an1n64x5 FILLER_327_1600 ();
 b15zdnd11an1n64x5 FILLER_327_1664 ();
 b15zdnd11an1n64x5 FILLER_327_1728 ();
 b15zdnd11an1n64x5 FILLER_327_1792 ();
 b15zdnd11an1n64x5 FILLER_327_1856 ();
 b15zdnd11an1n64x5 FILLER_327_1920 ();
 b15zdnd11an1n64x5 FILLER_327_1984 ();
 b15zdnd11an1n64x5 FILLER_327_2048 ();
 b15zdnd11an1n64x5 FILLER_327_2112 ();
 b15zdnd11an1n64x5 FILLER_327_2176 ();
 b15zdnd11an1n32x5 FILLER_327_2240 ();
 b15zdnd11an1n08x5 FILLER_327_2272 ();
 b15zdnd11an1n04x5 FILLER_327_2280 ();
 b15zdnd11an1n64x5 FILLER_328_8 ();
 b15zdnd11an1n64x5 FILLER_328_72 ();
 b15zdnd11an1n64x5 FILLER_328_136 ();
 b15zdnd11an1n64x5 FILLER_328_200 ();
 b15zdnd11an1n64x5 FILLER_328_264 ();
 b15zdnd11an1n64x5 FILLER_328_328 ();
 b15zdnd11an1n64x5 FILLER_328_392 ();
 b15zdnd11an1n64x5 FILLER_328_456 ();
 b15zdnd11an1n64x5 FILLER_328_520 ();
 b15zdnd11an1n64x5 FILLER_328_584 ();
 b15zdnd11an1n64x5 FILLER_328_648 ();
 b15zdnd11an1n04x5 FILLER_328_712 ();
 b15zdnd00an1n02x5 FILLER_328_716 ();
 b15zdnd11an1n64x5 FILLER_328_726 ();
 b15zdnd11an1n64x5 FILLER_328_790 ();
 b15zdnd11an1n64x5 FILLER_328_854 ();
 b15zdnd11an1n64x5 FILLER_328_918 ();
 b15zdnd11an1n64x5 FILLER_328_982 ();
 b15zdnd11an1n64x5 FILLER_328_1046 ();
 b15zdnd11an1n64x5 FILLER_328_1110 ();
 b15zdnd11an1n64x5 FILLER_328_1174 ();
 b15zdnd11an1n64x5 FILLER_328_1238 ();
 b15zdnd11an1n64x5 FILLER_328_1302 ();
 b15zdnd11an1n64x5 FILLER_328_1366 ();
 b15zdnd11an1n64x5 FILLER_328_1430 ();
 b15zdnd11an1n64x5 FILLER_328_1494 ();
 b15zdnd11an1n64x5 FILLER_328_1558 ();
 b15zdnd11an1n64x5 FILLER_328_1622 ();
 b15zdnd11an1n64x5 FILLER_328_1686 ();
 b15zdnd11an1n64x5 FILLER_328_1750 ();
 b15zdnd11an1n64x5 FILLER_328_1814 ();
 b15zdnd11an1n64x5 FILLER_328_1878 ();
 b15zdnd11an1n64x5 FILLER_328_1942 ();
 b15zdnd11an1n64x5 FILLER_328_2006 ();
 b15zdnd11an1n64x5 FILLER_328_2070 ();
 b15zdnd11an1n16x5 FILLER_328_2134 ();
 b15zdnd11an1n04x5 FILLER_328_2150 ();
 b15zdnd11an1n64x5 FILLER_328_2162 ();
 b15zdnd11an1n32x5 FILLER_328_2226 ();
 b15zdnd11an1n16x5 FILLER_328_2258 ();
 b15zdnd00an1n02x5 FILLER_328_2274 ();
 b15zdnd11an1n64x5 FILLER_329_0 ();
 b15zdnd11an1n64x5 FILLER_329_64 ();
 b15zdnd11an1n64x5 FILLER_329_128 ();
 b15zdnd11an1n64x5 FILLER_329_192 ();
 b15zdnd11an1n64x5 FILLER_329_256 ();
 b15zdnd11an1n64x5 FILLER_329_320 ();
 b15zdnd11an1n64x5 FILLER_329_384 ();
 b15zdnd11an1n64x5 FILLER_329_448 ();
 b15zdnd11an1n64x5 FILLER_329_512 ();
 b15zdnd11an1n64x5 FILLER_329_576 ();
 b15zdnd11an1n64x5 FILLER_329_640 ();
 b15zdnd11an1n64x5 FILLER_329_704 ();
 b15zdnd11an1n64x5 FILLER_329_768 ();
 b15zdnd11an1n64x5 FILLER_329_832 ();
 b15zdnd11an1n64x5 FILLER_329_896 ();
 b15zdnd11an1n64x5 FILLER_329_960 ();
 b15zdnd11an1n64x5 FILLER_329_1024 ();
 b15zdnd11an1n64x5 FILLER_329_1088 ();
 b15zdnd11an1n64x5 FILLER_329_1152 ();
 b15zdnd11an1n64x5 FILLER_329_1216 ();
 b15zdnd11an1n64x5 FILLER_329_1280 ();
 b15zdnd11an1n64x5 FILLER_329_1344 ();
 b15zdnd11an1n64x5 FILLER_329_1408 ();
 b15zdnd11an1n64x5 FILLER_329_1472 ();
 b15zdnd11an1n64x5 FILLER_329_1536 ();
 b15zdnd11an1n64x5 FILLER_329_1600 ();
 b15zdnd11an1n64x5 FILLER_329_1664 ();
 b15zdnd11an1n64x5 FILLER_329_1728 ();
 b15zdnd11an1n64x5 FILLER_329_1792 ();
 b15zdnd11an1n32x5 FILLER_329_1856 ();
 b15zdnd11an1n16x5 FILLER_329_1888 ();
 b15zdnd11an1n08x5 FILLER_329_1904 ();
 b15zdnd11an1n04x5 FILLER_329_1912 ();
 b15zdnd00an1n02x5 FILLER_329_1916 ();
 b15zdnd00an1n01x5 FILLER_329_1918 ();
 b15zdnd11an1n64x5 FILLER_329_1928 ();
 b15zdnd11an1n64x5 FILLER_329_1992 ();
 b15zdnd11an1n64x5 FILLER_329_2056 ();
 b15zdnd11an1n64x5 FILLER_329_2120 ();
 b15zdnd11an1n64x5 FILLER_329_2184 ();
 b15zdnd11an1n32x5 FILLER_329_2248 ();
 b15zdnd11an1n04x5 FILLER_329_2280 ();
 b15zdnd11an1n64x5 FILLER_330_8 ();
 b15zdnd11an1n64x5 FILLER_330_72 ();
 b15zdnd11an1n64x5 FILLER_330_136 ();
 b15zdnd11an1n64x5 FILLER_330_200 ();
 b15zdnd11an1n64x5 FILLER_330_264 ();
 b15zdnd11an1n64x5 FILLER_330_328 ();
 b15zdnd11an1n64x5 FILLER_330_392 ();
 b15zdnd11an1n64x5 FILLER_330_456 ();
 b15zdnd11an1n64x5 FILLER_330_520 ();
 b15zdnd11an1n64x5 FILLER_330_584 ();
 b15zdnd11an1n64x5 FILLER_330_648 ();
 b15zdnd11an1n04x5 FILLER_330_712 ();
 b15zdnd00an1n02x5 FILLER_330_716 ();
 b15zdnd11an1n64x5 FILLER_330_726 ();
 b15zdnd11an1n64x5 FILLER_330_790 ();
 b15zdnd11an1n64x5 FILLER_330_854 ();
 b15zdnd11an1n64x5 FILLER_330_918 ();
 b15zdnd11an1n64x5 FILLER_330_982 ();
 b15zdnd11an1n64x5 FILLER_330_1046 ();
 b15zdnd11an1n64x5 FILLER_330_1110 ();
 b15zdnd11an1n64x5 FILLER_330_1174 ();
 b15zdnd11an1n64x5 FILLER_330_1238 ();
 b15zdnd11an1n64x5 FILLER_330_1302 ();
 b15zdnd11an1n64x5 FILLER_330_1366 ();
 b15zdnd11an1n64x5 FILLER_330_1430 ();
 b15zdnd11an1n64x5 FILLER_330_1494 ();
 b15zdnd11an1n64x5 FILLER_330_1558 ();
 b15zdnd11an1n64x5 FILLER_330_1622 ();
 b15zdnd11an1n64x5 FILLER_330_1686 ();
 b15zdnd11an1n64x5 FILLER_330_1750 ();
 b15zdnd11an1n64x5 FILLER_330_1814 ();
 b15zdnd11an1n64x5 FILLER_330_1878 ();
 b15zdnd11an1n64x5 FILLER_330_1942 ();
 b15zdnd11an1n64x5 FILLER_330_2006 ();
 b15zdnd11an1n64x5 FILLER_330_2070 ();
 b15zdnd11an1n16x5 FILLER_330_2134 ();
 b15zdnd11an1n04x5 FILLER_330_2150 ();
 b15zdnd11an1n64x5 FILLER_330_2162 ();
 b15zdnd11an1n32x5 FILLER_330_2226 ();
 b15zdnd11an1n16x5 FILLER_330_2258 ();
 b15zdnd00an1n02x5 FILLER_330_2274 ();
 b15zdnd11an1n64x5 FILLER_331_0 ();
 b15zdnd11an1n64x5 FILLER_331_64 ();
 b15zdnd11an1n64x5 FILLER_331_128 ();
 b15zdnd11an1n64x5 FILLER_331_192 ();
 b15zdnd11an1n64x5 FILLER_331_256 ();
 b15zdnd11an1n64x5 FILLER_331_320 ();
 b15zdnd11an1n64x5 FILLER_331_384 ();
 b15zdnd11an1n64x5 FILLER_331_448 ();
 b15zdnd11an1n64x5 FILLER_331_512 ();
 b15zdnd11an1n64x5 FILLER_331_576 ();
 b15zdnd11an1n64x5 FILLER_331_640 ();
 b15zdnd11an1n64x5 FILLER_331_704 ();
 b15zdnd11an1n64x5 FILLER_331_768 ();
 b15zdnd11an1n64x5 FILLER_331_832 ();
 b15zdnd11an1n64x5 FILLER_331_896 ();
 b15zdnd11an1n64x5 FILLER_331_960 ();
 b15zdnd11an1n64x5 FILLER_331_1024 ();
 b15zdnd11an1n64x5 FILLER_331_1088 ();
 b15zdnd11an1n64x5 FILLER_331_1152 ();
 b15zdnd11an1n64x5 FILLER_331_1216 ();
 b15zdnd11an1n64x5 FILLER_331_1280 ();
 b15zdnd11an1n64x5 FILLER_331_1344 ();
 b15zdnd11an1n64x5 FILLER_331_1408 ();
 b15zdnd11an1n64x5 FILLER_331_1472 ();
 b15zdnd11an1n64x5 FILLER_331_1536 ();
 b15zdnd11an1n64x5 FILLER_331_1600 ();
 b15zdnd11an1n64x5 FILLER_331_1664 ();
 b15zdnd11an1n64x5 FILLER_331_1728 ();
 b15zdnd11an1n64x5 FILLER_331_1792 ();
 b15zdnd11an1n64x5 FILLER_331_1856 ();
 b15zdnd11an1n64x5 FILLER_331_1920 ();
 b15zdnd11an1n64x5 FILLER_331_1984 ();
 b15zdnd11an1n64x5 FILLER_331_2048 ();
 b15zdnd11an1n64x5 FILLER_331_2112 ();
 b15zdnd11an1n64x5 FILLER_331_2176 ();
 b15zdnd11an1n32x5 FILLER_331_2240 ();
 b15zdnd11an1n08x5 FILLER_331_2272 ();
 b15zdnd11an1n04x5 FILLER_331_2280 ();
 b15zdnd11an1n64x5 FILLER_332_8 ();
 b15zdnd11an1n64x5 FILLER_332_72 ();
 b15zdnd11an1n64x5 FILLER_332_136 ();
 b15zdnd11an1n64x5 FILLER_332_200 ();
 b15zdnd11an1n64x5 FILLER_332_264 ();
 b15zdnd11an1n64x5 FILLER_332_328 ();
 b15zdnd11an1n64x5 FILLER_332_392 ();
 b15zdnd11an1n64x5 FILLER_332_456 ();
 b15zdnd11an1n64x5 FILLER_332_520 ();
 b15zdnd11an1n64x5 FILLER_332_584 ();
 b15zdnd11an1n64x5 FILLER_332_648 ();
 b15zdnd11an1n04x5 FILLER_332_712 ();
 b15zdnd00an1n02x5 FILLER_332_716 ();
 b15zdnd11an1n64x5 FILLER_332_726 ();
 b15zdnd11an1n64x5 FILLER_332_790 ();
 b15zdnd11an1n64x5 FILLER_332_854 ();
 b15zdnd11an1n64x5 FILLER_332_918 ();
 b15zdnd11an1n64x5 FILLER_332_982 ();
 b15zdnd11an1n64x5 FILLER_332_1046 ();
 b15zdnd11an1n64x5 FILLER_332_1110 ();
 b15zdnd11an1n64x5 FILLER_332_1174 ();
 b15zdnd11an1n64x5 FILLER_332_1238 ();
 b15zdnd11an1n64x5 FILLER_332_1302 ();
 b15zdnd11an1n64x5 FILLER_332_1366 ();
 b15zdnd11an1n64x5 FILLER_332_1430 ();
 b15zdnd11an1n64x5 FILLER_332_1494 ();
 b15zdnd11an1n64x5 FILLER_332_1558 ();
 b15zdnd11an1n64x5 FILLER_332_1622 ();
 b15zdnd11an1n64x5 FILLER_332_1686 ();
 b15zdnd11an1n64x5 FILLER_332_1750 ();
 b15zdnd11an1n64x5 FILLER_332_1814 ();
 b15zdnd11an1n64x5 FILLER_332_1878 ();
 b15zdnd11an1n64x5 FILLER_332_1942 ();
 b15zdnd11an1n64x5 FILLER_332_2006 ();
 b15zdnd11an1n64x5 FILLER_332_2070 ();
 b15zdnd11an1n16x5 FILLER_332_2134 ();
 b15zdnd11an1n04x5 FILLER_332_2150 ();
 b15zdnd11an1n64x5 FILLER_332_2162 ();
 b15zdnd11an1n32x5 FILLER_332_2226 ();
 b15zdnd11an1n16x5 FILLER_332_2258 ();
 b15zdnd00an1n02x5 FILLER_332_2274 ();
 b15zdnd11an1n64x5 FILLER_333_0 ();
 b15zdnd11an1n64x5 FILLER_333_64 ();
 b15zdnd11an1n64x5 FILLER_333_128 ();
 b15zdnd11an1n64x5 FILLER_333_192 ();
 b15zdnd11an1n64x5 FILLER_333_256 ();
 b15zdnd11an1n64x5 FILLER_333_320 ();
 b15zdnd11an1n64x5 FILLER_333_384 ();
 b15zdnd11an1n64x5 FILLER_333_448 ();
 b15zdnd11an1n64x5 FILLER_333_512 ();
 b15zdnd11an1n64x5 FILLER_333_576 ();
 b15zdnd11an1n64x5 FILLER_333_640 ();
 b15zdnd11an1n64x5 FILLER_333_704 ();
 b15zdnd11an1n64x5 FILLER_333_768 ();
 b15zdnd11an1n64x5 FILLER_333_832 ();
 b15zdnd11an1n64x5 FILLER_333_896 ();
 b15zdnd11an1n64x5 FILLER_333_960 ();
 b15zdnd11an1n64x5 FILLER_333_1024 ();
 b15zdnd11an1n64x5 FILLER_333_1088 ();
 b15zdnd11an1n64x5 FILLER_333_1152 ();
 b15zdnd11an1n64x5 FILLER_333_1216 ();
 b15zdnd11an1n64x5 FILLER_333_1280 ();
 b15zdnd11an1n64x5 FILLER_333_1344 ();
 b15zdnd11an1n64x5 FILLER_333_1408 ();
 b15zdnd11an1n64x5 FILLER_333_1472 ();
 b15zdnd11an1n64x5 FILLER_333_1536 ();
 b15zdnd11an1n64x5 FILLER_333_1600 ();
 b15zdnd11an1n64x5 FILLER_333_1664 ();
 b15zdnd11an1n64x5 FILLER_333_1728 ();
 b15zdnd11an1n64x5 FILLER_333_1792 ();
 b15zdnd11an1n64x5 FILLER_333_1856 ();
 b15zdnd11an1n64x5 FILLER_333_1920 ();
 b15zdnd11an1n64x5 FILLER_333_1984 ();
 b15zdnd11an1n64x5 FILLER_333_2048 ();
 b15zdnd11an1n64x5 FILLER_333_2112 ();
 b15zdnd11an1n64x5 FILLER_333_2176 ();
 b15zdnd11an1n32x5 FILLER_333_2240 ();
 b15zdnd11an1n08x5 FILLER_333_2272 ();
 b15zdnd11an1n04x5 FILLER_333_2280 ();
 b15zdnd11an1n64x5 FILLER_334_8 ();
 b15zdnd11an1n64x5 FILLER_334_72 ();
 b15zdnd11an1n64x5 FILLER_334_136 ();
 b15zdnd11an1n64x5 FILLER_334_200 ();
 b15zdnd11an1n64x5 FILLER_334_264 ();
 b15zdnd11an1n64x5 FILLER_334_328 ();
 b15zdnd11an1n64x5 FILLER_334_392 ();
 b15zdnd11an1n64x5 FILLER_334_456 ();
 b15zdnd11an1n64x5 FILLER_334_520 ();
 b15zdnd11an1n64x5 FILLER_334_584 ();
 b15zdnd11an1n64x5 FILLER_334_648 ();
 b15zdnd11an1n04x5 FILLER_334_712 ();
 b15zdnd00an1n02x5 FILLER_334_716 ();
 b15zdnd11an1n64x5 FILLER_334_726 ();
 b15zdnd11an1n64x5 FILLER_334_790 ();
 b15zdnd11an1n64x5 FILLER_334_854 ();
 b15zdnd11an1n64x5 FILLER_334_918 ();
 b15zdnd11an1n64x5 FILLER_334_982 ();
 b15zdnd11an1n64x5 FILLER_334_1046 ();
 b15zdnd11an1n64x5 FILLER_334_1110 ();
 b15zdnd11an1n64x5 FILLER_334_1174 ();
 b15zdnd11an1n64x5 FILLER_334_1238 ();
 b15zdnd11an1n64x5 FILLER_334_1302 ();
 b15zdnd11an1n64x5 FILLER_334_1366 ();
 b15zdnd11an1n64x5 FILLER_334_1430 ();
 b15zdnd11an1n64x5 FILLER_334_1494 ();
 b15zdnd11an1n64x5 FILLER_334_1558 ();
 b15zdnd11an1n64x5 FILLER_334_1622 ();
 b15zdnd11an1n64x5 FILLER_334_1686 ();
 b15zdnd11an1n64x5 FILLER_334_1750 ();
 b15zdnd11an1n64x5 FILLER_334_1814 ();
 b15zdnd11an1n64x5 FILLER_334_1878 ();
 b15zdnd11an1n64x5 FILLER_334_1942 ();
 b15zdnd11an1n64x5 FILLER_334_2006 ();
 b15zdnd11an1n64x5 FILLER_334_2070 ();
 b15zdnd11an1n16x5 FILLER_334_2134 ();
 b15zdnd11an1n04x5 FILLER_334_2150 ();
 b15zdnd11an1n64x5 FILLER_334_2162 ();
 b15zdnd11an1n32x5 FILLER_334_2226 ();
 b15zdnd11an1n16x5 FILLER_334_2258 ();
 b15zdnd00an1n02x5 FILLER_334_2274 ();
 b15zdnd11an1n64x5 FILLER_335_0 ();
 b15zdnd11an1n64x5 FILLER_335_64 ();
 b15zdnd11an1n64x5 FILLER_335_128 ();
 b15zdnd11an1n64x5 FILLER_335_192 ();
 b15zdnd11an1n64x5 FILLER_335_256 ();
 b15zdnd11an1n64x5 FILLER_335_320 ();
 b15zdnd11an1n64x5 FILLER_335_384 ();
 b15zdnd11an1n64x5 FILLER_335_448 ();
 b15zdnd11an1n64x5 FILLER_335_512 ();
 b15zdnd11an1n64x5 FILLER_335_576 ();
 b15zdnd11an1n64x5 FILLER_335_640 ();
 b15zdnd11an1n64x5 FILLER_335_704 ();
 b15zdnd11an1n64x5 FILLER_335_768 ();
 b15zdnd11an1n64x5 FILLER_335_832 ();
 b15zdnd11an1n64x5 FILLER_335_896 ();
 b15zdnd11an1n64x5 FILLER_335_960 ();
 b15zdnd11an1n64x5 FILLER_335_1024 ();
 b15zdnd11an1n64x5 FILLER_335_1088 ();
 b15zdnd11an1n64x5 FILLER_335_1152 ();
 b15zdnd11an1n64x5 FILLER_335_1216 ();
 b15zdnd11an1n64x5 FILLER_335_1280 ();
 b15zdnd11an1n64x5 FILLER_335_1344 ();
 b15zdnd11an1n64x5 FILLER_335_1408 ();
 b15zdnd11an1n64x5 FILLER_335_1472 ();
 b15zdnd11an1n64x5 FILLER_335_1536 ();
 b15zdnd11an1n64x5 FILLER_335_1600 ();
 b15zdnd11an1n64x5 FILLER_335_1664 ();
 b15zdnd11an1n64x5 FILLER_335_1728 ();
 b15zdnd11an1n64x5 FILLER_335_1792 ();
 b15zdnd11an1n64x5 FILLER_335_1856 ();
 b15zdnd11an1n64x5 FILLER_335_1920 ();
 b15zdnd11an1n64x5 FILLER_335_1984 ();
 b15zdnd11an1n64x5 FILLER_335_2048 ();
 b15zdnd11an1n64x5 FILLER_335_2112 ();
 b15zdnd11an1n64x5 FILLER_335_2176 ();
 b15zdnd11an1n32x5 FILLER_335_2240 ();
 b15zdnd11an1n08x5 FILLER_335_2272 ();
 b15zdnd11an1n04x5 FILLER_335_2280 ();
 b15zdnd11an1n64x5 FILLER_336_8 ();
 b15zdnd11an1n64x5 FILLER_336_72 ();
 b15zdnd11an1n64x5 FILLER_336_136 ();
 b15zdnd11an1n64x5 FILLER_336_200 ();
 b15zdnd11an1n64x5 FILLER_336_264 ();
 b15zdnd11an1n64x5 FILLER_336_328 ();
 b15zdnd11an1n64x5 FILLER_336_392 ();
 b15zdnd11an1n64x5 FILLER_336_456 ();
 b15zdnd11an1n64x5 FILLER_336_520 ();
 b15zdnd11an1n64x5 FILLER_336_584 ();
 b15zdnd11an1n64x5 FILLER_336_648 ();
 b15zdnd11an1n04x5 FILLER_336_712 ();
 b15zdnd00an1n02x5 FILLER_336_716 ();
 b15zdnd11an1n64x5 FILLER_336_726 ();
 b15zdnd11an1n64x5 FILLER_336_790 ();
 b15zdnd11an1n64x5 FILLER_336_854 ();
 b15zdnd11an1n64x5 FILLER_336_918 ();
 b15zdnd11an1n64x5 FILLER_336_982 ();
 b15zdnd11an1n64x5 FILLER_336_1046 ();
 b15zdnd11an1n64x5 FILLER_336_1110 ();
 b15zdnd11an1n64x5 FILLER_336_1174 ();
 b15zdnd11an1n64x5 FILLER_336_1238 ();
 b15zdnd11an1n64x5 FILLER_336_1302 ();
 b15zdnd11an1n64x5 FILLER_336_1366 ();
 b15zdnd11an1n64x5 FILLER_336_1430 ();
 b15zdnd11an1n64x5 FILLER_336_1494 ();
 b15zdnd11an1n64x5 FILLER_336_1558 ();
 b15zdnd11an1n64x5 FILLER_336_1622 ();
 b15zdnd11an1n64x5 FILLER_336_1686 ();
 b15zdnd11an1n64x5 FILLER_336_1750 ();
 b15zdnd11an1n64x5 FILLER_336_1814 ();
 b15zdnd11an1n64x5 FILLER_336_1878 ();
 b15zdnd11an1n64x5 FILLER_336_1942 ();
 b15zdnd11an1n64x5 FILLER_336_2006 ();
 b15zdnd11an1n64x5 FILLER_336_2070 ();
 b15zdnd11an1n16x5 FILLER_336_2134 ();
 b15zdnd11an1n04x5 FILLER_336_2150 ();
 b15zdnd11an1n64x5 FILLER_336_2162 ();
 b15zdnd11an1n32x5 FILLER_336_2226 ();
 b15zdnd11an1n16x5 FILLER_336_2258 ();
 b15zdnd00an1n02x5 FILLER_336_2274 ();
 b15zdnd11an1n64x5 FILLER_337_0 ();
 b15zdnd11an1n64x5 FILLER_337_64 ();
 b15zdnd11an1n64x5 FILLER_337_128 ();
 b15zdnd11an1n64x5 FILLER_337_192 ();
 b15zdnd11an1n64x5 FILLER_337_256 ();
 b15zdnd11an1n64x5 FILLER_337_320 ();
 b15zdnd11an1n64x5 FILLER_337_384 ();
 b15zdnd11an1n64x5 FILLER_337_448 ();
 b15zdnd11an1n64x5 FILLER_337_512 ();
 b15zdnd11an1n64x5 FILLER_337_576 ();
 b15zdnd11an1n64x5 FILLER_337_640 ();
 b15zdnd11an1n64x5 FILLER_337_704 ();
 b15zdnd11an1n64x5 FILLER_337_768 ();
 b15zdnd11an1n64x5 FILLER_337_832 ();
 b15zdnd11an1n64x5 FILLER_337_896 ();
 b15zdnd11an1n64x5 FILLER_337_960 ();
 b15zdnd11an1n64x5 FILLER_337_1024 ();
 b15zdnd11an1n64x5 FILLER_337_1088 ();
 b15zdnd11an1n64x5 FILLER_337_1152 ();
 b15zdnd11an1n64x5 FILLER_337_1216 ();
 b15zdnd11an1n64x5 FILLER_337_1280 ();
 b15zdnd11an1n64x5 FILLER_337_1344 ();
 b15zdnd11an1n64x5 FILLER_337_1408 ();
 b15zdnd11an1n64x5 FILLER_337_1472 ();
 b15zdnd11an1n64x5 FILLER_337_1536 ();
 b15zdnd11an1n64x5 FILLER_337_1600 ();
 b15zdnd11an1n64x5 FILLER_337_1664 ();
 b15zdnd11an1n64x5 FILLER_337_1728 ();
 b15zdnd11an1n64x5 FILLER_337_1792 ();
 b15zdnd11an1n64x5 FILLER_337_1856 ();
 b15zdnd11an1n64x5 FILLER_337_1920 ();
 b15zdnd11an1n64x5 FILLER_337_1984 ();
 b15zdnd11an1n64x5 FILLER_337_2048 ();
 b15zdnd11an1n64x5 FILLER_337_2112 ();
 b15zdnd11an1n64x5 FILLER_337_2176 ();
 b15zdnd11an1n32x5 FILLER_337_2240 ();
 b15zdnd11an1n08x5 FILLER_337_2272 ();
 b15zdnd11an1n04x5 FILLER_337_2280 ();
 b15zdnd11an1n64x5 FILLER_338_8 ();
 b15zdnd11an1n64x5 FILLER_338_72 ();
 b15zdnd11an1n64x5 FILLER_338_136 ();
 b15zdnd11an1n64x5 FILLER_338_200 ();
 b15zdnd11an1n64x5 FILLER_338_264 ();
 b15zdnd11an1n64x5 FILLER_338_328 ();
 b15zdnd11an1n64x5 FILLER_338_392 ();
 b15zdnd11an1n64x5 FILLER_338_456 ();
 b15zdnd11an1n64x5 FILLER_338_520 ();
 b15zdnd11an1n64x5 FILLER_338_584 ();
 b15zdnd11an1n64x5 FILLER_338_648 ();
 b15zdnd11an1n04x5 FILLER_338_712 ();
 b15zdnd00an1n02x5 FILLER_338_716 ();
 b15zdnd11an1n64x5 FILLER_338_726 ();
 b15zdnd11an1n64x5 FILLER_338_790 ();
 b15zdnd11an1n64x5 FILLER_338_854 ();
 b15zdnd11an1n64x5 FILLER_338_918 ();
 b15zdnd11an1n64x5 FILLER_338_982 ();
 b15zdnd11an1n64x5 FILLER_338_1046 ();
 b15zdnd11an1n64x5 FILLER_338_1110 ();
 b15zdnd11an1n64x5 FILLER_338_1174 ();
 b15zdnd11an1n64x5 FILLER_338_1238 ();
 b15zdnd11an1n64x5 FILLER_338_1302 ();
 b15zdnd11an1n64x5 FILLER_338_1366 ();
 b15zdnd11an1n64x5 FILLER_338_1430 ();
 b15zdnd11an1n64x5 FILLER_338_1494 ();
 b15zdnd11an1n64x5 FILLER_338_1558 ();
 b15zdnd11an1n64x5 FILLER_338_1622 ();
 b15zdnd11an1n64x5 FILLER_338_1686 ();
 b15zdnd11an1n64x5 FILLER_338_1750 ();
 b15zdnd11an1n64x5 FILLER_338_1814 ();
 b15zdnd11an1n64x5 FILLER_338_1878 ();
 b15zdnd11an1n64x5 FILLER_338_1942 ();
 b15zdnd11an1n64x5 FILLER_338_2006 ();
 b15zdnd11an1n64x5 FILLER_338_2070 ();
 b15zdnd11an1n16x5 FILLER_338_2134 ();
 b15zdnd11an1n04x5 FILLER_338_2150 ();
 b15zdnd11an1n64x5 FILLER_338_2162 ();
 b15zdnd11an1n32x5 FILLER_338_2226 ();
 b15zdnd11an1n16x5 FILLER_338_2258 ();
 b15zdnd00an1n02x5 FILLER_338_2274 ();
 b15zdnd11an1n64x5 FILLER_339_0 ();
 b15zdnd11an1n64x5 FILLER_339_64 ();
 b15zdnd11an1n64x5 FILLER_339_128 ();
 b15zdnd11an1n64x5 FILLER_339_192 ();
 b15zdnd11an1n64x5 FILLER_339_256 ();
 b15zdnd11an1n64x5 FILLER_339_320 ();
 b15zdnd11an1n64x5 FILLER_339_384 ();
 b15zdnd11an1n64x5 FILLER_339_448 ();
 b15zdnd11an1n64x5 FILLER_339_512 ();
 b15zdnd11an1n64x5 FILLER_339_576 ();
 b15zdnd11an1n64x5 FILLER_339_640 ();
 b15zdnd11an1n64x5 FILLER_339_704 ();
 b15zdnd11an1n64x5 FILLER_339_768 ();
 b15zdnd11an1n64x5 FILLER_339_832 ();
 b15zdnd11an1n64x5 FILLER_339_896 ();
 b15zdnd11an1n64x5 FILLER_339_960 ();
 b15zdnd11an1n64x5 FILLER_339_1024 ();
 b15zdnd11an1n64x5 FILLER_339_1088 ();
 b15zdnd11an1n64x5 FILLER_339_1152 ();
 b15zdnd11an1n64x5 FILLER_339_1216 ();
 b15zdnd11an1n64x5 FILLER_339_1280 ();
 b15zdnd11an1n64x5 FILLER_339_1344 ();
 b15zdnd11an1n64x5 FILLER_339_1408 ();
 b15zdnd11an1n64x5 FILLER_339_1472 ();
 b15zdnd11an1n64x5 FILLER_339_1536 ();
 b15zdnd11an1n64x5 FILLER_339_1600 ();
 b15zdnd11an1n64x5 FILLER_339_1664 ();
 b15zdnd11an1n64x5 FILLER_339_1728 ();
 b15zdnd11an1n64x5 FILLER_339_1792 ();
 b15zdnd11an1n64x5 FILLER_339_1856 ();
 b15zdnd11an1n64x5 FILLER_339_1920 ();
 b15zdnd11an1n64x5 FILLER_339_1984 ();
 b15zdnd11an1n64x5 FILLER_339_2048 ();
 b15zdnd11an1n64x5 FILLER_339_2112 ();
 b15zdnd11an1n64x5 FILLER_339_2176 ();
 b15zdnd11an1n32x5 FILLER_339_2240 ();
 b15zdnd11an1n08x5 FILLER_339_2272 ();
 b15zdnd11an1n04x5 FILLER_339_2280 ();
 b15zdnd11an1n64x5 FILLER_340_8 ();
 b15zdnd11an1n64x5 FILLER_340_72 ();
 b15zdnd11an1n64x5 FILLER_340_136 ();
 b15zdnd11an1n64x5 FILLER_340_200 ();
 b15zdnd11an1n64x5 FILLER_340_264 ();
 b15zdnd11an1n64x5 FILLER_340_328 ();
 b15zdnd11an1n64x5 FILLER_340_392 ();
 b15zdnd11an1n64x5 FILLER_340_456 ();
 b15zdnd11an1n64x5 FILLER_340_520 ();
 b15zdnd11an1n64x5 FILLER_340_584 ();
 b15zdnd11an1n64x5 FILLER_340_648 ();
 b15zdnd11an1n04x5 FILLER_340_712 ();
 b15zdnd00an1n02x5 FILLER_340_716 ();
 b15zdnd11an1n64x5 FILLER_340_726 ();
 b15zdnd11an1n64x5 FILLER_340_790 ();
 b15zdnd11an1n64x5 FILLER_340_854 ();
 b15zdnd11an1n64x5 FILLER_340_918 ();
 b15zdnd11an1n64x5 FILLER_340_982 ();
 b15zdnd11an1n64x5 FILLER_340_1046 ();
 b15zdnd11an1n64x5 FILLER_340_1110 ();
 b15zdnd11an1n64x5 FILLER_340_1174 ();
 b15zdnd11an1n64x5 FILLER_340_1238 ();
 b15zdnd11an1n64x5 FILLER_340_1302 ();
 b15zdnd11an1n64x5 FILLER_340_1366 ();
 b15zdnd11an1n64x5 FILLER_340_1430 ();
 b15zdnd11an1n64x5 FILLER_340_1494 ();
 b15zdnd11an1n64x5 FILLER_340_1558 ();
 b15zdnd11an1n64x5 FILLER_340_1622 ();
 b15zdnd11an1n64x5 FILLER_340_1686 ();
 b15zdnd11an1n64x5 FILLER_340_1750 ();
 b15zdnd11an1n64x5 FILLER_340_1814 ();
 b15zdnd11an1n64x5 FILLER_340_1878 ();
 b15zdnd11an1n64x5 FILLER_340_1942 ();
 b15zdnd11an1n64x5 FILLER_340_2006 ();
 b15zdnd11an1n64x5 FILLER_340_2070 ();
 b15zdnd11an1n16x5 FILLER_340_2134 ();
 b15zdnd11an1n04x5 FILLER_340_2150 ();
 b15zdnd11an1n64x5 FILLER_340_2162 ();
 b15zdnd11an1n32x5 FILLER_340_2226 ();
 b15zdnd11an1n16x5 FILLER_340_2258 ();
 b15zdnd00an1n02x5 FILLER_340_2274 ();
 b15zdnd11an1n64x5 FILLER_341_0 ();
 b15zdnd11an1n64x5 FILLER_341_64 ();
 b15zdnd11an1n64x5 FILLER_341_128 ();
 b15zdnd11an1n64x5 FILLER_341_192 ();
 b15zdnd11an1n64x5 FILLER_341_256 ();
 b15zdnd11an1n64x5 FILLER_341_320 ();
 b15zdnd11an1n64x5 FILLER_341_384 ();
 b15zdnd11an1n64x5 FILLER_341_448 ();
 b15zdnd11an1n64x5 FILLER_341_512 ();
 b15zdnd11an1n64x5 FILLER_341_576 ();
 b15zdnd11an1n64x5 FILLER_341_640 ();
 b15zdnd11an1n64x5 FILLER_341_704 ();
 b15zdnd11an1n64x5 FILLER_341_768 ();
 b15zdnd11an1n64x5 FILLER_341_832 ();
 b15zdnd11an1n64x5 FILLER_341_896 ();
 b15zdnd11an1n64x5 FILLER_341_960 ();
 b15zdnd11an1n64x5 FILLER_341_1024 ();
 b15zdnd11an1n64x5 FILLER_341_1088 ();
 b15zdnd11an1n64x5 FILLER_341_1152 ();
 b15zdnd11an1n64x5 FILLER_341_1216 ();
 b15zdnd11an1n64x5 FILLER_341_1280 ();
 b15zdnd11an1n64x5 FILLER_341_1344 ();
 b15zdnd11an1n64x5 FILLER_341_1408 ();
 b15zdnd11an1n64x5 FILLER_341_1472 ();
 b15zdnd11an1n64x5 FILLER_341_1536 ();
 b15zdnd11an1n64x5 FILLER_341_1600 ();
 b15zdnd11an1n64x5 FILLER_341_1664 ();
 b15zdnd11an1n64x5 FILLER_341_1728 ();
 b15zdnd11an1n64x5 FILLER_341_1792 ();
 b15zdnd11an1n64x5 FILLER_341_1856 ();
 b15zdnd11an1n64x5 FILLER_341_1920 ();
 b15zdnd11an1n64x5 FILLER_341_1984 ();
 b15zdnd11an1n64x5 FILLER_341_2048 ();
 b15zdnd11an1n64x5 FILLER_341_2112 ();
 b15zdnd11an1n64x5 FILLER_341_2176 ();
 b15zdnd11an1n32x5 FILLER_341_2240 ();
 b15zdnd11an1n08x5 FILLER_341_2272 ();
 b15zdnd11an1n04x5 FILLER_341_2280 ();
 b15zdnd11an1n64x5 FILLER_342_8 ();
 b15zdnd11an1n64x5 FILLER_342_72 ();
 b15zdnd11an1n64x5 FILLER_342_136 ();
 b15zdnd11an1n64x5 FILLER_342_200 ();
 b15zdnd11an1n64x5 FILLER_342_264 ();
 b15zdnd11an1n64x5 FILLER_342_328 ();
 b15zdnd11an1n64x5 FILLER_342_392 ();
 b15zdnd11an1n64x5 FILLER_342_456 ();
 b15zdnd11an1n64x5 FILLER_342_520 ();
 b15zdnd11an1n64x5 FILLER_342_584 ();
 b15zdnd11an1n64x5 FILLER_342_648 ();
 b15zdnd11an1n04x5 FILLER_342_712 ();
 b15zdnd00an1n02x5 FILLER_342_716 ();
 b15zdnd11an1n64x5 FILLER_342_726 ();
 b15zdnd11an1n64x5 FILLER_342_790 ();
 b15zdnd11an1n64x5 FILLER_342_854 ();
 b15zdnd11an1n64x5 FILLER_342_918 ();
 b15zdnd11an1n64x5 FILLER_342_982 ();
 b15zdnd11an1n64x5 FILLER_342_1046 ();
 b15zdnd11an1n64x5 FILLER_342_1110 ();
 b15zdnd11an1n64x5 FILLER_342_1174 ();
 b15zdnd11an1n64x5 FILLER_342_1238 ();
 b15zdnd11an1n64x5 FILLER_342_1302 ();
 b15zdnd11an1n64x5 FILLER_342_1366 ();
 b15zdnd11an1n64x5 FILLER_342_1430 ();
 b15zdnd11an1n64x5 FILLER_342_1494 ();
 b15zdnd11an1n64x5 FILLER_342_1558 ();
 b15zdnd11an1n64x5 FILLER_342_1622 ();
 b15zdnd11an1n64x5 FILLER_342_1686 ();
 b15zdnd11an1n64x5 FILLER_342_1750 ();
 b15zdnd11an1n64x5 FILLER_342_1814 ();
 b15zdnd11an1n64x5 FILLER_342_1878 ();
 b15zdnd11an1n64x5 FILLER_342_1942 ();
 b15zdnd11an1n64x5 FILLER_342_2006 ();
 b15zdnd11an1n64x5 FILLER_342_2070 ();
 b15zdnd11an1n16x5 FILLER_342_2134 ();
 b15zdnd11an1n04x5 FILLER_342_2150 ();
 b15zdnd11an1n64x5 FILLER_342_2162 ();
 b15zdnd11an1n32x5 FILLER_342_2226 ();
 b15zdnd11an1n16x5 FILLER_342_2258 ();
 b15zdnd00an1n02x5 FILLER_342_2274 ();
 b15zdnd11an1n64x5 FILLER_343_0 ();
 b15zdnd11an1n64x5 FILLER_343_64 ();
 b15zdnd11an1n64x5 FILLER_343_128 ();
 b15zdnd11an1n64x5 FILLER_343_192 ();
 b15zdnd11an1n64x5 FILLER_343_256 ();
 b15zdnd11an1n64x5 FILLER_343_320 ();
 b15zdnd11an1n64x5 FILLER_343_384 ();
 b15zdnd11an1n64x5 FILLER_343_448 ();
 b15zdnd11an1n64x5 FILLER_343_512 ();
 b15zdnd11an1n64x5 FILLER_343_576 ();
 b15zdnd11an1n64x5 FILLER_343_640 ();
 b15zdnd11an1n64x5 FILLER_343_704 ();
 b15zdnd11an1n64x5 FILLER_343_768 ();
 b15zdnd11an1n64x5 FILLER_343_832 ();
 b15zdnd11an1n64x5 FILLER_343_896 ();
 b15zdnd11an1n64x5 FILLER_343_960 ();
 b15zdnd11an1n64x5 FILLER_343_1024 ();
 b15zdnd11an1n64x5 FILLER_343_1088 ();
 b15zdnd11an1n64x5 FILLER_343_1152 ();
 b15zdnd11an1n64x5 FILLER_343_1216 ();
 b15zdnd11an1n64x5 FILLER_343_1280 ();
 b15zdnd11an1n64x5 FILLER_343_1344 ();
 b15zdnd11an1n64x5 FILLER_343_1408 ();
 b15zdnd11an1n64x5 FILLER_343_1472 ();
 b15zdnd11an1n64x5 FILLER_343_1536 ();
 b15zdnd11an1n64x5 FILLER_343_1600 ();
 b15zdnd11an1n64x5 FILLER_343_1664 ();
 b15zdnd11an1n64x5 FILLER_343_1728 ();
 b15zdnd11an1n64x5 FILLER_343_1792 ();
 b15zdnd11an1n64x5 FILLER_343_1856 ();
 b15zdnd11an1n64x5 FILLER_343_1920 ();
 b15zdnd11an1n64x5 FILLER_343_1984 ();
 b15zdnd11an1n64x5 FILLER_343_2048 ();
 b15zdnd11an1n64x5 FILLER_343_2112 ();
 b15zdnd11an1n64x5 FILLER_343_2176 ();
 b15zdnd11an1n32x5 FILLER_343_2240 ();
 b15zdnd11an1n08x5 FILLER_343_2272 ();
 b15zdnd11an1n04x5 FILLER_343_2280 ();
 b15zdnd11an1n64x5 FILLER_344_8 ();
 b15zdnd11an1n64x5 FILLER_344_72 ();
 b15zdnd11an1n64x5 FILLER_344_136 ();
 b15zdnd11an1n64x5 FILLER_344_200 ();
 b15zdnd11an1n64x5 FILLER_344_264 ();
 b15zdnd11an1n64x5 FILLER_344_328 ();
 b15zdnd11an1n64x5 FILLER_344_392 ();
 b15zdnd11an1n64x5 FILLER_344_456 ();
 b15zdnd11an1n64x5 FILLER_344_520 ();
 b15zdnd11an1n64x5 FILLER_344_584 ();
 b15zdnd11an1n64x5 FILLER_344_648 ();
 b15zdnd11an1n04x5 FILLER_344_712 ();
 b15zdnd00an1n02x5 FILLER_344_716 ();
 b15zdnd11an1n64x5 FILLER_344_726 ();
 b15zdnd11an1n64x5 FILLER_344_790 ();
 b15zdnd11an1n64x5 FILLER_344_854 ();
 b15zdnd11an1n64x5 FILLER_344_918 ();
 b15zdnd11an1n64x5 FILLER_344_982 ();
 b15zdnd11an1n64x5 FILLER_344_1046 ();
 b15zdnd11an1n64x5 FILLER_344_1110 ();
 b15zdnd11an1n64x5 FILLER_344_1174 ();
 b15zdnd11an1n64x5 FILLER_344_1238 ();
 b15zdnd11an1n64x5 FILLER_344_1302 ();
 b15zdnd11an1n64x5 FILLER_344_1366 ();
 b15zdnd11an1n64x5 FILLER_344_1430 ();
 b15zdnd11an1n64x5 FILLER_344_1494 ();
 b15zdnd11an1n64x5 FILLER_344_1558 ();
 b15zdnd11an1n64x5 FILLER_344_1622 ();
 b15zdnd11an1n64x5 FILLER_344_1686 ();
 b15zdnd11an1n64x5 FILLER_344_1750 ();
 b15zdnd11an1n64x5 FILLER_344_1814 ();
 b15zdnd11an1n64x5 FILLER_344_1878 ();
 b15zdnd11an1n64x5 FILLER_344_1942 ();
 b15zdnd11an1n64x5 FILLER_344_2006 ();
 b15zdnd11an1n64x5 FILLER_344_2070 ();
 b15zdnd11an1n16x5 FILLER_344_2134 ();
 b15zdnd11an1n04x5 FILLER_344_2150 ();
 b15zdnd11an1n64x5 FILLER_344_2162 ();
 b15zdnd11an1n32x5 FILLER_344_2226 ();
 b15zdnd11an1n16x5 FILLER_344_2258 ();
 b15zdnd00an1n02x5 FILLER_344_2274 ();
 b15zdnd11an1n64x5 FILLER_345_0 ();
 b15zdnd11an1n64x5 FILLER_345_64 ();
 b15zdnd11an1n64x5 FILLER_345_128 ();
 b15zdnd11an1n64x5 FILLER_345_192 ();
 b15zdnd11an1n64x5 FILLER_345_256 ();
 b15zdnd11an1n64x5 FILLER_345_320 ();
 b15zdnd11an1n64x5 FILLER_345_384 ();
 b15zdnd11an1n64x5 FILLER_345_448 ();
 b15zdnd11an1n64x5 FILLER_345_512 ();
 b15zdnd11an1n64x5 FILLER_345_576 ();
 b15zdnd11an1n64x5 FILLER_345_640 ();
 b15zdnd11an1n64x5 FILLER_345_704 ();
 b15zdnd11an1n64x5 FILLER_345_768 ();
 b15zdnd11an1n64x5 FILLER_345_832 ();
 b15zdnd11an1n64x5 FILLER_345_896 ();
 b15zdnd11an1n64x5 FILLER_345_960 ();
 b15zdnd11an1n64x5 FILLER_345_1024 ();
 b15zdnd11an1n64x5 FILLER_345_1088 ();
 b15zdnd11an1n64x5 FILLER_345_1152 ();
 b15zdnd11an1n64x5 FILLER_345_1216 ();
 b15zdnd11an1n64x5 FILLER_345_1280 ();
 b15zdnd11an1n64x5 FILLER_345_1344 ();
 b15zdnd11an1n64x5 FILLER_345_1408 ();
 b15zdnd11an1n64x5 FILLER_345_1472 ();
 b15zdnd11an1n64x5 FILLER_345_1536 ();
 b15zdnd11an1n64x5 FILLER_345_1600 ();
 b15zdnd11an1n64x5 FILLER_345_1664 ();
 b15zdnd11an1n64x5 FILLER_345_1728 ();
 b15zdnd11an1n64x5 FILLER_345_1792 ();
 b15zdnd11an1n64x5 FILLER_345_1856 ();
 b15zdnd11an1n64x5 FILLER_345_1920 ();
 b15zdnd11an1n64x5 FILLER_345_1984 ();
 b15zdnd11an1n64x5 FILLER_345_2048 ();
 b15zdnd11an1n64x5 FILLER_345_2112 ();
 b15zdnd11an1n64x5 FILLER_345_2176 ();
 b15zdnd11an1n32x5 FILLER_345_2240 ();
 b15zdnd11an1n08x5 FILLER_345_2272 ();
 b15zdnd11an1n04x5 FILLER_345_2280 ();
 b15zdnd11an1n64x5 FILLER_346_8 ();
 b15zdnd11an1n64x5 FILLER_346_72 ();
 b15zdnd11an1n64x5 FILLER_346_136 ();
 b15zdnd11an1n64x5 FILLER_346_200 ();
 b15zdnd11an1n64x5 FILLER_346_264 ();
 b15zdnd11an1n64x5 FILLER_346_328 ();
 b15zdnd11an1n64x5 FILLER_346_392 ();
 b15zdnd11an1n64x5 FILLER_346_456 ();
 b15zdnd11an1n64x5 FILLER_346_520 ();
 b15zdnd11an1n64x5 FILLER_346_584 ();
 b15zdnd11an1n64x5 FILLER_346_648 ();
 b15zdnd11an1n04x5 FILLER_346_712 ();
 b15zdnd00an1n02x5 FILLER_346_716 ();
 b15zdnd11an1n64x5 FILLER_346_726 ();
 b15zdnd11an1n64x5 FILLER_346_790 ();
 b15zdnd11an1n64x5 FILLER_346_854 ();
 b15zdnd11an1n64x5 FILLER_346_918 ();
 b15zdnd11an1n64x5 FILLER_346_982 ();
 b15zdnd11an1n64x5 FILLER_346_1046 ();
 b15zdnd11an1n64x5 FILLER_346_1110 ();
 b15zdnd11an1n64x5 FILLER_346_1174 ();
 b15zdnd11an1n64x5 FILLER_346_1238 ();
 b15zdnd11an1n64x5 FILLER_346_1302 ();
 b15zdnd11an1n64x5 FILLER_346_1366 ();
 b15zdnd11an1n64x5 FILLER_346_1430 ();
 b15zdnd11an1n64x5 FILLER_346_1494 ();
 b15zdnd11an1n64x5 FILLER_346_1558 ();
 b15zdnd11an1n64x5 FILLER_346_1622 ();
 b15zdnd11an1n64x5 FILLER_346_1686 ();
 b15zdnd11an1n64x5 FILLER_346_1750 ();
 b15zdnd11an1n64x5 FILLER_346_1814 ();
 b15zdnd11an1n64x5 FILLER_346_1878 ();
 b15zdnd11an1n64x5 FILLER_346_1942 ();
 b15zdnd11an1n64x5 FILLER_346_2006 ();
 b15zdnd11an1n64x5 FILLER_346_2070 ();
 b15zdnd11an1n16x5 FILLER_346_2134 ();
 b15zdnd11an1n04x5 FILLER_346_2150 ();
 b15zdnd11an1n64x5 FILLER_346_2162 ();
 b15zdnd11an1n32x5 FILLER_346_2226 ();
 b15zdnd11an1n16x5 FILLER_346_2258 ();
 b15zdnd00an1n02x5 FILLER_346_2274 ();
 b15zdnd11an1n64x5 FILLER_347_0 ();
 b15zdnd11an1n64x5 FILLER_347_64 ();
 b15zdnd11an1n64x5 FILLER_347_128 ();
 b15zdnd11an1n64x5 FILLER_347_192 ();
 b15zdnd11an1n64x5 FILLER_347_256 ();
 b15zdnd11an1n64x5 FILLER_347_320 ();
 b15zdnd11an1n64x5 FILLER_347_384 ();
 b15zdnd11an1n64x5 FILLER_347_448 ();
 b15zdnd11an1n64x5 FILLER_347_512 ();
 b15zdnd11an1n64x5 FILLER_347_576 ();
 b15zdnd11an1n64x5 FILLER_347_640 ();
 b15zdnd11an1n64x5 FILLER_347_704 ();
 b15zdnd11an1n64x5 FILLER_347_768 ();
 b15zdnd11an1n64x5 FILLER_347_832 ();
 b15zdnd11an1n64x5 FILLER_347_896 ();
 b15zdnd11an1n64x5 FILLER_347_960 ();
 b15zdnd11an1n64x5 FILLER_347_1024 ();
 b15zdnd11an1n64x5 FILLER_347_1088 ();
 b15zdnd11an1n64x5 FILLER_347_1152 ();
 b15zdnd11an1n64x5 FILLER_347_1216 ();
 b15zdnd11an1n64x5 FILLER_347_1280 ();
 b15zdnd11an1n64x5 FILLER_347_1344 ();
 b15zdnd11an1n64x5 FILLER_347_1408 ();
 b15zdnd11an1n64x5 FILLER_347_1472 ();
 b15zdnd11an1n64x5 FILLER_347_1536 ();
 b15zdnd11an1n64x5 FILLER_347_1600 ();
 b15zdnd11an1n64x5 FILLER_347_1664 ();
 b15zdnd11an1n64x5 FILLER_347_1728 ();
 b15zdnd11an1n64x5 FILLER_347_1792 ();
 b15zdnd11an1n64x5 FILLER_347_1856 ();
 b15zdnd11an1n64x5 FILLER_347_1920 ();
 b15zdnd11an1n64x5 FILLER_347_1984 ();
 b15zdnd11an1n64x5 FILLER_347_2048 ();
 b15zdnd11an1n64x5 FILLER_347_2112 ();
 b15zdnd11an1n64x5 FILLER_347_2176 ();
 b15zdnd11an1n32x5 FILLER_347_2240 ();
 b15zdnd11an1n08x5 FILLER_347_2272 ();
 b15zdnd11an1n04x5 FILLER_347_2280 ();
 b15zdnd11an1n64x5 FILLER_348_8 ();
 b15zdnd11an1n64x5 FILLER_348_72 ();
 b15zdnd11an1n64x5 FILLER_348_136 ();
 b15zdnd11an1n64x5 FILLER_348_200 ();
 b15zdnd11an1n64x5 FILLER_348_264 ();
 b15zdnd11an1n64x5 FILLER_348_328 ();
 b15zdnd11an1n64x5 FILLER_348_392 ();
 b15zdnd11an1n64x5 FILLER_348_456 ();
 b15zdnd11an1n64x5 FILLER_348_520 ();
 b15zdnd11an1n64x5 FILLER_348_584 ();
 b15zdnd11an1n64x5 FILLER_348_648 ();
 b15zdnd11an1n04x5 FILLER_348_712 ();
 b15zdnd00an1n02x5 FILLER_348_716 ();
 b15zdnd11an1n64x5 FILLER_348_726 ();
 b15zdnd11an1n64x5 FILLER_348_790 ();
 b15zdnd11an1n64x5 FILLER_348_854 ();
 b15zdnd11an1n64x5 FILLER_348_918 ();
 b15zdnd11an1n64x5 FILLER_348_982 ();
 b15zdnd11an1n64x5 FILLER_348_1046 ();
 b15zdnd11an1n64x5 FILLER_348_1110 ();
 b15zdnd11an1n64x5 FILLER_348_1174 ();
 b15zdnd11an1n64x5 FILLER_348_1238 ();
 b15zdnd11an1n64x5 FILLER_348_1302 ();
 b15zdnd11an1n64x5 FILLER_348_1366 ();
 b15zdnd11an1n64x5 FILLER_348_1430 ();
 b15zdnd11an1n64x5 FILLER_348_1494 ();
 b15zdnd11an1n64x5 FILLER_348_1558 ();
 b15zdnd11an1n64x5 FILLER_348_1622 ();
 b15zdnd11an1n64x5 FILLER_348_1686 ();
 b15zdnd11an1n64x5 FILLER_348_1750 ();
 b15zdnd11an1n64x5 FILLER_348_1814 ();
 b15zdnd11an1n64x5 FILLER_348_1878 ();
 b15zdnd11an1n64x5 FILLER_348_1942 ();
 b15zdnd11an1n64x5 FILLER_348_2006 ();
 b15zdnd11an1n64x5 FILLER_348_2070 ();
 b15zdnd11an1n16x5 FILLER_348_2134 ();
 b15zdnd11an1n04x5 FILLER_348_2150 ();
 b15zdnd11an1n64x5 FILLER_348_2162 ();
 b15zdnd11an1n32x5 FILLER_348_2226 ();
 b15zdnd11an1n16x5 FILLER_348_2258 ();
 b15zdnd00an1n02x5 FILLER_348_2274 ();
 b15zdnd11an1n64x5 FILLER_349_0 ();
 b15zdnd11an1n64x5 FILLER_349_64 ();
 b15zdnd11an1n64x5 FILLER_349_128 ();
 b15zdnd11an1n64x5 FILLER_349_192 ();
 b15zdnd11an1n64x5 FILLER_349_256 ();
 b15zdnd11an1n64x5 FILLER_349_320 ();
 b15zdnd11an1n64x5 FILLER_349_384 ();
 b15zdnd11an1n64x5 FILLER_349_448 ();
 b15zdnd11an1n64x5 FILLER_349_512 ();
 b15zdnd11an1n64x5 FILLER_349_576 ();
 b15zdnd11an1n64x5 FILLER_349_640 ();
 b15zdnd11an1n64x5 FILLER_349_704 ();
 b15zdnd11an1n64x5 FILLER_349_768 ();
 b15zdnd11an1n64x5 FILLER_349_832 ();
 b15zdnd11an1n64x5 FILLER_349_896 ();
 b15zdnd11an1n64x5 FILLER_349_960 ();
 b15zdnd11an1n64x5 FILLER_349_1024 ();
 b15zdnd11an1n64x5 FILLER_349_1088 ();
 b15zdnd11an1n64x5 FILLER_349_1152 ();
 b15zdnd11an1n64x5 FILLER_349_1216 ();
 b15zdnd11an1n64x5 FILLER_349_1280 ();
 b15zdnd11an1n64x5 FILLER_349_1344 ();
 b15zdnd11an1n64x5 FILLER_349_1408 ();
 b15zdnd11an1n64x5 FILLER_349_1472 ();
 b15zdnd11an1n64x5 FILLER_349_1536 ();
 b15zdnd11an1n64x5 FILLER_349_1600 ();
 b15zdnd11an1n64x5 FILLER_349_1664 ();
 b15zdnd11an1n64x5 FILLER_349_1728 ();
 b15zdnd11an1n64x5 FILLER_349_1792 ();
 b15zdnd11an1n64x5 FILLER_349_1856 ();
 b15zdnd11an1n64x5 FILLER_349_1920 ();
 b15zdnd11an1n64x5 FILLER_349_1984 ();
 b15zdnd11an1n64x5 FILLER_349_2048 ();
 b15zdnd11an1n64x5 FILLER_349_2112 ();
 b15zdnd11an1n64x5 FILLER_349_2176 ();
 b15zdnd11an1n32x5 FILLER_349_2240 ();
 b15zdnd11an1n08x5 FILLER_349_2272 ();
 b15zdnd11an1n04x5 FILLER_349_2280 ();
 b15zdnd11an1n64x5 FILLER_350_8 ();
 b15zdnd11an1n64x5 FILLER_350_72 ();
 b15zdnd11an1n64x5 FILLER_350_136 ();
 b15zdnd11an1n64x5 FILLER_350_200 ();
 b15zdnd11an1n64x5 FILLER_350_264 ();
 b15zdnd11an1n64x5 FILLER_350_328 ();
 b15zdnd11an1n64x5 FILLER_350_392 ();
 b15zdnd11an1n64x5 FILLER_350_456 ();
 b15zdnd11an1n64x5 FILLER_350_520 ();
 b15zdnd11an1n64x5 FILLER_350_584 ();
 b15zdnd11an1n64x5 FILLER_350_648 ();
 b15zdnd11an1n04x5 FILLER_350_712 ();
 b15zdnd00an1n02x5 FILLER_350_716 ();
 b15zdnd11an1n64x5 FILLER_350_726 ();
 b15zdnd11an1n64x5 FILLER_350_790 ();
 b15zdnd11an1n64x5 FILLER_350_854 ();
 b15zdnd11an1n64x5 FILLER_350_918 ();
 b15zdnd11an1n64x5 FILLER_350_982 ();
 b15zdnd11an1n64x5 FILLER_350_1046 ();
 b15zdnd11an1n64x5 FILLER_350_1110 ();
 b15zdnd11an1n64x5 FILLER_350_1174 ();
 b15zdnd11an1n64x5 FILLER_350_1238 ();
 b15zdnd11an1n64x5 FILLER_350_1302 ();
 b15zdnd11an1n64x5 FILLER_350_1366 ();
 b15zdnd11an1n64x5 FILLER_350_1430 ();
 b15zdnd11an1n64x5 FILLER_350_1494 ();
 b15zdnd11an1n64x5 FILLER_350_1558 ();
 b15zdnd11an1n64x5 FILLER_350_1622 ();
 b15zdnd11an1n64x5 FILLER_350_1686 ();
 b15zdnd11an1n64x5 FILLER_350_1750 ();
 b15zdnd11an1n64x5 FILLER_350_1814 ();
 b15zdnd11an1n64x5 FILLER_350_1878 ();
 b15zdnd11an1n64x5 FILLER_350_1942 ();
 b15zdnd11an1n64x5 FILLER_350_2006 ();
 b15zdnd11an1n64x5 FILLER_350_2070 ();
 b15zdnd11an1n16x5 FILLER_350_2134 ();
 b15zdnd11an1n04x5 FILLER_350_2150 ();
 b15zdnd11an1n64x5 FILLER_350_2162 ();
 b15zdnd11an1n32x5 FILLER_350_2226 ();
 b15zdnd11an1n16x5 FILLER_350_2258 ();
 b15zdnd00an1n02x5 FILLER_350_2274 ();
 b15zdnd11an1n64x5 FILLER_351_0 ();
 b15zdnd11an1n64x5 FILLER_351_64 ();
 b15zdnd11an1n64x5 FILLER_351_128 ();
 b15zdnd11an1n64x5 FILLER_351_192 ();
 b15zdnd11an1n64x5 FILLER_351_256 ();
 b15zdnd11an1n64x5 FILLER_351_320 ();
 b15zdnd11an1n64x5 FILLER_351_384 ();
 b15zdnd11an1n64x5 FILLER_351_448 ();
 b15zdnd11an1n64x5 FILLER_351_512 ();
 b15zdnd11an1n64x5 FILLER_351_576 ();
 b15zdnd11an1n64x5 FILLER_351_640 ();
 b15zdnd11an1n64x5 FILLER_351_704 ();
 b15zdnd11an1n64x5 FILLER_351_768 ();
 b15zdnd11an1n64x5 FILLER_351_832 ();
 b15zdnd11an1n64x5 FILLER_351_896 ();
 b15zdnd11an1n64x5 FILLER_351_960 ();
 b15zdnd11an1n64x5 FILLER_351_1024 ();
 b15zdnd11an1n64x5 FILLER_351_1088 ();
 b15zdnd11an1n64x5 FILLER_351_1152 ();
 b15zdnd11an1n64x5 FILLER_351_1216 ();
 b15zdnd11an1n64x5 FILLER_351_1280 ();
 b15zdnd11an1n64x5 FILLER_351_1344 ();
 b15zdnd11an1n64x5 FILLER_351_1408 ();
 b15zdnd11an1n64x5 FILLER_351_1472 ();
 b15zdnd11an1n64x5 FILLER_351_1536 ();
 b15zdnd11an1n64x5 FILLER_351_1600 ();
 b15zdnd11an1n64x5 FILLER_351_1664 ();
 b15zdnd11an1n64x5 FILLER_351_1728 ();
 b15zdnd11an1n64x5 FILLER_351_1792 ();
 b15zdnd11an1n64x5 FILLER_351_1856 ();
 b15zdnd11an1n64x5 FILLER_351_1920 ();
 b15zdnd11an1n64x5 FILLER_351_1984 ();
 b15zdnd11an1n64x5 FILLER_351_2048 ();
 b15zdnd11an1n64x5 FILLER_351_2112 ();
 b15zdnd11an1n64x5 FILLER_351_2176 ();
 b15zdnd11an1n32x5 FILLER_351_2240 ();
 b15zdnd11an1n08x5 FILLER_351_2272 ();
 b15zdnd11an1n04x5 FILLER_351_2280 ();
 b15zdnd11an1n64x5 FILLER_352_8 ();
 b15zdnd11an1n64x5 FILLER_352_72 ();
 b15zdnd11an1n64x5 FILLER_352_136 ();
 b15zdnd11an1n64x5 FILLER_352_200 ();
 b15zdnd11an1n64x5 FILLER_352_264 ();
 b15zdnd11an1n64x5 FILLER_352_328 ();
 b15zdnd11an1n64x5 FILLER_352_392 ();
 b15zdnd11an1n64x5 FILLER_352_456 ();
 b15zdnd11an1n64x5 FILLER_352_520 ();
 b15zdnd11an1n64x5 FILLER_352_584 ();
 b15zdnd11an1n64x5 FILLER_352_648 ();
 b15zdnd11an1n04x5 FILLER_352_712 ();
 b15zdnd00an1n02x5 FILLER_352_716 ();
 b15zdnd11an1n64x5 FILLER_352_726 ();
 b15zdnd11an1n64x5 FILLER_352_790 ();
 b15zdnd11an1n64x5 FILLER_352_854 ();
 b15zdnd11an1n64x5 FILLER_352_918 ();
 b15zdnd11an1n64x5 FILLER_352_982 ();
 b15zdnd11an1n64x5 FILLER_352_1046 ();
 b15zdnd11an1n64x5 FILLER_352_1110 ();
 b15zdnd11an1n64x5 FILLER_352_1174 ();
 b15zdnd11an1n64x5 FILLER_352_1238 ();
 b15zdnd11an1n64x5 FILLER_352_1302 ();
 b15zdnd11an1n64x5 FILLER_352_1366 ();
 b15zdnd11an1n64x5 FILLER_352_1430 ();
 b15zdnd11an1n64x5 FILLER_352_1494 ();
 b15zdnd11an1n64x5 FILLER_352_1558 ();
 b15zdnd11an1n64x5 FILLER_352_1622 ();
 b15zdnd11an1n64x5 FILLER_352_1686 ();
 b15zdnd11an1n64x5 FILLER_352_1750 ();
 b15zdnd11an1n64x5 FILLER_352_1814 ();
 b15zdnd11an1n64x5 FILLER_352_1878 ();
 b15zdnd11an1n64x5 FILLER_352_1942 ();
 b15zdnd11an1n64x5 FILLER_352_2006 ();
 b15zdnd11an1n64x5 FILLER_352_2070 ();
 b15zdnd11an1n16x5 FILLER_352_2134 ();
 b15zdnd11an1n04x5 FILLER_352_2150 ();
 b15zdnd11an1n64x5 FILLER_352_2162 ();
 b15zdnd11an1n32x5 FILLER_352_2226 ();
 b15zdnd11an1n16x5 FILLER_352_2258 ();
 b15zdnd00an1n02x5 FILLER_352_2274 ();
 b15zdnd11an1n64x5 FILLER_353_0 ();
 b15zdnd11an1n64x5 FILLER_353_64 ();
 b15zdnd11an1n64x5 FILLER_353_128 ();
 b15zdnd11an1n64x5 FILLER_353_192 ();
 b15zdnd11an1n64x5 FILLER_353_256 ();
 b15zdnd11an1n64x5 FILLER_353_320 ();
 b15zdnd11an1n64x5 FILLER_353_384 ();
 b15zdnd11an1n64x5 FILLER_353_448 ();
 b15zdnd11an1n64x5 FILLER_353_512 ();
 b15zdnd11an1n64x5 FILLER_353_576 ();
 b15zdnd11an1n64x5 FILLER_353_640 ();
 b15zdnd11an1n64x5 FILLER_353_704 ();
 b15zdnd11an1n64x5 FILLER_353_768 ();
 b15zdnd11an1n64x5 FILLER_353_832 ();
 b15zdnd11an1n64x5 FILLER_353_896 ();
 b15zdnd11an1n64x5 FILLER_353_960 ();
 b15zdnd11an1n64x5 FILLER_353_1024 ();
 b15zdnd11an1n64x5 FILLER_353_1088 ();
 b15zdnd11an1n64x5 FILLER_353_1152 ();
 b15zdnd11an1n64x5 FILLER_353_1216 ();
 b15zdnd11an1n64x5 FILLER_353_1280 ();
 b15zdnd11an1n64x5 FILLER_353_1344 ();
 b15zdnd11an1n64x5 FILLER_353_1408 ();
 b15zdnd11an1n64x5 FILLER_353_1472 ();
 b15zdnd11an1n64x5 FILLER_353_1536 ();
 b15zdnd11an1n64x5 FILLER_353_1600 ();
 b15zdnd11an1n64x5 FILLER_353_1664 ();
 b15zdnd11an1n64x5 FILLER_353_1728 ();
 b15zdnd11an1n64x5 FILLER_353_1792 ();
 b15zdnd11an1n64x5 FILLER_353_1856 ();
 b15zdnd11an1n64x5 FILLER_353_1920 ();
 b15zdnd11an1n64x5 FILLER_353_1984 ();
 b15zdnd11an1n64x5 FILLER_353_2048 ();
 b15zdnd11an1n64x5 FILLER_353_2112 ();
 b15zdnd11an1n64x5 FILLER_353_2176 ();
 b15zdnd11an1n32x5 FILLER_353_2240 ();
 b15zdnd11an1n08x5 FILLER_353_2272 ();
 b15zdnd11an1n04x5 FILLER_353_2280 ();
 b15zdnd11an1n64x5 FILLER_354_8 ();
 b15zdnd11an1n64x5 FILLER_354_72 ();
 b15zdnd11an1n64x5 FILLER_354_136 ();
 b15zdnd11an1n64x5 FILLER_354_200 ();
 b15zdnd11an1n64x5 FILLER_354_264 ();
 b15zdnd11an1n64x5 FILLER_354_328 ();
 b15zdnd11an1n64x5 FILLER_354_392 ();
 b15zdnd11an1n64x5 FILLER_354_456 ();
 b15zdnd11an1n64x5 FILLER_354_520 ();
 b15zdnd11an1n64x5 FILLER_354_584 ();
 b15zdnd11an1n64x5 FILLER_354_648 ();
 b15zdnd11an1n04x5 FILLER_354_712 ();
 b15zdnd00an1n02x5 FILLER_354_716 ();
 b15zdnd11an1n64x5 FILLER_354_726 ();
 b15zdnd11an1n64x5 FILLER_354_790 ();
 b15zdnd11an1n64x5 FILLER_354_854 ();
 b15zdnd11an1n64x5 FILLER_354_918 ();
 b15zdnd11an1n64x5 FILLER_354_982 ();
 b15zdnd11an1n64x5 FILLER_354_1046 ();
 b15zdnd11an1n64x5 FILLER_354_1110 ();
 b15zdnd11an1n64x5 FILLER_354_1174 ();
 b15zdnd11an1n64x5 FILLER_354_1238 ();
 b15zdnd11an1n64x5 FILLER_354_1302 ();
 b15zdnd11an1n64x5 FILLER_354_1366 ();
 b15zdnd11an1n64x5 FILLER_354_1430 ();
 b15zdnd11an1n64x5 FILLER_354_1494 ();
 b15zdnd11an1n64x5 FILLER_354_1558 ();
 b15zdnd11an1n64x5 FILLER_354_1622 ();
 b15zdnd11an1n64x5 FILLER_354_1686 ();
 b15zdnd11an1n64x5 FILLER_354_1750 ();
 b15zdnd11an1n64x5 FILLER_354_1814 ();
 b15zdnd11an1n64x5 FILLER_354_1878 ();
 b15zdnd11an1n64x5 FILLER_354_1942 ();
 b15zdnd11an1n64x5 FILLER_354_2006 ();
 b15zdnd11an1n64x5 FILLER_354_2070 ();
 b15zdnd11an1n16x5 FILLER_354_2134 ();
 b15zdnd11an1n04x5 FILLER_354_2150 ();
 b15zdnd11an1n64x5 FILLER_354_2162 ();
 b15zdnd11an1n32x5 FILLER_354_2226 ();
 b15zdnd11an1n16x5 FILLER_354_2258 ();
 b15zdnd00an1n02x5 FILLER_354_2274 ();
 b15zdnd11an1n64x5 FILLER_355_0 ();
 b15zdnd11an1n64x5 FILLER_355_64 ();
 b15zdnd11an1n64x5 FILLER_355_128 ();
 b15zdnd11an1n64x5 FILLER_355_192 ();
 b15zdnd11an1n64x5 FILLER_355_256 ();
 b15zdnd11an1n64x5 FILLER_355_320 ();
 b15zdnd11an1n64x5 FILLER_355_384 ();
 b15zdnd11an1n64x5 FILLER_355_448 ();
 b15zdnd11an1n64x5 FILLER_355_512 ();
 b15zdnd11an1n64x5 FILLER_355_576 ();
 b15zdnd11an1n64x5 FILLER_355_640 ();
 b15zdnd11an1n64x5 FILLER_355_704 ();
 b15zdnd11an1n64x5 FILLER_355_768 ();
 b15zdnd11an1n64x5 FILLER_355_832 ();
 b15zdnd11an1n64x5 FILLER_355_896 ();
 b15zdnd11an1n64x5 FILLER_355_960 ();
 b15zdnd11an1n64x5 FILLER_355_1024 ();
 b15zdnd11an1n64x5 FILLER_355_1088 ();
 b15zdnd11an1n64x5 FILLER_355_1152 ();
 b15zdnd11an1n64x5 FILLER_355_1216 ();
 b15zdnd11an1n64x5 FILLER_355_1280 ();
 b15zdnd11an1n64x5 FILLER_355_1344 ();
 b15zdnd11an1n64x5 FILLER_355_1408 ();
 b15zdnd11an1n64x5 FILLER_355_1472 ();
 b15zdnd11an1n64x5 FILLER_355_1536 ();
 b15zdnd11an1n64x5 FILLER_355_1600 ();
 b15zdnd11an1n64x5 FILLER_355_1664 ();
 b15zdnd11an1n64x5 FILLER_355_1728 ();
 b15zdnd11an1n64x5 FILLER_355_1792 ();
 b15zdnd11an1n64x5 FILLER_355_1856 ();
 b15zdnd11an1n64x5 FILLER_355_1920 ();
 b15zdnd11an1n64x5 FILLER_355_1984 ();
 b15zdnd11an1n64x5 FILLER_355_2048 ();
 b15zdnd11an1n64x5 FILLER_355_2112 ();
 b15zdnd11an1n64x5 FILLER_355_2176 ();
 b15zdnd11an1n32x5 FILLER_355_2240 ();
 b15zdnd11an1n08x5 FILLER_355_2272 ();
 b15zdnd11an1n04x5 FILLER_355_2280 ();
 b15zdnd11an1n64x5 FILLER_356_8 ();
 b15zdnd11an1n64x5 FILLER_356_72 ();
 b15zdnd11an1n64x5 FILLER_356_136 ();
 b15zdnd11an1n64x5 FILLER_356_200 ();
 b15zdnd11an1n64x5 FILLER_356_264 ();
 b15zdnd11an1n64x5 FILLER_356_328 ();
 b15zdnd11an1n64x5 FILLER_356_392 ();
 b15zdnd11an1n64x5 FILLER_356_456 ();
 b15zdnd11an1n64x5 FILLER_356_520 ();
 b15zdnd11an1n64x5 FILLER_356_584 ();
 b15zdnd11an1n64x5 FILLER_356_648 ();
 b15zdnd11an1n04x5 FILLER_356_712 ();
 b15zdnd00an1n02x5 FILLER_356_716 ();
 b15zdnd11an1n64x5 FILLER_356_726 ();
 b15zdnd11an1n64x5 FILLER_356_790 ();
 b15zdnd11an1n64x5 FILLER_356_854 ();
 b15zdnd11an1n64x5 FILLER_356_918 ();
 b15zdnd11an1n64x5 FILLER_356_982 ();
 b15zdnd11an1n64x5 FILLER_356_1046 ();
 b15zdnd11an1n64x5 FILLER_356_1110 ();
 b15zdnd11an1n64x5 FILLER_356_1174 ();
 b15zdnd11an1n64x5 FILLER_356_1238 ();
 b15zdnd11an1n64x5 FILLER_356_1302 ();
 b15zdnd11an1n64x5 FILLER_356_1366 ();
 b15zdnd11an1n64x5 FILLER_356_1430 ();
 b15zdnd11an1n64x5 FILLER_356_1494 ();
 b15zdnd11an1n64x5 FILLER_356_1558 ();
 b15zdnd11an1n64x5 FILLER_356_1622 ();
 b15zdnd11an1n64x5 FILLER_356_1686 ();
 b15zdnd11an1n64x5 FILLER_356_1750 ();
 b15zdnd11an1n64x5 FILLER_356_1814 ();
 b15zdnd11an1n64x5 FILLER_356_1878 ();
 b15zdnd11an1n64x5 FILLER_356_1942 ();
 b15zdnd11an1n64x5 FILLER_356_2006 ();
 b15zdnd11an1n64x5 FILLER_356_2070 ();
 b15zdnd11an1n16x5 FILLER_356_2134 ();
 b15zdnd11an1n04x5 FILLER_356_2150 ();
 b15zdnd11an1n64x5 FILLER_356_2162 ();
 b15zdnd11an1n32x5 FILLER_356_2226 ();
 b15zdnd11an1n16x5 FILLER_356_2258 ();
 b15zdnd00an1n02x5 FILLER_356_2274 ();
 b15zdnd11an1n64x5 FILLER_357_0 ();
 b15zdnd11an1n64x5 FILLER_357_64 ();
 b15zdnd11an1n64x5 FILLER_357_128 ();
 b15zdnd11an1n64x5 FILLER_357_192 ();
 b15zdnd11an1n64x5 FILLER_357_256 ();
 b15zdnd11an1n64x5 FILLER_357_320 ();
 b15zdnd11an1n64x5 FILLER_357_384 ();
 b15zdnd11an1n64x5 FILLER_357_448 ();
 b15zdnd11an1n64x5 FILLER_357_512 ();
 b15zdnd11an1n64x5 FILLER_357_576 ();
 b15zdnd11an1n64x5 FILLER_357_640 ();
 b15zdnd11an1n64x5 FILLER_357_704 ();
 b15zdnd11an1n64x5 FILLER_357_768 ();
 b15zdnd11an1n64x5 FILLER_357_832 ();
 b15zdnd11an1n64x5 FILLER_357_896 ();
 b15zdnd11an1n64x5 FILLER_357_960 ();
 b15zdnd11an1n64x5 FILLER_357_1024 ();
 b15zdnd11an1n64x5 FILLER_357_1088 ();
 b15zdnd11an1n64x5 FILLER_357_1152 ();
 b15zdnd11an1n64x5 FILLER_357_1216 ();
 b15zdnd11an1n64x5 FILLER_357_1280 ();
 b15zdnd11an1n64x5 FILLER_357_1344 ();
 b15zdnd11an1n64x5 FILLER_357_1408 ();
 b15zdnd11an1n64x5 FILLER_357_1472 ();
 b15zdnd11an1n64x5 FILLER_357_1536 ();
 b15zdnd11an1n64x5 FILLER_357_1600 ();
 b15zdnd11an1n64x5 FILLER_357_1664 ();
 b15zdnd11an1n64x5 FILLER_357_1728 ();
 b15zdnd11an1n64x5 FILLER_357_1792 ();
 b15zdnd11an1n64x5 FILLER_357_1856 ();
 b15zdnd11an1n64x5 FILLER_357_1920 ();
 b15zdnd11an1n64x5 FILLER_357_1984 ();
 b15zdnd11an1n64x5 FILLER_357_2048 ();
 b15zdnd11an1n64x5 FILLER_357_2112 ();
 b15zdnd11an1n64x5 FILLER_357_2176 ();
 b15zdnd11an1n32x5 FILLER_357_2240 ();
 b15zdnd11an1n08x5 FILLER_357_2272 ();
 b15zdnd11an1n04x5 FILLER_357_2280 ();
 b15zdnd11an1n64x5 FILLER_358_8 ();
 b15zdnd11an1n64x5 FILLER_358_72 ();
 b15zdnd11an1n64x5 FILLER_358_136 ();
 b15zdnd11an1n64x5 FILLER_358_200 ();
 b15zdnd11an1n64x5 FILLER_358_264 ();
 b15zdnd11an1n64x5 FILLER_358_328 ();
 b15zdnd11an1n64x5 FILLER_358_392 ();
 b15zdnd11an1n64x5 FILLER_358_456 ();
 b15zdnd11an1n64x5 FILLER_358_520 ();
 b15zdnd11an1n64x5 FILLER_358_584 ();
 b15zdnd11an1n64x5 FILLER_358_648 ();
 b15zdnd11an1n04x5 FILLER_358_712 ();
 b15zdnd00an1n02x5 FILLER_358_716 ();
 b15zdnd11an1n64x5 FILLER_358_726 ();
 b15zdnd11an1n64x5 FILLER_358_790 ();
 b15zdnd11an1n64x5 FILLER_358_854 ();
 b15zdnd11an1n64x5 FILLER_358_918 ();
 b15zdnd11an1n64x5 FILLER_358_982 ();
 b15zdnd11an1n64x5 FILLER_358_1046 ();
 b15zdnd11an1n64x5 FILLER_358_1110 ();
 b15zdnd11an1n64x5 FILLER_358_1174 ();
 b15zdnd11an1n64x5 FILLER_358_1238 ();
 b15zdnd11an1n64x5 FILLER_358_1302 ();
 b15zdnd11an1n64x5 FILLER_358_1366 ();
 b15zdnd11an1n64x5 FILLER_358_1430 ();
 b15zdnd11an1n64x5 FILLER_358_1494 ();
 b15zdnd11an1n64x5 FILLER_358_1558 ();
 b15zdnd11an1n64x5 FILLER_358_1622 ();
 b15zdnd11an1n64x5 FILLER_358_1686 ();
 b15zdnd11an1n64x5 FILLER_358_1750 ();
 b15zdnd11an1n64x5 FILLER_358_1814 ();
 b15zdnd11an1n64x5 FILLER_358_1878 ();
 b15zdnd11an1n64x5 FILLER_358_1942 ();
 b15zdnd11an1n64x5 FILLER_358_2006 ();
 b15zdnd11an1n64x5 FILLER_358_2070 ();
 b15zdnd11an1n16x5 FILLER_358_2134 ();
 b15zdnd11an1n04x5 FILLER_358_2150 ();
 b15zdnd11an1n64x5 FILLER_358_2162 ();
 b15zdnd11an1n32x5 FILLER_358_2226 ();
 b15zdnd11an1n16x5 FILLER_358_2258 ();
 b15zdnd00an1n02x5 FILLER_358_2274 ();
 b15zdnd11an1n64x5 FILLER_359_0 ();
 b15zdnd11an1n64x5 FILLER_359_64 ();
 b15zdnd11an1n64x5 FILLER_359_128 ();
 b15zdnd11an1n64x5 FILLER_359_192 ();
 b15zdnd11an1n64x5 FILLER_359_256 ();
 b15zdnd11an1n64x5 FILLER_359_320 ();
 b15zdnd11an1n64x5 FILLER_359_384 ();
 b15zdnd11an1n64x5 FILLER_359_448 ();
 b15zdnd11an1n64x5 FILLER_359_512 ();
 b15zdnd11an1n64x5 FILLER_359_576 ();
 b15zdnd11an1n64x5 FILLER_359_640 ();
 b15zdnd11an1n64x5 FILLER_359_704 ();
 b15zdnd11an1n64x5 FILLER_359_768 ();
 b15zdnd11an1n64x5 FILLER_359_832 ();
 b15zdnd11an1n64x5 FILLER_359_896 ();
 b15zdnd11an1n64x5 FILLER_359_960 ();
 b15zdnd11an1n64x5 FILLER_359_1024 ();
 b15zdnd11an1n64x5 FILLER_359_1088 ();
 b15zdnd11an1n64x5 FILLER_359_1152 ();
 b15zdnd11an1n64x5 FILLER_359_1216 ();
 b15zdnd11an1n64x5 FILLER_359_1280 ();
 b15zdnd11an1n64x5 FILLER_359_1344 ();
 b15zdnd11an1n64x5 FILLER_359_1408 ();
 b15zdnd11an1n64x5 FILLER_359_1472 ();
 b15zdnd11an1n64x5 FILLER_359_1536 ();
 b15zdnd11an1n64x5 FILLER_359_1600 ();
 b15zdnd11an1n64x5 FILLER_359_1664 ();
 b15zdnd11an1n64x5 FILLER_359_1728 ();
 b15zdnd11an1n64x5 FILLER_359_1792 ();
 b15zdnd11an1n64x5 FILLER_359_1856 ();
 b15zdnd11an1n64x5 FILLER_359_1920 ();
 b15zdnd11an1n64x5 FILLER_359_1984 ();
 b15zdnd11an1n64x5 FILLER_359_2048 ();
 b15zdnd11an1n64x5 FILLER_359_2112 ();
 b15zdnd11an1n64x5 FILLER_359_2176 ();
 b15zdnd11an1n32x5 FILLER_359_2240 ();
 b15zdnd11an1n08x5 FILLER_359_2272 ();
 b15zdnd11an1n04x5 FILLER_359_2280 ();
 b15zdnd11an1n64x5 FILLER_360_8 ();
 b15zdnd11an1n64x5 FILLER_360_72 ();
 b15zdnd11an1n64x5 FILLER_360_136 ();
 b15zdnd11an1n64x5 FILLER_360_200 ();
 b15zdnd11an1n64x5 FILLER_360_264 ();
 b15zdnd11an1n64x5 FILLER_360_328 ();
 b15zdnd11an1n64x5 FILLER_360_392 ();
 b15zdnd11an1n64x5 FILLER_360_456 ();
 b15zdnd11an1n64x5 FILLER_360_520 ();
 b15zdnd11an1n64x5 FILLER_360_584 ();
 b15zdnd11an1n64x5 FILLER_360_648 ();
 b15zdnd11an1n04x5 FILLER_360_712 ();
 b15zdnd00an1n02x5 FILLER_360_716 ();
 b15zdnd11an1n64x5 FILLER_360_726 ();
 b15zdnd11an1n64x5 FILLER_360_790 ();
 b15zdnd11an1n64x5 FILLER_360_854 ();
 b15zdnd11an1n64x5 FILLER_360_918 ();
 b15zdnd11an1n64x5 FILLER_360_982 ();
 b15zdnd11an1n64x5 FILLER_360_1046 ();
 b15zdnd11an1n64x5 FILLER_360_1110 ();
 b15zdnd11an1n64x5 FILLER_360_1174 ();
 b15zdnd11an1n64x5 FILLER_360_1238 ();
 b15zdnd11an1n64x5 FILLER_360_1302 ();
 b15zdnd11an1n64x5 FILLER_360_1366 ();
 b15zdnd11an1n64x5 FILLER_360_1430 ();
 b15zdnd11an1n64x5 FILLER_360_1494 ();
 b15zdnd11an1n64x5 FILLER_360_1558 ();
 b15zdnd11an1n64x5 FILLER_360_1622 ();
 b15zdnd11an1n64x5 FILLER_360_1686 ();
 b15zdnd11an1n64x5 FILLER_360_1750 ();
 b15zdnd11an1n64x5 FILLER_360_1814 ();
 b15zdnd11an1n64x5 FILLER_360_1878 ();
 b15zdnd11an1n64x5 FILLER_360_1942 ();
 b15zdnd11an1n64x5 FILLER_360_2006 ();
 b15zdnd11an1n64x5 FILLER_360_2070 ();
 b15zdnd11an1n16x5 FILLER_360_2134 ();
 b15zdnd11an1n04x5 FILLER_360_2150 ();
 b15zdnd11an1n64x5 FILLER_360_2162 ();
 b15zdnd11an1n32x5 FILLER_360_2226 ();
 b15zdnd11an1n16x5 FILLER_360_2258 ();
 b15zdnd00an1n02x5 FILLER_360_2274 ();
 b15zdnd11an1n64x5 FILLER_361_0 ();
 b15zdnd11an1n64x5 FILLER_361_64 ();
 b15zdnd11an1n64x5 FILLER_361_128 ();
 b15zdnd11an1n64x5 FILLER_361_192 ();
 b15zdnd11an1n64x5 FILLER_361_256 ();
 b15zdnd11an1n64x5 FILLER_361_320 ();
 b15zdnd11an1n64x5 FILLER_361_384 ();
 b15zdnd11an1n64x5 FILLER_361_448 ();
 b15zdnd11an1n64x5 FILLER_361_512 ();
 b15zdnd11an1n64x5 FILLER_361_576 ();
 b15zdnd11an1n64x5 FILLER_361_640 ();
 b15zdnd11an1n64x5 FILLER_361_704 ();
 b15zdnd11an1n64x5 FILLER_361_768 ();
 b15zdnd11an1n64x5 FILLER_361_832 ();
 b15zdnd11an1n64x5 FILLER_361_896 ();
 b15zdnd11an1n64x5 FILLER_361_960 ();
 b15zdnd11an1n64x5 FILLER_361_1024 ();
 b15zdnd11an1n64x5 FILLER_361_1088 ();
 b15zdnd11an1n64x5 FILLER_361_1152 ();
 b15zdnd11an1n64x5 FILLER_361_1216 ();
 b15zdnd11an1n64x5 FILLER_361_1280 ();
 b15zdnd11an1n64x5 FILLER_361_1344 ();
 b15zdnd11an1n64x5 FILLER_361_1408 ();
 b15zdnd11an1n64x5 FILLER_361_1472 ();
 b15zdnd11an1n64x5 FILLER_361_1536 ();
 b15zdnd11an1n64x5 FILLER_361_1600 ();
 b15zdnd11an1n64x5 FILLER_361_1664 ();
 b15zdnd11an1n64x5 FILLER_361_1728 ();
 b15zdnd11an1n64x5 FILLER_361_1792 ();
 b15zdnd11an1n64x5 FILLER_361_1856 ();
 b15zdnd11an1n64x5 FILLER_361_1920 ();
 b15zdnd11an1n64x5 FILLER_361_1984 ();
 b15zdnd11an1n64x5 FILLER_361_2048 ();
 b15zdnd11an1n64x5 FILLER_361_2112 ();
 b15zdnd11an1n64x5 FILLER_361_2176 ();
 b15zdnd11an1n32x5 FILLER_361_2240 ();
 b15zdnd11an1n08x5 FILLER_361_2272 ();
 b15zdnd11an1n04x5 FILLER_361_2280 ();
 b15zdnd11an1n64x5 FILLER_362_8 ();
 b15zdnd11an1n64x5 FILLER_362_72 ();
 b15zdnd11an1n64x5 FILLER_362_136 ();
 b15zdnd11an1n64x5 FILLER_362_200 ();
 b15zdnd11an1n64x5 FILLER_362_264 ();
 b15zdnd11an1n64x5 FILLER_362_328 ();
 b15zdnd11an1n64x5 FILLER_362_392 ();
 b15zdnd11an1n64x5 FILLER_362_456 ();
 b15zdnd11an1n64x5 FILLER_362_520 ();
 b15zdnd11an1n64x5 FILLER_362_584 ();
 b15zdnd11an1n64x5 FILLER_362_648 ();
 b15zdnd11an1n04x5 FILLER_362_712 ();
 b15zdnd00an1n02x5 FILLER_362_716 ();
 b15zdnd11an1n64x5 FILLER_362_726 ();
 b15zdnd11an1n64x5 FILLER_362_790 ();
 b15zdnd11an1n64x5 FILLER_362_854 ();
 b15zdnd11an1n64x5 FILLER_362_918 ();
 b15zdnd11an1n64x5 FILLER_362_982 ();
 b15zdnd11an1n64x5 FILLER_362_1046 ();
 b15zdnd11an1n64x5 FILLER_362_1110 ();
 b15zdnd11an1n64x5 FILLER_362_1174 ();
 b15zdnd11an1n64x5 FILLER_362_1238 ();
 b15zdnd11an1n64x5 FILLER_362_1302 ();
 b15zdnd11an1n64x5 FILLER_362_1366 ();
 b15zdnd11an1n64x5 FILLER_362_1430 ();
 b15zdnd11an1n64x5 FILLER_362_1494 ();
 b15zdnd11an1n64x5 FILLER_362_1558 ();
 b15zdnd11an1n64x5 FILLER_362_1622 ();
 b15zdnd11an1n64x5 FILLER_362_1686 ();
 b15zdnd11an1n64x5 FILLER_362_1750 ();
 b15zdnd11an1n64x5 FILLER_362_1814 ();
 b15zdnd11an1n64x5 FILLER_362_1878 ();
 b15zdnd11an1n64x5 FILLER_362_1942 ();
 b15zdnd11an1n64x5 FILLER_362_2006 ();
 b15zdnd11an1n64x5 FILLER_362_2070 ();
 b15zdnd11an1n16x5 FILLER_362_2134 ();
 b15zdnd11an1n04x5 FILLER_362_2150 ();
 b15zdnd11an1n64x5 FILLER_362_2162 ();
 b15zdnd11an1n32x5 FILLER_362_2226 ();
 b15zdnd11an1n16x5 FILLER_362_2258 ();
 b15zdnd00an1n02x5 FILLER_362_2274 ();
 b15zdnd11an1n64x5 FILLER_363_0 ();
 b15zdnd11an1n64x5 FILLER_363_64 ();
 b15zdnd11an1n64x5 FILLER_363_128 ();
 b15zdnd11an1n64x5 FILLER_363_192 ();
 b15zdnd11an1n64x5 FILLER_363_256 ();
 b15zdnd11an1n64x5 FILLER_363_320 ();
 b15zdnd11an1n64x5 FILLER_363_384 ();
 b15zdnd11an1n64x5 FILLER_363_448 ();
 b15zdnd11an1n64x5 FILLER_363_512 ();
 b15zdnd11an1n64x5 FILLER_363_576 ();
 b15zdnd11an1n64x5 FILLER_363_640 ();
 b15zdnd11an1n64x5 FILLER_363_704 ();
 b15zdnd11an1n64x5 FILLER_363_768 ();
 b15zdnd11an1n64x5 FILLER_363_832 ();
 b15zdnd11an1n64x5 FILLER_363_896 ();
 b15zdnd11an1n64x5 FILLER_363_960 ();
 b15zdnd11an1n64x5 FILLER_363_1024 ();
 b15zdnd11an1n64x5 FILLER_363_1088 ();
 b15zdnd11an1n64x5 FILLER_363_1152 ();
 b15zdnd11an1n64x5 FILLER_363_1216 ();
 b15zdnd11an1n64x5 FILLER_363_1280 ();
 b15zdnd11an1n64x5 FILLER_363_1344 ();
 b15zdnd11an1n64x5 FILLER_363_1408 ();
 b15zdnd11an1n64x5 FILLER_363_1472 ();
 b15zdnd11an1n64x5 FILLER_363_1536 ();
 b15zdnd11an1n64x5 FILLER_363_1600 ();
 b15zdnd11an1n64x5 FILLER_363_1664 ();
 b15zdnd11an1n64x5 FILLER_363_1728 ();
 b15zdnd11an1n64x5 FILLER_363_1792 ();
 b15zdnd11an1n64x5 FILLER_363_1856 ();
 b15zdnd11an1n64x5 FILLER_363_1920 ();
 b15zdnd11an1n64x5 FILLER_363_1984 ();
 b15zdnd11an1n64x5 FILLER_363_2048 ();
 b15zdnd11an1n64x5 FILLER_363_2112 ();
 b15zdnd11an1n64x5 FILLER_363_2176 ();
 b15zdnd11an1n32x5 FILLER_363_2240 ();
 b15zdnd11an1n08x5 FILLER_363_2272 ();
 b15zdnd11an1n04x5 FILLER_363_2280 ();
 b15zdnd11an1n64x5 FILLER_364_8 ();
 b15zdnd11an1n64x5 FILLER_364_72 ();
 b15zdnd11an1n64x5 FILLER_364_136 ();
 b15zdnd11an1n64x5 FILLER_364_200 ();
 b15zdnd11an1n64x5 FILLER_364_264 ();
 b15zdnd11an1n64x5 FILLER_364_328 ();
 b15zdnd11an1n64x5 FILLER_364_392 ();
 b15zdnd11an1n64x5 FILLER_364_456 ();
 b15zdnd11an1n64x5 FILLER_364_520 ();
 b15zdnd11an1n64x5 FILLER_364_584 ();
 b15zdnd11an1n64x5 FILLER_364_648 ();
 b15zdnd11an1n04x5 FILLER_364_712 ();
 b15zdnd00an1n02x5 FILLER_364_716 ();
 b15zdnd11an1n64x5 FILLER_364_726 ();
 b15zdnd11an1n64x5 FILLER_364_790 ();
 b15zdnd11an1n64x5 FILLER_364_854 ();
 b15zdnd11an1n64x5 FILLER_364_918 ();
 b15zdnd11an1n64x5 FILLER_364_982 ();
 b15zdnd11an1n64x5 FILLER_364_1046 ();
 b15zdnd11an1n64x5 FILLER_364_1110 ();
 b15zdnd11an1n64x5 FILLER_364_1174 ();
 b15zdnd11an1n64x5 FILLER_364_1238 ();
 b15zdnd11an1n64x5 FILLER_364_1302 ();
 b15zdnd11an1n64x5 FILLER_364_1366 ();
 b15zdnd11an1n64x5 FILLER_364_1430 ();
 b15zdnd11an1n64x5 FILLER_364_1494 ();
 b15zdnd11an1n64x5 FILLER_364_1558 ();
 b15zdnd11an1n64x5 FILLER_364_1622 ();
 b15zdnd11an1n64x5 FILLER_364_1686 ();
 b15zdnd11an1n64x5 FILLER_364_1750 ();
 b15zdnd11an1n64x5 FILLER_364_1814 ();
 b15zdnd11an1n64x5 FILLER_364_1878 ();
 b15zdnd11an1n64x5 FILLER_364_1942 ();
 b15zdnd11an1n64x5 FILLER_364_2006 ();
 b15zdnd11an1n64x5 FILLER_364_2070 ();
 b15zdnd11an1n16x5 FILLER_364_2134 ();
 b15zdnd11an1n04x5 FILLER_364_2150 ();
 b15zdnd11an1n64x5 FILLER_364_2162 ();
 b15zdnd11an1n32x5 FILLER_364_2226 ();
 b15zdnd11an1n16x5 FILLER_364_2258 ();
 b15zdnd00an1n02x5 FILLER_364_2274 ();
 b15zdnd11an1n64x5 FILLER_365_0 ();
 b15zdnd11an1n64x5 FILLER_365_64 ();
 b15zdnd11an1n64x5 FILLER_365_128 ();
 b15zdnd11an1n64x5 FILLER_365_192 ();
 b15zdnd11an1n64x5 FILLER_365_256 ();
 b15zdnd11an1n64x5 FILLER_365_320 ();
 b15zdnd11an1n64x5 FILLER_365_384 ();
 b15zdnd11an1n64x5 FILLER_365_448 ();
 b15zdnd11an1n64x5 FILLER_365_512 ();
 b15zdnd11an1n64x5 FILLER_365_576 ();
 b15zdnd11an1n64x5 FILLER_365_640 ();
 b15zdnd11an1n64x5 FILLER_365_704 ();
 b15zdnd11an1n64x5 FILLER_365_768 ();
 b15zdnd11an1n64x5 FILLER_365_832 ();
 b15zdnd11an1n64x5 FILLER_365_896 ();
 b15zdnd11an1n64x5 FILLER_365_960 ();
 b15zdnd11an1n64x5 FILLER_365_1024 ();
 b15zdnd11an1n64x5 FILLER_365_1088 ();
 b15zdnd11an1n64x5 FILLER_365_1152 ();
 b15zdnd11an1n64x5 FILLER_365_1216 ();
 b15zdnd11an1n64x5 FILLER_365_1280 ();
 b15zdnd11an1n64x5 FILLER_365_1344 ();
 b15zdnd11an1n64x5 FILLER_365_1408 ();
 b15zdnd11an1n64x5 FILLER_365_1472 ();
 b15zdnd11an1n64x5 FILLER_365_1536 ();
 b15zdnd11an1n64x5 FILLER_365_1600 ();
 b15zdnd11an1n64x5 FILLER_365_1664 ();
 b15zdnd11an1n64x5 FILLER_365_1728 ();
 b15zdnd11an1n64x5 FILLER_365_1792 ();
 b15zdnd11an1n64x5 FILLER_365_1856 ();
 b15zdnd11an1n64x5 FILLER_365_1920 ();
 b15zdnd11an1n64x5 FILLER_365_1984 ();
 b15zdnd11an1n64x5 FILLER_365_2048 ();
 b15zdnd11an1n64x5 FILLER_365_2112 ();
 b15zdnd11an1n64x5 FILLER_365_2176 ();
 b15zdnd11an1n32x5 FILLER_365_2240 ();
 b15zdnd11an1n08x5 FILLER_365_2272 ();
 b15zdnd11an1n04x5 FILLER_365_2280 ();
 b15zdnd11an1n64x5 FILLER_366_8 ();
 b15zdnd11an1n64x5 FILLER_366_72 ();
 b15zdnd11an1n64x5 FILLER_366_136 ();
 b15zdnd11an1n64x5 FILLER_366_200 ();
 b15zdnd11an1n64x5 FILLER_366_264 ();
 b15zdnd11an1n64x5 FILLER_366_328 ();
 b15zdnd11an1n64x5 FILLER_366_392 ();
 b15zdnd11an1n64x5 FILLER_366_456 ();
 b15zdnd11an1n64x5 FILLER_366_520 ();
 b15zdnd11an1n64x5 FILLER_366_584 ();
 b15zdnd11an1n64x5 FILLER_366_648 ();
 b15zdnd11an1n04x5 FILLER_366_712 ();
 b15zdnd00an1n02x5 FILLER_366_716 ();
 b15zdnd11an1n64x5 FILLER_366_726 ();
 b15zdnd11an1n64x5 FILLER_366_790 ();
 b15zdnd11an1n64x5 FILLER_366_854 ();
 b15zdnd11an1n64x5 FILLER_366_918 ();
 b15zdnd11an1n64x5 FILLER_366_982 ();
 b15zdnd11an1n64x5 FILLER_366_1046 ();
 b15zdnd11an1n64x5 FILLER_366_1110 ();
 b15zdnd11an1n64x5 FILLER_366_1174 ();
 b15zdnd11an1n64x5 FILLER_366_1238 ();
 b15zdnd11an1n64x5 FILLER_366_1302 ();
 b15zdnd11an1n64x5 FILLER_366_1366 ();
 b15zdnd11an1n64x5 FILLER_366_1430 ();
 b15zdnd11an1n64x5 FILLER_366_1494 ();
 b15zdnd11an1n64x5 FILLER_366_1558 ();
 b15zdnd11an1n64x5 FILLER_366_1622 ();
 b15zdnd11an1n64x5 FILLER_366_1686 ();
 b15zdnd11an1n64x5 FILLER_366_1750 ();
 b15zdnd11an1n64x5 FILLER_366_1814 ();
 b15zdnd11an1n64x5 FILLER_366_1878 ();
 b15zdnd11an1n64x5 FILLER_366_1942 ();
 b15zdnd11an1n64x5 FILLER_366_2006 ();
 b15zdnd11an1n64x5 FILLER_366_2070 ();
 b15zdnd11an1n16x5 FILLER_366_2134 ();
 b15zdnd11an1n04x5 FILLER_366_2150 ();
 b15zdnd11an1n64x5 FILLER_366_2162 ();
 b15zdnd11an1n32x5 FILLER_366_2226 ();
 b15zdnd11an1n16x5 FILLER_366_2258 ();
 b15zdnd00an1n02x5 FILLER_366_2274 ();
 b15zdnd11an1n64x5 FILLER_367_0 ();
 b15zdnd11an1n64x5 FILLER_367_64 ();
 b15zdnd11an1n64x5 FILLER_367_128 ();
 b15zdnd11an1n64x5 FILLER_367_192 ();
 b15zdnd11an1n64x5 FILLER_367_256 ();
 b15zdnd11an1n64x5 FILLER_367_320 ();
 b15zdnd11an1n64x5 FILLER_367_384 ();
 b15zdnd11an1n64x5 FILLER_367_448 ();
 b15zdnd11an1n64x5 FILLER_367_512 ();
 b15zdnd11an1n64x5 FILLER_367_576 ();
 b15zdnd11an1n64x5 FILLER_367_640 ();
 b15zdnd11an1n64x5 FILLER_367_704 ();
 b15zdnd11an1n64x5 FILLER_367_768 ();
 b15zdnd11an1n64x5 FILLER_367_832 ();
 b15zdnd11an1n64x5 FILLER_367_896 ();
 b15zdnd11an1n64x5 FILLER_367_960 ();
 b15zdnd11an1n64x5 FILLER_367_1024 ();
 b15zdnd11an1n64x5 FILLER_367_1088 ();
 b15zdnd11an1n64x5 FILLER_367_1152 ();
 b15zdnd11an1n64x5 FILLER_367_1216 ();
 b15zdnd11an1n64x5 FILLER_367_1280 ();
 b15zdnd11an1n64x5 FILLER_367_1344 ();
 b15zdnd11an1n64x5 FILLER_367_1408 ();
 b15zdnd11an1n64x5 FILLER_367_1472 ();
 b15zdnd11an1n64x5 FILLER_367_1536 ();
 b15zdnd11an1n64x5 FILLER_367_1600 ();
 b15zdnd11an1n64x5 FILLER_367_1664 ();
 b15zdnd11an1n64x5 FILLER_367_1728 ();
 b15zdnd11an1n64x5 FILLER_367_1792 ();
 b15zdnd11an1n64x5 FILLER_367_1856 ();
 b15zdnd11an1n64x5 FILLER_367_1920 ();
 b15zdnd11an1n64x5 FILLER_367_1984 ();
 b15zdnd11an1n64x5 FILLER_367_2048 ();
 b15zdnd11an1n64x5 FILLER_367_2112 ();
 b15zdnd11an1n64x5 FILLER_367_2176 ();
 b15zdnd11an1n32x5 FILLER_367_2240 ();
 b15zdnd11an1n08x5 FILLER_367_2272 ();
 b15zdnd11an1n04x5 FILLER_367_2280 ();
 b15zdnd11an1n64x5 FILLER_368_8 ();
 b15zdnd11an1n64x5 FILLER_368_72 ();
 b15zdnd11an1n64x5 FILLER_368_136 ();
 b15zdnd11an1n64x5 FILLER_368_200 ();
 b15zdnd11an1n64x5 FILLER_368_264 ();
 b15zdnd11an1n64x5 FILLER_368_328 ();
 b15zdnd11an1n64x5 FILLER_368_392 ();
 b15zdnd11an1n64x5 FILLER_368_456 ();
 b15zdnd11an1n64x5 FILLER_368_520 ();
 b15zdnd11an1n64x5 FILLER_368_584 ();
 b15zdnd11an1n64x5 FILLER_368_648 ();
 b15zdnd11an1n04x5 FILLER_368_712 ();
 b15zdnd00an1n02x5 FILLER_368_716 ();
 b15zdnd11an1n64x5 FILLER_368_726 ();
 b15zdnd11an1n64x5 FILLER_368_790 ();
 b15zdnd11an1n64x5 FILLER_368_854 ();
 b15zdnd11an1n64x5 FILLER_368_918 ();
 b15zdnd11an1n64x5 FILLER_368_982 ();
 b15zdnd11an1n64x5 FILLER_368_1046 ();
 b15zdnd11an1n64x5 FILLER_368_1110 ();
 b15zdnd11an1n64x5 FILLER_368_1174 ();
 b15zdnd11an1n64x5 FILLER_368_1238 ();
 b15zdnd11an1n64x5 FILLER_368_1302 ();
 b15zdnd11an1n64x5 FILLER_368_1366 ();
 b15zdnd11an1n64x5 FILLER_368_1430 ();
 b15zdnd11an1n64x5 FILLER_368_1494 ();
 b15zdnd11an1n64x5 FILLER_368_1558 ();
 b15zdnd11an1n64x5 FILLER_368_1622 ();
 b15zdnd11an1n64x5 FILLER_368_1686 ();
 b15zdnd11an1n64x5 FILLER_368_1750 ();
 b15zdnd11an1n64x5 FILLER_368_1814 ();
 b15zdnd11an1n64x5 FILLER_368_1878 ();
 b15zdnd11an1n64x5 FILLER_368_1942 ();
 b15zdnd11an1n64x5 FILLER_368_2006 ();
 b15zdnd11an1n64x5 FILLER_368_2070 ();
 b15zdnd11an1n16x5 FILLER_368_2134 ();
 b15zdnd11an1n04x5 FILLER_368_2150 ();
 b15zdnd11an1n64x5 FILLER_368_2162 ();
 b15zdnd11an1n32x5 FILLER_368_2226 ();
 b15zdnd11an1n16x5 FILLER_368_2258 ();
 b15zdnd00an1n02x5 FILLER_368_2274 ();
 b15zdnd11an1n64x5 FILLER_369_0 ();
 b15zdnd11an1n64x5 FILLER_369_64 ();
 b15zdnd11an1n64x5 FILLER_369_128 ();
 b15zdnd11an1n64x5 FILLER_369_192 ();
 b15zdnd11an1n64x5 FILLER_369_256 ();
 b15zdnd11an1n64x5 FILLER_369_320 ();
 b15zdnd11an1n64x5 FILLER_369_384 ();
 b15zdnd11an1n64x5 FILLER_369_448 ();
 b15zdnd11an1n64x5 FILLER_369_512 ();
 b15zdnd11an1n64x5 FILLER_369_576 ();
 b15zdnd11an1n64x5 FILLER_369_640 ();
 b15zdnd11an1n64x5 FILLER_369_704 ();
 b15zdnd11an1n64x5 FILLER_369_768 ();
 b15zdnd11an1n64x5 FILLER_369_832 ();
 b15zdnd11an1n64x5 FILLER_369_896 ();
 b15zdnd11an1n64x5 FILLER_369_960 ();
 b15zdnd11an1n64x5 FILLER_369_1024 ();
 b15zdnd11an1n64x5 FILLER_369_1088 ();
 b15zdnd11an1n64x5 FILLER_369_1152 ();
 b15zdnd11an1n64x5 FILLER_369_1216 ();
 b15zdnd11an1n64x5 FILLER_369_1280 ();
 b15zdnd11an1n64x5 FILLER_369_1344 ();
 b15zdnd11an1n64x5 FILLER_369_1408 ();
 b15zdnd11an1n64x5 FILLER_369_1472 ();
 b15zdnd11an1n64x5 FILLER_369_1536 ();
 b15zdnd11an1n64x5 FILLER_369_1600 ();
 b15zdnd11an1n64x5 FILLER_369_1664 ();
 b15zdnd11an1n64x5 FILLER_369_1728 ();
 b15zdnd11an1n64x5 FILLER_369_1792 ();
 b15zdnd11an1n64x5 FILLER_369_1856 ();
 b15zdnd11an1n64x5 FILLER_369_1920 ();
 b15zdnd11an1n64x5 FILLER_369_1984 ();
 b15zdnd11an1n64x5 FILLER_369_2048 ();
 b15zdnd11an1n64x5 FILLER_369_2112 ();
 b15zdnd11an1n64x5 FILLER_369_2176 ();
 b15zdnd11an1n32x5 FILLER_369_2240 ();
 b15zdnd11an1n08x5 FILLER_369_2272 ();
 b15zdnd11an1n04x5 FILLER_369_2280 ();
 b15zdnd11an1n64x5 FILLER_370_8 ();
 b15zdnd11an1n64x5 FILLER_370_72 ();
 b15zdnd11an1n64x5 FILLER_370_136 ();
 b15zdnd11an1n64x5 FILLER_370_200 ();
 b15zdnd11an1n64x5 FILLER_370_264 ();
 b15zdnd11an1n64x5 FILLER_370_328 ();
 b15zdnd11an1n64x5 FILLER_370_392 ();
 b15zdnd11an1n64x5 FILLER_370_456 ();
 b15zdnd11an1n64x5 FILLER_370_520 ();
 b15zdnd11an1n64x5 FILLER_370_584 ();
 b15zdnd11an1n64x5 FILLER_370_648 ();
 b15zdnd11an1n04x5 FILLER_370_712 ();
 b15zdnd00an1n02x5 FILLER_370_716 ();
 b15zdnd11an1n64x5 FILLER_370_726 ();
 b15zdnd11an1n64x5 FILLER_370_790 ();
 b15zdnd11an1n64x5 FILLER_370_854 ();
 b15zdnd11an1n64x5 FILLER_370_918 ();
 b15zdnd11an1n64x5 FILLER_370_982 ();
 b15zdnd11an1n64x5 FILLER_370_1046 ();
 b15zdnd11an1n64x5 FILLER_370_1110 ();
 b15zdnd11an1n64x5 FILLER_370_1174 ();
 b15zdnd11an1n64x5 FILLER_370_1238 ();
 b15zdnd11an1n64x5 FILLER_370_1302 ();
 b15zdnd11an1n64x5 FILLER_370_1366 ();
 b15zdnd11an1n64x5 FILLER_370_1430 ();
 b15zdnd11an1n64x5 FILLER_370_1494 ();
 b15zdnd11an1n64x5 FILLER_370_1558 ();
 b15zdnd11an1n64x5 FILLER_370_1622 ();
 b15zdnd11an1n64x5 FILLER_370_1686 ();
 b15zdnd11an1n64x5 FILLER_370_1750 ();
 b15zdnd11an1n64x5 FILLER_370_1814 ();
 b15zdnd11an1n64x5 FILLER_370_1878 ();
 b15zdnd11an1n64x5 FILLER_370_1942 ();
 b15zdnd11an1n64x5 FILLER_370_2006 ();
 b15zdnd11an1n64x5 FILLER_370_2070 ();
 b15zdnd11an1n16x5 FILLER_370_2134 ();
 b15zdnd11an1n04x5 FILLER_370_2150 ();
 b15zdnd11an1n64x5 FILLER_370_2162 ();
 b15zdnd11an1n32x5 FILLER_370_2226 ();
 b15zdnd11an1n16x5 FILLER_370_2258 ();
 b15zdnd00an1n02x5 FILLER_370_2274 ();
 b15zdnd11an1n64x5 FILLER_371_0 ();
 b15zdnd11an1n64x5 FILLER_371_64 ();
 b15zdnd11an1n64x5 FILLER_371_128 ();
 b15zdnd11an1n64x5 FILLER_371_192 ();
 b15zdnd11an1n64x5 FILLER_371_256 ();
 b15zdnd11an1n64x5 FILLER_371_320 ();
 b15zdnd11an1n64x5 FILLER_371_384 ();
 b15zdnd11an1n64x5 FILLER_371_448 ();
 b15zdnd11an1n64x5 FILLER_371_512 ();
 b15zdnd11an1n64x5 FILLER_371_576 ();
 b15zdnd11an1n64x5 FILLER_371_640 ();
 b15zdnd11an1n64x5 FILLER_371_704 ();
 b15zdnd11an1n64x5 FILLER_371_768 ();
 b15zdnd11an1n64x5 FILLER_371_832 ();
 b15zdnd11an1n64x5 FILLER_371_896 ();
 b15zdnd11an1n64x5 FILLER_371_960 ();
 b15zdnd11an1n64x5 FILLER_371_1024 ();
 b15zdnd11an1n64x5 FILLER_371_1088 ();
 b15zdnd11an1n64x5 FILLER_371_1152 ();
 b15zdnd11an1n64x5 FILLER_371_1216 ();
 b15zdnd11an1n64x5 FILLER_371_1280 ();
 b15zdnd11an1n64x5 FILLER_371_1344 ();
 b15zdnd11an1n64x5 FILLER_371_1408 ();
 b15zdnd11an1n64x5 FILLER_371_1472 ();
 b15zdnd11an1n64x5 FILLER_371_1536 ();
 b15zdnd11an1n64x5 FILLER_371_1600 ();
 b15zdnd11an1n64x5 FILLER_371_1664 ();
 b15zdnd11an1n64x5 FILLER_371_1728 ();
 b15zdnd11an1n64x5 FILLER_371_1792 ();
 b15zdnd11an1n64x5 FILLER_371_1856 ();
 b15zdnd11an1n64x5 FILLER_371_1920 ();
 b15zdnd11an1n64x5 FILLER_371_1984 ();
 b15zdnd11an1n64x5 FILLER_371_2048 ();
 b15zdnd11an1n64x5 FILLER_371_2112 ();
 b15zdnd11an1n64x5 FILLER_371_2176 ();
 b15zdnd11an1n32x5 FILLER_371_2240 ();
 b15zdnd11an1n08x5 FILLER_371_2272 ();
 b15zdnd11an1n04x5 FILLER_371_2280 ();
 b15zdnd11an1n64x5 FILLER_372_8 ();
 b15zdnd11an1n64x5 FILLER_372_72 ();
 b15zdnd11an1n64x5 FILLER_372_136 ();
 b15zdnd11an1n64x5 FILLER_372_200 ();
 b15zdnd11an1n64x5 FILLER_372_264 ();
 b15zdnd11an1n64x5 FILLER_372_328 ();
 b15zdnd11an1n64x5 FILLER_372_392 ();
 b15zdnd11an1n64x5 FILLER_372_456 ();
 b15zdnd11an1n64x5 FILLER_372_520 ();
 b15zdnd11an1n64x5 FILLER_372_584 ();
 b15zdnd11an1n64x5 FILLER_372_648 ();
 b15zdnd11an1n04x5 FILLER_372_712 ();
 b15zdnd00an1n02x5 FILLER_372_716 ();
 b15zdnd11an1n64x5 FILLER_372_726 ();
 b15zdnd11an1n64x5 FILLER_372_790 ();
 b15zdnd11an1n64x5 FILLER_372_854 ();
 b15zdnd11an1n64x5 FILLER_372_918 ();
 b15zdnd11an1n64x5 FILLER_372_982 ();
 b15zdnd11an1n64x5 FILLER_372_1046 ();
 b15zdnd11an1n64x5 FILLER_372_1110 ();
 b15zdnd11an1n64x5 FILLER_372_1174 ();
 b15zdnd11an1n64x5 FILLER_372_1238 ();
 b15zdnd11an1n64x5 FILLER_372_1302 ();
 b15zdnd11an1n64x5 FILLER_372_1366 ();
 b15zdnd11an1n64x5 FILLER_372_1430 ();
 b15zdnd11an1n64x5 FILLER_372_1494 ();
 b15zdnd11an1n64x5 FILLER_372_1558 ();
 b15zdnd11an1n64x5 FILLER_372_1622 ();
 b15zdnd11an1n64x5 FILLER_372_1686 ();
 b15zdnd11an1n64x5 FILLER_372_1750 ();
 b15zdnd11an1n64x5 FILLER_372_1814 ();
 b15zdnd11an1n64x5 FILLER_372_1878 ();
 b15zdnd11an1n64x5 FILLER_372_1942 ();
 b15zdnd11an1n64x5 FILLER_372_2006 ();
 b15zdnd11an1n64x5 FILLER_372_2070 ();
 b15zdnd11an1n16x5 FILLER_372_2134 ();
 b15zdnd11an1n04x5 FILLER_372_2150 ();
 b15zdnd11an1n64x5 FILLER_372_2162 ();
 b15zdnd11an1n32x5 FILLER_372_2226 ();
 b15zdnd11an1n16x5 FILLER_372_2258 ();
 b15zdnd00an1n02x5 FILLER_372_2274 ();
 b15zdnd11an1n64x5 FILLER_373_0 ();
 b15zdnd11an1n64x5 FILLER_373_64 ();
 b15zdnd11an1n64x5 FILLER_373_128 ();
 b15zdnd11an1n64x5 FILLER_373_192 ();
 b15zdnd11an1n64x5 FILLER_373_256 ();
 b15zdnd11an1n64x5 FILLER_373_320 ();
 b15zdnd11an1n64x5 FILLER_373_384 ();
 b15zdnd11an1n64x5 FILLER_373_448 ();
 b15zdnd11an1n64x5 FILLER_373_512 ();
 b15zdnd11an1n64x5 FILLER_373_576 ();
 b15zdnd11an1n64x5 FILLER_373_640 ();
 b15zdnd11an1n64x5 FILLER_373_704 ();
 b15zdnd11an1n64x5 FILLER_373_768 ();
 b15zdnd11an1n64x5 FILLER_373_832 ();
 b15zdnd11an1n64x5 FILLER_373_896 ();
 b15zdnd11an1n64x5 FILLER_373_960 ();
 b15zdnd11an1n64x5 FILLER_373_1024 ();
 b15zdnd11an1n64x5 FILLER_373_1088 ();
 b15zdnd11an1n64x5 FILLER_373_1152 ();
 b15zdnd11an1n64x5 FILLER_373_1216 ();
 b15zdnd11an1n64x5 FILLER_373_1280 ();
 b15zdnd11an1n64x5 FILLER_373_1344 ();
 b15zdnd11an1n64x5 FILLER_373_1408 ();
 b15zdnd11an1n64x5 FILLER_373_1472 ();
 b15zdnd11an1n64x5 FILLER_373_1536 ();
 b15zdnd11an1n64x5 FILLER_373_1600 ();
 b15zdnd11an1n64x5 FILLER_373_1664 ();
 b15zdnd11an1n64x5 FILLER_373_1728 ();
 b15zdnd11an1n64x5 FILLER_373_1792 ();
 b15zdnd11an1n64x5 FILLER_373_1856 ();
 b15zdnd11an1n64x5 FILLER_373_1920 ();
 b15zdnd11an1n64x5 FILLER_373_1984 ();
 b15zdnd11an1n64x5 FILLER_373_2048 ();
 b15zdnd11an1n64x5 FILLER_373_2112 ();
 b15zdnd11an1n64x5 FILLER_373_2176 ();
 b15zdnd11an1n32x5 FILLER_373_2240 ();
 b15zdnd11an1n08x5 FILLER_373_2272 ();
 b15zdnd11an1n04x5 FILLER_373_2280 ();
 b15zdnd11an1n64x5 FILLER_374_8 ();
 b15zdnd11an1n64x5 FILLER_374_72 ();
 b15zdnd11an1n64x5 FILLER_374_136 ();
 b15zdnd11an1n64x5 FILLER_374_200 ();
 b15zdnd11an1n64x5 FILLER_374_264 ();
 b15zdnd11an1n64x5 FILLER_374_328 ();
 b15zdnd11an1n64x5 FILLER_374_392 ();
 b15zdnd11an1n64x5 FILLER_374_456 ();
 b15zdnd11an1n64x5 FILLER_374_520 ();
 b15zdnd11an1n64x5 FILLER_374_584 ();
 b15zdnd11an1n64x5 FILLER_374_648 ();
 b15zdnd11an1n04x5 FILLER_374_712 ();
 b15zdnd00an1n02x5 FILLER_374_716 ();
 b15zdnd11an1n64x5 FILLER_374_726 ();
 b15zdnd11an1n64x5 FILLER_374_790 ();
 b15zdnd11an1n64x5 FILLER_374_854 ();
 b15zdnd11an1n64x5 FILLER_374_918 ();
 b15zdnd11an1n64x5 FILLER_374_982 ();
 b15zdnd11an1n64x5 FILLER_374_1046 ();
 b15zdnd11an1n64x5 FILLER_374_1110 ();
 b15zdnd11an1n64x5 FILLER_374_1174 ();
 b15zdnd11an1n64x5 FILLER_374_1238 ();
 b15zdnd11an1n64x5 FILLER_374_1302 ();
 b15zdnd11an1n64x5 FILLER_374_1366 ();
 b15zdnd11an1n64x5 FILLER_374_1430 ();
 b15zdnd11an1n64x5 FILLER_374_1494 ();
 b15zdnd11an1n64x5 FILLER_374_1558 ();
 b15zdnd11an1n64x5 FILLER_374_1622 ();
 b15zdnd11an1n64x5 FILLER_374_1686 ();
 b15zdnd11an1n64x5 FILLER_374_1750 ();
 b15zdnd11an1n64x5 FILLER_374_1814 ();
 b15zdnd11an1n64x5 FILLER_374_1878 ();
 b15zdnd11an1n64x5 FILLER_374_1942 ();
 b15zdnd11an1n64x5 FILLER_374_2006 ();
 b15zdnd11an1n64x5 FILLER_374_2070 ();
 b15zdnd11an1n16x5 FILLER_374_2134 ();
 b15zdnd11an1n04x5 FILLER_374_2150 ();
 b15zdnd11an1n64x5 FILLER_374_2162 ();
 b15zdnd11an1n32x5 FILLER_374_2226 ();
 b15zdnd11an1n16x5 FILLER_374_2258 ();
 b15zdnd00an1n02x5 FILLER_374_2274 ();
 b15zdnd11an1n64x5 FILLER_375_0 ();
 b15zdnd11an1n64x5 FILLER_375_64 ();
 b15zdnd11an1n64x5 FILLER_375_128 ();
 b15zdnd11an1n64x5 FILLER_375_192 ();
 b15zdnd11an1n64x5 FILLER_375_256 ();
 b15zdnd11an1n64x5 FILLER_375_320 ();
 b15zdnd11an1n64x5 FILLER_375_384 ();
 b15zdnd11an1n64x5 FILLER_375_448 ();
 b15zdnd11an1n64x5 FILLER_375_512 ();
 b15zdnd11an1n64x5 FILLER_375_576 ();
 b15zdnd11an1n64x5 FILLER_375_640 ();
 b15zdnd11an1n64x5 FILLER_375_704 ();
 b15zdnd11an1n64x5 FILLER_375_768 ();
 b15zdnd11an1n64x5 FILLER_375_832 ();
 b15zdnd11an1n64x5 FILLER_375_896 ();
 b15zdnd11an1n64x5 FILLER_375_960 ();
 b15zdnd11an1n64x5 FILLER_375_1024 ();
 b15zdnd11an1n64x5 FILLER_375_1088 ();
 b15zdnd11an1n64x5 FILLER_375_1152 ();
 b15zdnd11an1n64x5 FILLER_375_1216 ();
 b15zdnd11an1n64x5 FILLER_375_1280 ();
 b15zdnd11an1n64x5 FILLER_375_1344 ();
 b15zdnd11an1n64x5 FILLER_375_1408 ();
 b15zdnd11an1n64x5 FILLER_375_1472 ();
 b15zdnd11an1n64x5 FILLER_375_1536 ();
 b15zdnd11an1n64x5 FILLER_375_1600 ();
 b15zdnd11an1n64x5 FILLER_375_1664 ();
 b15zdnd11an1n64x5 FILLER_375_1728 ();
 b15zdnd11an1n64x5 FILLER_375_1792 ();
 b15zdnd11an1n64x5 FILLER_375_1856 ();
 b15zdnd11an1n64x5 FILLER_375_1920 ();
 b15zdnd11an1n64x5 FILLER_375_1984 ();
 b15zdnd11an1n64x5 FILLER_375_2048 ();
 b15zdnd11an1n64x5 FILLER_375_2112 ();
 b15zdnd11an1n64x5 FILLER_375_2176 ();
 b15zdnd11an1n32x5 FILLER_375_2240 ();
 b15zdnd11an1n08x5 FILLER_375_2272 ();
 b15zdnd11an1n04x5 FILLER_375_2280 ();
 b15zdnd11an1n64x5 FILLER_376_8 ();
 b15zdnd11an1n64x5 FILLER_376_72 ();
 b15zdnd11an1n64x5 FILLER_376_136 ();
 b15zdnd11an1n64x5 FILLER_376_200 ();
 b15zdnd11an1n64x5 FILLER_376_264 ();
 b15zdnd11an1n64x5 FILLER_376_328 ();
 b15zdnd11an1n64x5 FILLER_376_392 ();
 b15zdnd11an1n64x5 FILLER_376_456 ();
 b15zdnd11an1n64x5 FILLER_376_520 ();
 b15zdnd11an1n64x5 FILLER_376_584 ();
 b15zdnd11an1n64x5 FILLER_376_648 ();
 b15zdnd11an1n04x5 FILLER_376_712 ();
 b15zdnd00an1n02x5 FILLER_376_716 ();
 b15zdnd11an1n64x5 FILLER_376_726 ();
 b15zdnd11an1n64x5 FILLER_376_790 ();
 b15zdnd11an1n64x5 FILLER_376_854 ();
 b15zdnd11an1n64x5 FILLER_376_918 ();
 b15zdnd11an1n64x5 FILLER_376_982 ();
 b15zdnd11an1n64x5 FILLER_376_1046 ();
 b15zdnd11an1n64x5 FILLER_376_1110 ();
 b15zdnd11an1n64x5 FILLER_376_1174 ();
 b15zdnd11an1n64x5 FILLER_376_1238 ();
 b15zdnd11an1n64x5 FILLER_376_1302 ();
 b15zdnd11an1n64x5 FILLER_376_1366 ();
 b15zdnd11an1n64x5 FILLER_376_1430 ();
 b15zdnd11an1n64x5 FILLER_376_1494 ();
 b15zdnd11an1n64x5 FILLER_376_1558 ();
 b15zdnd11an1n64x5 FILLER_376_1622 ();
 b15zdnd11an1n64x5 FILLER_376_1686 ();
 b15zdnd11an1n64x5 FILLER_376_1750 ();
 b15zdnd11an1n64x5 FILLER_376_1814 ();
 b15zdnd11an1n64x5 FILLER_376_1878 ();
 b15zdnd11an1n64x5 FILLER_376_1942 ();
 b15zdnd11an1n64x5 FILLER_376_2006 ();
 b15zdnd11an1n64x5 FILLER_376_2070 ();
 b15zdnd11an1n16x5 FILLER_376_2134 ();
 b15zdnd11an1n04x5 FILLER_376_2150 ();
 b15zdnd11an1n64x5 FILLER_376_2162 ();
 b15zdnd11an1n32x5 FILLER_376_2226 ();
 b15zdnd11an1n16x5 FILLER_376_2258 ();
 b15zdnd00an1n02x5 FILLER_376_2274 ();
 b15zdnd11an1n64x5 FILLER_377_0 ();
 b15zdnd11an1n64x5 FILLER_377_64 ();
 b15zdnd11an1n64x5 FILLER_377_128 ();
 b15zdnd11an1n64x5 FILLER_377_192 ();
 b15zdnd11an1n64x5 FILLER_377_256 ();
 b15zdnd11an1n64x5 FILLER_377_320 ();
 b15zdnd11an1n64x5 FILLER_377_384 ();
 b15zdnd11an1n64x5 FILLER_377_448 ();
 b15zdnd11an1n64x5 FILLER_377_512 ();
 b15zdnd11an1n64x5 FILLER_377_576 ();
 b15zdnd11an1n64x5 FILLER_377_640 ();
 b15zdnd11an1n64x5 FILLER_377_704 ();
 b15zdnd11an1n64x5 FILLER_377_768 ();
 b15zdnd11an1n64x5 FILLER_377_832 ();
 b15zdnd11an1n64x5 FILLER_377_896 ();
 b15zdnd11an1n64x5 FILLER_377_960 ();
 b15zdnd11an1n64x5 FILLER_377_1024 ();
 b15zdnd11an1n64x5 FILLER_377_1088 ();
 b15zdnd11an1n64x5 FILLER_377_1152 ();
 b15zdnd11an1n64x5 FILLER_377_1216 ();
 b15zdnd11an1n64x5 FILLER_377_1280 ();
 b15zdnd11an1n64x5 FILLER_377_1344 ();
 b15zdnd11an1n64x5 FILLER_377_1408 ();
 b15zdnd11an1n64x5 FILLER_377_1472 ();
 b15zdnd11an1n64x5 FILLER_377_1536 ();
 b15zdnd11an1n64x5 FILLER_377_1600 ();
 b15zdnd11an1n64x5 FILLER_377_1664 ();
 b15zdnd11an1n64x5 FILLER_377_1728 ();
 b15zdnd11an1n64x5 FILLER_377_1792 ();
 b15zdnd11an1n64x5 FILLER_377_1856 ();
 b15zdnd11an1n64x5 FILLER_377_1920 ();
 b15zdnd11an1n64x5 FILLER_377_1984 ();
 b15zdnd11an1n64x5 FILLER_377_2048 ();
 b15zdnd11an1n64x5 FILLER_377_2112 ();
 b15zdnd11an1n64x5 FILLER_377_2176 ();
 b15zdnd11an1n32x5 FILLER_377_2240 ();
 b15zdnd11an1n08x5 FILLER_377_2272 ();
 b15zdnd11an1n04x5 FILLER_377_2280 ();
 b15zdnd11an1n64x5 FILLER_378_8 ();
 b15zdnd11an1n64x5 FILLER_378_72 ();
 b15zdnd11an1n64x5 FILLER_378_136 ();
 b15zdnd11an1n64x5 FILLER_378_200 ();
 b15zdnd11an1n64x5 FILLER_378_264 ();
 b15zdnd11an1n64x5 FILLER_378_328 ();
 b15zdnd11an1n64x5 FILLER_378_392 ();
 b15zdnd11an1n64x5 FILLER_378_456 ();
 b15zdnd11an1n64x5 FILLER_378_520 ();
 b15zdnd11an1n64x5 FILLER_378_584 ();
 b15zdnd11an1n64x5 FILLER_378_648 ();
 b15zdnd11an1n04x5 FILLER_378_712 ();
 b15zdnd00an1n02x5 FILLER_378_716 ();
 b15zdnd11an1n64x5 FILLER_378_726 ();
 b15zdnd11an1n64x5 FILLER_378_790 ();
 b15zdnd11an1n64x5 FILLER_378_854 ();
 b15zdnd11an1n64x5 FILLER_378_918 ();
 b15zdnd11an1n64x5 FILLER_378_982 ();
 b15zdnd11an1n64x5 FILLER_378_1046 ();
 b15zdnd11an1n64x5 FILLER_378_1110 ();
 b15zdnd11an1n64x5 FILLER_378_1174 ();
 b15zdnd11an1n64x5 FILLER_378_1238 ();
 b15zdnd11an1n64x5 FILLER_378_1302 ();
 b15zdnd11an1n64x5 FILLER_378_1366 ();
 b15zdnd11an1n64x5 FILLER_378_1430 ();
 b15zdnd11an1n64x5 FILLER_378_1494 ();
 b15zdnd11an1n64x5 FILLER_378_1558 ();
 b15zdnd11an1n64x5 FILLER_378_1622 ();
 b15zdnd11an1n64x5 FILLER_378_1686 ();
 b15zdnd11an1n64x5 FILLER_378_1750 ();
 b15zdnd11an1n64x5 FILLER_378_1814 ();
 b15zdnd11an1n64x5 FILLER_378_1878 ();
 b15zdnd11an1n64x5 FILLER_378_1942 ();
 b15zdnd11an1n64x5 FILLER_378_2006 ();
 b15zdnd11an1n64x5 FILLER_378_2070 ();
 b15zdnd11an1n16x5 FILLER_378_2134 ();
 b15zdnd11an1n04x5 FILLER_378_2150 ();
 b15zdnd11an1n64x5 FILLER_378_2162 ();
 b15zdnd11an1n32x5 FILLER_378_2226 ();
 b15zdnd11an1n16x5 FILLER_378_2258 ();
 b15zdnd00an1n02x5 FILLER_378_2274 ();
 b15zdnd11an1n64x5 FILLER_379_0 ();
 b15zdnd11an1n64x5 FILLER_379_64 ();
 b15zdnd11an1n64x5 FILLER_379_128 ();
 b15zdnd11an1n64x5 FILLER_379_192 ();
 b15zdnd11an1n64x5 FILLER_379_256 ();
 b15zdnd11an1n64x5 FILLER_379_320 ();
 b15zdnd11an1n64x5 FILLER_379_384 ();
 b15zdnd11an1n64x5 FILLER_379_448 ();
 b15zdnd11an1n64x5 FILLER_379_512 ();
 b15zdnd11an1n64x5 FILLER_379_576 ();
 b15zdnd11an1n64x5 FILLER_379_640 ();
 b15zdnd11an1n64x5 FILLER_379_704 ();
 b15zdnd11an1n64x5 FILLER_379_768 ();
 b15zdnd11an1n64x5 FILLER_379_832 ();
 b15zdnd11an1n64x5 FILLER_379_896 ();
 b15zdnd11an1n64x5 FILLER_379_960 ();
 b15zdnd11an1n64x5 FILLER_379_1024 ();
 b15zdnd11an1n64x5 FILLER_379_1088 ();
 b15zdnd11an1n64x5 FILLER_379_1152 ();
 b15zdnd11an1n64x5 FILLER_379_1216 ();
 b15zdnd11an1n64x5 FILLER_379_1280 ();
 b15zdnd11an1n64x5 FILLER_379_1344 ();
 b15zdnd11an1n64x5 FILLER_379_1408 ();
 b15zdnd11an1n64x5 FILLER_379_1472 ();
 b15zdnd11an1n64x5 FILLER_379_1536 ();
 b15zdnd11an1n64x5 FILLER_379_1600 ();
 b15zdnd11an1n64x5 FILLER_379_1664 ();
 b15zdnd11an1n64x5 FILLER_379_1728 ();
 b15zdnd11an1n64x5 FILLER_379_1792 ();
 b15zdnd11an1n64x5 FILLER_379_1856 ();
 b15zdnd11an1n64x5 FILLER_379_1920 ();
 b15zdnd11an1n64x5 FILLER_379_1984 ();
 b15zdnd11an1n64x5 FILLER_379_2048 ();
 b15zdnd11an1n64x5 FILLER_379_2112 ();
 b15zdnd11an1n64x5 FILLER_379_2176 ();
 b15zdnd11an1n32x5 FILLER_379_2240 ();
 b15zdnd11an1n08x5 FILLER_379_2272 ();
 b15zdnd11an1n04x5 FILLER_379_2280 ();
 b15zdnd11an1n64x5 FILLER_380_8 ();
 b15zdnd11an1n64x5 FILLER_380_72 ();
 b15zdnd11an1n64x5 FILLER_380_136 ();
 b15zdnd11an1n64x5 FILLER_380_200 ();
 b15zdnd11an1n64x5 FILLER_380_264 ();
 b15zdnd11an1n64x5 FILLER_380_328 ();
 b15zdnd11an1n64x5 FILLER_380_392 ();
 b15zdnd11an1n64x5 FILLER_380_456 ();
 b15zdnd11an1n64x5 FILLER_380_520 ();
 b15zdnd11an1n64x5 FILLER_380_584 ();
 b15zdnd11an1n64x5 FILLER_380_648 ();
 b15zdnd11an1n04x5 FILLER_380_712 ();
 b15zdnd00an1n02x5 FILLER_380_716 ();
 b15zdnd11an1n64x5 FILLER_380_726 ();
 b15zdnd11an1n64x5 FILLER_380_790 ();
 b15zdnd11an1n64x5 FILLER_380_854 ();
 b15zdnd11an1n64x5 FILLER_380_918 ();
 b15zdnd11an1n64x5 FILLER_380_982 ();
 b15zdnd11an1n64x5 FILLER_380_1046 ();
 b15zdnd11an1n64x5 FILLER_380_1110 ();
 b15zdnd11an1n64x5 FILLER_380_1174 ();
 b15zdnd11an1n64x5 FILLER_380_1238 ();
 b15zdnd11an1n64x5 FILLER_380_1302 ();
 b15zdnd11an1n64x5 FILLER_380_1366 ();
 b15zdnd11an1n64x5 FILLER_380_1430 ();
 b15zdnd11an1n64x5 FILLER_380_1494 ();
 b15zdnd11an1n64x5 FILLER_380_1558 ();
 b15zdnd11an1n64x5 FILLER_380_1622 ();
 b15zdnd11an1n64x5 FILLER_380_1686 ();
 b15zdnd11an1n64x5 FILLER_380_1750 ();
 b15zdnd11an1n64x5 FILLER_380_1814 ();
 b15zdnd11an1n64x5 FILLER_380_1878 ();
 b15zdnd11an1n64x5 FILLER_380_1942 ();
 b15zdnd11an1n64x5 FILLER_380_2006 ();
 b15zdnd11an1n64x5 FILLER_380_2070 ();
 b15zdnd11an1n16x5 FILLER_380_2134 ();
 b15zdnd11an1n04x5 FILLER_380_2150 ();
 b15zdnd11an1n64x5 FILLER_380_2162 ();
 b15zdnd11an1n32x5 FILLER_380_2226 ();
 b15zdnd11an1n16x5 FILLER_380_2258 ();
 b15zdnd00an1n02x5 FILLER_380_2274 ();
 b15zdnd11an1n64x5 FILLER_381_0 ();
 b15zdnd11an1n64x5 FILLER_381_64 ();
 b15zdnd11an1n64x5 FILLER_381_128 ();
 b15zdnd11an1n64x5 FILLER_381_192 ();
 b15zdnd11an1n64x5 FILLER_381_256 ();
 b15zdnd11an1n64x5 FILLER_381_320 ();
 b15zdnd11an1n64x5 FILLER_381_384 ();
 b15zdnd11an1n64x5 FILLER_381_448 ();
 b15zdnd11an1n64x5 FILLER_381_512 ();
 b15zdnd11an1n64x5 FILLER_381_576 ();
 b15zdnd11an1n64x5 FILLER_381_640 ();
 b15zdnd11an1n64x5 FILLER_381_704 ();
 b15zdnd11an1n64x5 FILLER_381_768 ();
 b15zdnd11an1n64x5 FILLER_381_832 ();
 b15zdnd11an1n64x5 FILLER_381_896 ();
 b15zdnd11an1n64x5 FILLER_381_960 ();
 b15zdnd11an1n64x5 FILLER_381_1024 ();
 b15zdnd11an1n64x5 FILLER_381_1088 ();
 b15zdnd11an1n64x5 FILLER_381_1152 ();
 b15zdnd11an1n64x5 FILLER_381_1216 ();
 b15zdnd11an1n64x5 FILLER_381_1280 ();
 b15zdnd11an1n64x5 FILLER_381_1344 ();
 b15zdnd11an1n64x5 FILLER_381_1408 ();
 b15zdnd11an1n64x5 FILLER_381_1472 ();
 b15zdnd11an1n64x5 FILLER_381_1536 ();
 b15zdnd11an1n64x5 FILLER_381_1600 ();
 b15zdnd11an1n64x5 FILLER_381_1664 ();
 b15zdnd11an1n64x5 FILLER_381_1728 ();
 b15zdnd11an1n64x5 FILLER_381_1792 ();
 b15zdnd11an1n64x5 FILLER_381_1856 ();
 b15zdnd11an1n64x5 FILLER_381_1920 ();
 b15zdnd11an1n64x5 FILLER_381_1984 ();
 b15zdnd11an1n64x5 FILLER_381_2048 ();
 b15zdnd11an1n64x5 FILLER_381_2112 ();
 b15zdnd11an1n64x5 FILLER_381_2176 ();
 b15zdnd11an1n32x5 FILLER_381_2240 ();
 b15zdnd11an1n08x5 FILLER_381_2272 ();
 b15zdnd11an1n04x5 FILLER_381_2280 ();
 b15zdnd11an1n64x5 FILLER_382_8 ();
 b15zdnd11an1n64x5 FILLER_382_72 ();
 b15zdnd11an1n64x5 FILLER_382_136 ();
 b15zdnd11an1n64x5 FILLER_382_200 ();
 b15zdnd11an1n64x5 FILLER_382_264 ();
 b15zdnd11an1n64x5 FILLER_382_328 ();
 b15zdnd11an1n64x5 FILLER_382_392 ();
 b15zdnd11an1n64x5 FILLER_382_456 ();
 b15zdnd11an1n64x5 FILLER_382_520 ();
 b15zdnd11an1n64x5 FILLER_382_584 ();
 b15zdnd11an1n64x5 FILLER_382_648 ();
 b15zdnd11an1n04x5 FILLER_382_712 ();
 b15zdnd00an1n02x5 FILLER_382_716 ();
 b15zdnd11an1n64x5 FILLER_382_726 ();
 b15zdnd11an1n64x5 FILLER_382_790 ();
 b15zdnd11an1n64x5 FILLER_382_854 ();
 b15zdnd11an1n64x5 FILLER_382_918 ();
 b15zdnd11an1n64x5 FILLER_382_982 ();
 b15zdnd11an1n64x5 FILLER_382_1046 ();
 b15zdnd11an1n64x5 FILLER_382_1110 ();
 b15zdnd11an1n64x5 FILLER_382_1174 ();
 b15zdnd11an1n64x5 FILLER_382_1238 ();
 b15zdnd11an1n64x5 FILLER_382_1302 ();
 b15zdnd11an1n64x5 FILLER_382_1366 ();
 b15zdnd11an1n64x5 FILLER_382_1430 ();
 b15zdnd11an1n64x5 FILLER_382_1494 ();
 b15zdnd11an1n64x5 FILLER_382_1558 ();
 b15zdnd11an1n64x5 FILLER_382_1622 ();
 b15zdnd11an1n64x5 FILLER_382_1686 ();
 b15zdnd11an1n64x5 FILLER_382_1750 ();
 b15zdnd11an1n64x5 FILLER_382_1814 ();
 b15zdnd11an1n64x5 FILLER_382_1878 ();
 b15zdnd11an1n64x5 FILLER_382_1942 ();
 b15zdnd11an1n64x5 FILLER_382_2006 ();
 b15zdnd11an1n64x5 FILLER_382_2070 ();
 b15zdnd11an1n16x5 FILLER_382_2134 ();
 b15zdnd11an1n04x5 FILLER_382_2150 ();
 b15zdnd11an1n64x5 FILLER_382_2162 ();
 b15zdnd11an1n32x5 FILLER_382_2226 ();
 b15zdnd11an1n16x5 FILLER_382_2258 ();
 b15zdnd00an1n02x5 FILLER_382_2274 ();
 b15zdnd11an1n64x5 FILLER_383_0 ();
 b15zdnd11an1n64x5 FILLER_383_64 ();
 b15zdnd11an1n64x5 FILLER_383_128 ();
 b15zdnd11an1n64x5 FILLER_383_192 ();
 b15zdnd11an1n64x5 FILLER_383_256 ();
 b15zdnd11an1n64x5 FILLER_383_320 ();
 b15zdnd11an1n64x5 FILLER_383_384 ();
 b15zdnd11an1n64x5 FILLER_383_448 ();
 b15zdnd11an1n64x5 FILLER_383_512 ();
 b15zdnd11an1n64x5 FILLER_383_576 ();
 b15zdnd11an1n64x5 FILLER_383_640 ();
 b15zdnd11an1n64x5 FILLER_383_704 ();
 b15zdnd11an1n64x5 FILLER_383_768 ();
 b15zdnd11an1n64x5 FILLER_383_832 ();
 b15zdnd11an1n64x5 FILLER_383_896 ();
 b15zdnd11an1n64x5 FILLER_383_960 ();
 b15zdnd11an1n64x5 FILLER_383_1024 ();
 b15zdnd11an1n64x5 FILLER_383_1088 ();
 b15zdnd11an1n64x5 FILLER_383_1152 ();
 b15zdnd11an1n64x5 FILLER_383_1216 ();
 b15zdnd11an1n64x5 FILLER_383_1280 ();
 b15zdnd11an1n64x5 FILLER_383_1344 ();
 b15zdnd11an1n64x5 FILLER_383_1408 ();
 b15zdnd11an1n64x5 FILLER_383_1472 ();
 b15zdnd11an1n64x5 FILLER_383_1536 ();
 b15zdnd11an1n64x5 FILLER_383_1600 ();
 b15zdnd11an1n64x5 FILLER_383_1664 ();
 b15zdnd11an1n64x5 FILLER_383_1728 ();
 b15zdnd11an1n64x5 FILLER_383_1792 ();
 b15zdnd11an1n64x5 FILLER_383_1856 ();
 b15zdnd11an1n64x5 FILLER_383_1920 ();
 b15zdnd11an1n64x5 FILLER_383_1984 ();
 b15zdnd11an1n64x5 FILLER_383_2048 ();
 b15zdnd11an1n64x5 FILLER_383_2112 ();
 b15zdnd11an1n64x5 FILLER_383_2176 ();
 b15zdnd11an1n32x5 FILLER_383_2240 ();
 b15zdnd11an1n08x5 FILLER_383_2272 ();
 b15zdnd11an1n04x5 FILLER_383_2280 ();
 b15zdnd11an1n64x5 FILLER_384_8 ();
 b15zdnd11an1n64x5 FILLER_384_72 ();
 b15zdnd11an1n64x5 FILLER_384_136 ();
 b15zdnd11an1n64x5 FILLER_384_200 ();
 b15zdnd11an1n64x5 FILLER_384_264 ();
 b15zdnd11an1n64x5 FILLER_384_328 ();
 b15zdnd11an1n64x5 FILLER_384_392 ();
 b15zdnd11an1n64x5 FILLER_384_456 ();
 b15zdnd11an1n64x5 FILLER_384_520 ();
 b15zdnd11an1n64x5 FILLER_384_584 ();
 b15zdnd11an1n64x5 FILLER_384_648 ();
 b15zdnd11an1n04x5 FILLER_384_712 ();
 b15zdnd00an1n02x5 FILLER_384_716 ();
 b15zdnd11an1n64x5 FILLER_384_726 ();
 b15zdnd11an1n64x5 FILLER_384_790 ();
 b15zdnd11an1n64x5 FILLER_384_854 ();
 b15zdnd11an1n64x5 FILLER_384_918 ();
 b15zdnd11an1n64x5 FILLER_384_982 ();
 b15zdnd11an1n64x5 FILLER_384_1046 ();
 b15zdnd11an1n64x5 FILLER_384_1110 ();
 b15zdnd11an1n64x5 FILLER_384_1174 ();
 b15zdnd11an1n64x5 FILLER_384_1238 ();
 b15zdnd11an1n64x5 FILLER_384_1302 ();
 b15zdnd11an1n64x5 FILLER_384_1366 ();
 b15zdnd11an1n64x5 FILLER_384_1430 ();
 b15zdnd11an1n64x5 FILLER_384_1494 ();
 b15zdnd11an1n64x5 FILLER_384_1558 ();
 b15zdnd11an1n64x5 FILLER_384_1622 ();
 b15zdnd11an1n64x5 FILLER_384_1686 ();
 b15zdnd11an1n64x5 FILLER_384_1750 ();
 b15zdnd11an1n64x5 FILLER_384_1814 ();
 b15zdnd11an1n64x5 FILLER_384_1878 ();
 b15zdnd11an1n64x5 FILLER_384_1942 ();
 b15zdnd11an1n64x5 FILLER_384_2006 ();
 b15zdnd11an1n64x5 FILLER_384_2070 ();
 b15zdnd11an1n16x5 FILLER_384_2134 ();
 b15zdnd11an1n04x5 FILLER_384_2150 ();
 b15zdnd11an1n64x5 FILLER_384_2162 ();
 b15zdnd11an1n32x5 FILLER_384_2226 ();
 b15zdnd11an1n16x5 FILLER_384_2258 ();
 b15zdnd00an1n02x5 FILLER_384_2274 ();
 b15zdnd11an1n64x5 FILLER_385_0 ();
 b15zdnd11an1n64x5 FILLER_385_64 ();
 b15zdnd11an1n64x5 FILLER_385_128 ();
 b15zdnd11an1n64x5 FILLER_385_192 ();
 b15zdnd11an1n64x5 FILLER_385_256 ();
 b15zdnd11an1n64x5 FILLER_385_320 ();
 b15zdnd11an1n64x5 FILLER_385_384 ();
 b15zdnd11an1n64x5 FILLER_385_448 ();
 b15zdnd11an1n64x5 FILLER_385_512 ();
 b15zdnd11an1n64x5 FILLER_385_576 ();
 b15zdnd11an1n64x5 FILLER_385_640 ();
 b15zdnd11an1n64x5 FILLER_385_704 ();
 b15zdnd11an1n64x5 FILLER_385_768 ();
 b15zdnd11an1n64x5 FILLER_385_832 ();
 b15zdnd11an1n64x5 FILLER_385_896 ();
 b15zdnd11an1n64x5 FILLER_385_960 ();
 b15zdnd11an1n64x5 FILLER_385_1024 ();
 b15zdnd11an1n64x5 FILLER_385_1088 ();
 b15zdnd11an1n64x5 FILLER_385_1152 ();
 b15zdnd11an1n64x5 FILLER_385_1216 ();
 b15zdnd11an1n64x5 FILLER_385_1280 ();
 b15zdnd11an1n64x5 FILLER_385_1344 ();
 b15zdnd11an1n64x5 FILLER_385_1408 ();
 b15zdnd11an1n64x5 FILLER_385_1472 ();
 b15zdnd11an1n64x5 FILLER_385_1536 ();
 b15zdnd11an1n64x5 FILLER_385_1600 ();
 b15zdnd11an1n64x5 FILLER_385_1664 ();
 b15zdnd11an1n64x5 FILLER_385_1728 ();
 b15zdnd11an1n64x5 FILLER_385_1792 ();
 b15zdnd11an1n64x5 FILLER_385_1856 ();
 b15zdnd11an1n64x5 FILLER_385_1920 ();
 b15zdnd11an1n64x5 FILLER_385_1984 ();
 b15zdnd11an1n64x5 FILLER_385_2048 ();
 b15zdnd11an1n64x5 FILLER_385_2112 ();
 b15zdnd11an1n64x5 FILLER_385_2176 ();
 b15zdnd11an1n32x5 FILLER_385_2240 ();
 b15zdnd11an1n08x5 FILLER_385_2272 ();
 b15zdnd11an1n04x5 FILLER_385_2280 ();
 b15zdnd11an1n64x5 FILLER_386_8 ();
 b15zdnd11an1n64x5 FILLER_386_72 ();
 b15zdnd11an1n64x5 FILLER_386_136 ();
 b15zdnd11an1n64x5 FILLER_386_200 ();
 b15zdnd11an1n64x5 FILLER_386_264 ();
 b15zdnd11an1n64x5 FILLER_386_328 ();
 b15zdnd11an1n64x5 FILLER_386_392 ();
 b15zdnd11an1n64x5 FILLER_386_456 ();
 b15zdnd11an1n64x5 FILLER_386_520 ();
 b15zdnd11an1n64x5 FILLER_386_584 ();
 b15zdnd11an1n64x5 FILLER_386_648 ();
 b15zdnd11an1n04x5 FILLER_386_712 ();
 b15zdnd00an1n02x5 FILLER_386_716 ();
 b15zdnd11an1n64x5 FILLER_386_726 ();
 b15zdnd11an1n64x5 FILLER_386_790 ();
 b15zdnd11an1n64x5 FILLER_386_854 ();
 b15zdnd11an1n64x5 FILLER_386_918 ();
 b15zdnd11an1n08x5 FILLER_386_982 ();
 b15zdnd11an1n04x5 FILLER_386_990 ();
 b15zdnd00an1n02x5 FILLER_386_994 ();
 b15zdnd00an1n01x5 FILLER_386_996 ();
 b15zdnd11an1n16x5 FILLER_386_1001 ();
 b15zdnd11an1n04x5 FILLER_386_1017 ();
 b15zdnd00an1n02x5 FILLER_386_1021 ();
 b15zdnd11an1n64x5 FILLER_386_1027 ();
 b15zdnd11an1n64x5 FILLER_386_1091 ();
 b15zdnd11an1n64x5 FILLER_386_1155 ();
 b15zdnd11an1n64x5 FILLER_386_1219 ();
 b15zdnd11an1n64x5 FILLER_386_1283 ();
 b15zdnd11an1n64x5 FILLER_386_1347 ();
 b15zdnd11an1n64x5 FILLER_386_1411 ();
 b15zdnd11an1n64x5 FILLER_386_1475 ();
 b15zdnd11an1n64x5 FILLER_386_1539 ();
 b15zdnd11an1n64x5 FILLER_386_1603 ();
 b15zdnd11an1n64x5 FILLER_386_1667 ();
 b15zdnd11an1n64x5 FILLER_386_1731 ();
 b15zdnd11an1n64x5 FILLER_386_1795 ();
 b15zdnd11an1n64x5 FILLER_386_1859 ();
 b15zdnd11an1n64x5 FILLER_386_1923 ();
 b15zdnd11an1n64x5 FILLER_386_1987 ();
 b15zdnd11an1n64x5 FILLER_386_2051 ();
 b15zdnd11an1n32x5 FILLER_386_2115 ();
 b15zdnd11an1n04x5 FILLER_386_2147 ();
 b15zdnd00an1n02x5 FILLER_386_2151 ();
 b15zdnd00an1n01x5 FILLER_386_2153 ();
 b15zdnd11an1n64x5 FILLER_386_2162 ();
 b15zdnd11an1n32x5 FILLER_386_2226 ();
 b15zdnd11an1n16x5 FILLER_386_2258 ();
 b15zdnd00an1n02x5 FILLER_386_2274 ();
 b15zdnd11an1n64x5 FILLER_387_0 ();
 b15zdnd11an1n64x5 FILLER_387_64 ();
 b15zdnd11an1n64x5 FILLER_387_128 ();
 b15zdnd11an1n64x5 FILLER_387_192 ();
 b15zdnd11an1n64x5 FILLER_387_256 ();
 b15zdnd11an1n64x5 FILLER_387_320 ();
 b15zdnd11an1n64x5 FILLER_387_384 ();
 b15zdnd11an1n64x5 FILLER_387_448 ();
 b15zdnd11an1n64x5 FILLER_387_512 ();
 b15zdnd11an1n64x5 FILLER_387_576 ();
 b15zdnd11an1n64x5 FILLER_387_640 ();
 b15zdnd11an1n64x5 FILLER_387_704 ();
 b15zdnd11an1n64x5 FILLER_387_768 ();
 b15zdnd11an1n64x5 FILLER_387_832 ();
 b15zdnd11an1n16x5 FILLER_387_896 ();
 b15zdnd11an1n04x5 FILLER_387_912 ();
 b15zdnd11an1n32x5 FILLER_387_958 ();
 b15zdnd11an1n04x5 FILLER_387_990 ();
 b15zdnd00an1n02x5 FILLER_387_994 ();
 b15zdnd11an1n64x5 FILLER_387_1038 ();
 b15zdnd11an1n64x5 FILLER_387_1102 ();
 b15zdnd11an1n64x5 FILLER_387_1166 ();
 b15zdnd11an1n64x5 FILLER_387_1230 ();
 b15zdnd11an1n64x5 FILLER_387_1294 ();
 b15zdnd11an1n64x5 FILLER_387_1358 ();
 b15zdnd11an1n64x5 FILLER_387_1422 ();
 b15zdnd11an1n64x5 FILLER_387_1486 ();
 b15zdnd11an1n64x5 FILLER_387_1550 ();
 b15zdnd11an1n64x5 FILLER_387_1614 ();
 b15zdnd11an1n64x5 FILLER_387_1678 ();
 b15zdnd11an1n64x5 FILLER_387_1742 ();
 b15zdnd11an1n64x5 FILLER_387_1806 ();
 b15zdnd11an1n64x5 FILLER_387_1870 ();
 b15zdnd11an1n64x5 FILLER_387_1934 ();
 b15zdnd11an1n64x5 FILLER_387_1998 ();
 b15zdnd11an1n64x5 FILLER_387_2062 ();
 b15zdnd11an1n64x5 FILLER_387_2126 ();
 b15zdnd11an1n64x5 FILLER_387_2190 ();
 b15zdnd11an1n16x5 FILLER_387_2254 ();
 b15zdnd11an1n08x5 FILLER_387_2270 ();
 b15zdnd11an1n04x5 FILLER_387_2278 ();
 b15zdnd00an1n02x5 FILLER_387_2282 ();
 b15zdnd11an1n64x5 FILLER_388_8 ();
 b15zdnd11an1n64x5 FILLER_388_72 ();
 b15zdnd11an1n64x5 FILLER_388_136 ();
 b15zdnd11an1n64x5 FILLER_388_200 ();
 b15zdnd11an1n64x5 FILLER_388_264 ();
 b15zdnd11an1n64x5 FILLER_388_328 ();
 b15zdnd11an1n64x5 FILLER_388_392 ();
 b15zdnd11an1n64x5 FILLER_388_456 ();
 b15zdnd11an1n64x5 FILLER_388_520 ();
 b15zdnd11an1n64x5 FILLER_388_584 ();
 b15zdnd11an1n64x5 FILLER_388_648 ();
 b15zdnd11an1n04x5 FILLER_388_712 ();
 b15zdnd00an1n02x5 FILLER_388_716 ();
 b15zdnd11an1n64x5 FILLER_388_726 ();
 b15zdnd11an1n08x5 FILLER_388_790 ();
 b15zdnd11an1n04x5 FILLER_388_798 ();
 b15zdnd00an1n02x5 FILLER_388_802 ();
 b15zdnd11an1n64x5 FILLER_388_808 ();
 b15zdnd11an1n32x5 FILLER_388_872 ();
 b15zdnd11an1n08x5 FILLER_388_904 ();
 b15zdnd00an1n01x5 FILLER_388_912 ();
 b15zdnd11an1n04x5 FILLER_388_917 ();
 b15zdnd11an1n32x5 FILLER_388_963 ();
 b15zdnd11an1n08x5 FILLER_388_995 ();
 b15zdnd00an1n01x5 FILLER_388_1003 ();
 b15zdnd11an1n64x5 FILLER_388_1046 ();
 b15zdnd11an1n64x5 FILLER_388_1110 ();
 b15zdnd11an1n64x5 FILLER_388_1174 ();
 b15zdnd11an1n64x5 FILLER_388_1238 ();
 b15zdnd11an1n32x5 FILLER_388_1302 ();
 b15zdnd00an1n02x5 FILLER_388_1334 ();
 b15zdnd11an1n64x5 FILLER_388_1340 ();
 b15zdnd11an1n64x5 FILLER_388_1404 ();
 b15zdnd11an1n64x5 FILLER_388_1468 ();
 b15zdnd11an1n64x5 FILLER_388_1532 ();
 b15zdnd11an1n64x5 FILLER_388_1596 ();
 b15zdnd11an1n64x5 FILLER_388_1660 ();
 b15zdnd11an1n64x5 FILLER_388_1724 ();
 b15zdnd11an1n64x5 FILLER_388_1788 ();
 b15zdnd11an1n64x5 FILLER_388_1852 ();
 b15zdnd11an1n64x5 FILLER_388_1916 ();
 b15zdnd11an1n64x5 FILLER_388_1980 ();
 b15zdnd11an1n64x5 FILLER_388_2044 ();
 b15zdnd11an1n32x5 FILLER_388_2108 ();
 b15zdnd11an1n08x5 FILLER_388_2140 ();
 b15zdnd11an1n04x5 FILLER_388_2148 ();
 b15zdnd00an1n02x5 FILLER_388_2152 ();
 b15zdnd11an1n64x5 FILLER_388_2162 ();
 b15zdnd11an1n32x5 FILLER_388_2226 ();
 b15zdnd11an1n16x5 FILLER_388_2258 ();
 b15zdnd00an1n02x5 FILLER_388_2274 ();
 b15zdnd11an1n64x5 FILLER_389_0 ();
 b15zdnd11an1n64x5 FILLER_389_64 ();
 b15zdnd11an1n64x5 FILLER_389_128 ();
 b15zdnd11an1n64x5 FILLER_389_192 ();
 b15zdnd11an1n64x5 FILLER_389_256 ();
 b15zdnd11an1n64x5 FILLER_389_320 ();
 b15zdnd11an1n64x5 FILLER_389_384 ();
 b15zdnd11an1n64x5 FILLER_389_448 ();
 b15zdnd11an1n64x5 FILLER_389_512 ();
 b15zdnd11an1n64x5 FILLER_389_576 ();
 b15zdnd11an1n64x5 FILLER_389_640 ();
 b15zdnd11an1n64x5 FILLER_389_704 ();
 b15zdnd11an1n64x5 FILLER_389_768 ();
 b15zdnd11an1n64x5 FILLER_389_832 ();
 b15zdnd11an1n08x5 FILLER_389_896 ();
 b15zdnd11an1n04x5 FILLER_389_904 ();
 b15zdnd00an1n02x5 FILLER_389_908 ();
 b15zdnd11an1n04x5 FILLER_389_914 ();
 b15zdnd11an1n04x5 FILLER_389_922 ();
 b15zdnd11an1n32x5 FILLER_389_968 ();
 b15zdnd00an1n02x5 FILLER_389_1000 ();
 b15zdnd11an1n04x5 FILLER_389_1006 ();
 b15zdnd11an1n64x5 FILLER_389_1052 ();
 b15zdnd11an1n64x5 FILLER_389_1116 ();
 b15zdnd11an1n64x5 FILLER_389_1180 ();
 b15zdnd11an1n32x5 FILLER_389_1244 ();
 b15zdnd11an1n08x5 FILLER_389_1276 ();
 b15zdnd11an1n08x5 FILLER_389_1288 ();
 b15zdnd00an1n01x5 FILLER_389_1296 ();
 b15zdnd11an1n04x5 FILLER_389_1339 ();
 b15zdnd11an1n64x5 FILLER_389_1385 ();
 b15zdnd11an1n64x5 FILLER_389_1449 ();
 b15zdnd11an1n64x5 FILLER_389_1513 ();
 b15zdnd11an1n64x5 FILLER_389_1577 ();
 b15zdnd11an1n64x5 FILLER_389_1641 ();
 b15zdnd11an1n64x5 FILLER_389_1705 ();
 b15zdnd11an1n64x5 FILLER_389_1769 ();
 b15zdnd11an1n64x5 FILLER_389_1833 ();
 b15zdnd11an1n64x5 FILLER_389_1897 ();
 b15zdnd11an1n64x5 FILLER_389_1961 ();
 b15zdnd11an1n64x5 FILLER_389_2025 ();
 b15zdnd11an1n64x5 FILLER_389_2089 ();
 b15zdnd11an1n64x5 FILLER_389_2153 ();
 b15zdnd11an1n64x5 FILLER_389_2217 ();
 b15zdnd00an1n02x5 FILLER_389_2281 ();
 b15zdnd00an1n01x5 FILLER_389_2283 ();
endmodule
