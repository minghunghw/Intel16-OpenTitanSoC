
module dhm_lut (
        clk,
        reset_n,
        d_in,
        xor_out
);

input           clk;
input           reset_n;
input   [63:0]  d_in;
output          xor_out;

reg             xor_out;

////////////////////////////////////////////////////////////////////////////////

parameter LUT_WIDTH_IN  = 4;
parameter LUT_WIDTH_OUT = 4;

reg     [63:0]  lut_in;
reg     [63:0]  lut_out;
reg     [63:0]  lut;

// If lut_width=0, lut_mask=b00000000
// If lut_width=1, lut_mask=b00000001
// If lut_width=2, lut_mask=b00000011

wire    [63:0]  lut_mask_in  = (1 << LUT_WIDTH_IN  ) - 1;
wire    [63:0]  lut_mask_out = (1 << LUT_WIDTH_OUT ) - 1;

always @(posedge clk or negedge reset_n)
  begin
    if (!reset_n)
      begin
        lut_in  <= 0;
        lut_out <= 0;
        xor_out <= 0;
      end
    else
      begin
        lut_in  <= d_in & lut_mask_in;
        lut_out <= lut  & lut_mask_out;
        xor_out <= ^lut_out;
      end
  end

// Note that case content was generated by dhm_lut.tcl

always @ (lut_in or lut_mask_in)
  begin  
    case (lut_in)

      (64'he11b7f6503720372 & lut_mask_in) : lut = 64'h700b484f288dc659;
      (64'h8925fcb062156215 & lut_mask_in) : lut = 64'h43b991c1f4fbdd68;
      (64'h96e3271b6a266a26 & lut_mask_in) : lut = 64'hecb6b95e23451733;
      (64'hcbe0be7c11591159 & lut_mask_in) : lut = 64'h195e753da998e132;
      (64'h62f56d99fe3dfe3d & lut_mask_in) : lut = 64'h1a9abcb1f711e772;
      (64'h29e4838b7bfb7bfb & lut_mask_in) : lut = 64'h4546525859524b09;
      (64'h5f360611c3edc3ed & lut_mask_in) : lut = 64'h258f4692df6c0cab;
      (64'h7d23f82508260826 & lut_mask_in) : lut = 64'hd221294e1a1098a7;
      (64'hd6877e0207eb07eb & lut_mask_in) : lut = 64'h8f32c9adbae36efd;
      (64'h97ad4133eec1eec1 & lut_mask_in) : lut = 64'hcef0678673d40a9b;
      (64'h5bc60b6de34ce34c & lut_mask_in) : lut = 64'hc454a7fc5808474e;
      (64'hb60689cf97619761 & lut_mask_in) : lut = 64'h9c7bcb27de7864f4;
      (64'h1b9c6ef37a917a91 & lut_mask_in) : lut = 64'h97ebd23cc631b5a6;
      (64'h6396dc60d556d556 & lut_mask_in) : lut = 64'he7aadd02f1ae2ce3;
      (64'h8f3b6b8f2fb32fb3 & lut_mask_in) : lut = 64'h77342315b6a17184;
      (64'h5f5027d2bc53bc53 & lut_mask_in) : lut = 64'h6db5ab8405dfa2d7;
      (64'hc9d19d3b1d741d74 & lut_mask_in) : lut = 64'he26e95063773f80d;
      (64'h805cc5cab2dbb2db & lut_mask_in) : lut = 64'h0125ac125778389b;
      (64'h530d35065b085b08 & lut_mask_in) : lut = 64'h3a9942b7584595f6;
      (64'h44db1351a367a367 & lut_mask_in) : lut = 64'hbbf69292633e9072;
      (64'h1b1544e1e880e880 & lut_mask_in) : lut = 64'h5dc42227a4421f6a;
      (64'h681c0f0e4b434b43 & lut_mask_in) : lut = 64'hb22df4e4c9b24467;
      (64'hd978cf8743d543d5 & lut_mask_in) : lut = 64'hc336af06301c6329;
      (64'h0051255560a360a3 & lut_mask_in) : lut = 64'hb27d02990fa4f843;
      (64'hc516377c8aa78aa7 & lut_mask_in) : lut = 64'hc72fceb126982b27;
      (64'h3dede0fd02600260 & lut_mask_in) : lut = 64'h749cc4b5a60dc634;
      (64'h53e2e186ffdcffdc & lut_mask_in) : lut = 64'ha2dc7b996b8f4f2a;
      (64'h48764ade034d034d & lut_mask_in) : lut = 64'h1e9e6ddecb1f6989;
      (64'h8c8a46d9d7add7ad & lut_mask_in) : lut = 64'h3b3efd6a5f61e00c;
      (64'h94636646da3bda3b & lut_mask_in) : lut = 64'h4d06cb7c5886f67c;
      (64'hac51d069778e778e & lut_mask_in) : lut = 64'hbcd594cbca553619;
      (64'h29a145d70db90db9 & lut_mask_in) : lut = 64'h8c40f20acf5d4467;
      (64'h83e6df8cfa0cfa0c & lut_mask_in) : lut = 64'hd012835b3ae89a9b;
      (64'h8b8d7514325e325e & lut_mask_in) : lut = 64'he300c7b307f6e118;
      (64'hc7c33579db62db62 & lut_mask_in) : lut = 64'h6dabd6557341f064;
      (64'hde2b127524eb24eb & lut_mask_in) : lut = 64'h8840ec489bcd0c74;
      (64'hc61b29edccf8ccf8 & lut_mask_in) : lut = 64'hda6efa97ceb546b7;
      (64'hec3185a8bab9bab9 & lut_mask_in) : lut = 64'hc5f98edae533a89d;
      (64'h2cca745bfc5cfc5c & lut_mask_in) : lut = 64'hb9d77aee0e628703;
      (64'hd7b5f4872ef32ef3 & lut_mask_in) : lut = 64'hf2b7f76091d0ea22;
      (64'h1966d6eb7ff07ff0 & lut_mask_in) : lut = 64'h9bd976aecaaea5da;
      (64'h6734d84478487848 & lut_mask_in) : lut = 64'h9f1cbc782b418b09;
      (64'hbd371930f892f892 & lut_mask_in) : lut = 64'h170f1b11e30391eb;
      (64'h8b77050c73657365 & lut_mask_in) : lut = 64'h03290e499e513bb7;
      (64'hdf23a96318851885 & lut_mask_in) : lut = 64'h7ee7f9c703369398;
      (64'hbde19afaf95df95d & lut_mask_in) : lut = 64'h933d459202f1000f;
      (64'h3da1a10063e663e6 & lut_mask_in) : lut = 64'h863d41cb48562891;
      (64'h97820f64ae40ae40 & lut_mask_in) : lut = 64'h670f59a1427d1831;
      (64'habac30c406d306d3 & lut_mask_in) : lut = 64'h722fca7b4af3cc37;
      (64'h0bc798513b323b32 & lut_mask_in) : lut = 64'hb555ab08fe6563ff;
      (64'h765c02da77ff77ff & lut_mask_in) : lut = 64'h6e6cc069dd92a749;
      (64'h9a59818e19131913 & lut_mask_in) : lut = 64'h1aba45817d586433;
      (64'hbecab8416a586a58 & lut_mask_in) : lut = 64'ha9e992d042a5f096;
      (64'hf4520583cbd9cbd9 & lut_mask_in) : lut = 64'h18a9e724c4174157;
      (64'h23a7262050ff50ff & lut_mask_in) : lut = 64'h52a7437f9389ccc4;
      (64'h85e28065c74ec74e & lut_mask_in) : lut = 64'ha4374393cc5ef90d;
      (64'h41142992d418d418 & lut_mask_in) : lut = 64'hf0823beb8f97ad77;
      (64'h6e0ff9367cb57cb5 & lut_mask_in) : lut = 64'h6234187f9a0aaaec;
      (64'h912d47ea5e795e79 & lut_mask_in) : lut = 64'hb0e8953845f32598;
      (64'h2e4287139a549a54 & lut_mask_in) : lut = 64'hb5a2088a7c8106ad;
      (64'h211e9fef06360636 & lut_mask_in) : lut = 64'h13dbee2ed55159d9;
      (64'h5c2e986acfa5cfa5 & lut_mask_in) : lut = 64'hccb8605af1a4001b;
      (64'h99ae7eb45b155b15 & lut_mask_in) : lut = 64'h04d6012c25c6a988;
      (64'haf2a887cce5dce5d & lut_mask_in) : lut = 64'h9f31f77eadf21934;
      (64'h9b3e60b3465e465e & lut_mask_in) : lut = 64'hc2c9820300a12f57;
      (64'h2ba3578adc1cdc1c & lut_mask_in) : lut = 64'h7b417340305e0ee6;
      (64'hc3effbcef375f375 & lut_mask_in) : lut = 64'h5e6a297383fc8cd7;
      (64'hb530b32ec6fbc6fb & lut_mask_in) : lut = 64'hf4c72d9209ef8113;
      (64'h435a4635ae4bae4b & lut_mask_in) : lut = 64'h3fd7f37f8cc9cfad;
      (64'h60894247d5ced5ce & lut_mask_in) : lut = 64'h6cfa4626d3c1dc6a;
      (64'h6a4998faf60cf60c & lut_mask_in) : lut = 64'h9a1dd8f86a73fe93;
      (64'h4058f31ab496b496 & lut_mask_in) : lut = 64'hfac5eb96d66a7515;
      (64'h446fb36f12e112e1 & lut_mask_in) : lut = 64'h0a2b65e6a642d67c;
      (64'h5df5926d896f896f & lut_mask_in) : lut = 64'h418ddec0b80e9592;
      (64'hb33ab34df50af50a & lut_mask_in) : lut = 64'h96a0e73d7baad070;
      (64'h8df2ed936b066b06 & lut_mask_in) : lut = 64'h4163e11dcb6e3650;
      (64'h015be4db6b346b34 & lut_mask_in) : lut = 64'hdff0d1c1391d246c;
      (64'h29610a0a61b161b1 & lut_mask_in) : lut = 64'hac2af2e503edc15a;
      (64'hcd98360ad640d640 & lut_mask_in) : lut = 64'h6f4e8ac0071bd043;
      (64'h458b71bd3d743d74 & lut_mask_in) : lut = 64'h03487de07bd7cfb5;
      (64'h4d0fa94eb9e8b9e8 & lut_mask_in) : lut = 64'h1866472d08ca4473;
      (64'h8f5cee376e7e6e7e & lut_mask_in) : lut = 64'h624a3c5acfee10fe;
      (64'he1aa0a6a1ddf1ddf & lut_mask_in) : lut = 64'h2be8e6e2a0969830;
      (64'heac2af0239523952 & lut_mask_in) : lut = 64'h8d77b3e92e2575fc;
      (64'h3b6bc1244f414f41 & lut_mask_in) : lut = 64'h80fa9f1efb8f112a;
      (64'h6fd8a8dd3eab3eab & lut_mask_in) : lut = 64'h06629d2583a0e183;
      (64'h254b184860856085 & lut_mask_in) : lut = 64'h541bd1bb3afd946f;
      (64'hff04c6aecebaceba & lut_mask_in) : lut = 64'h4d8c46f4db288abe;
      (64'h9bd24da550925092 & lut_mask_in) : lut = 64'hc4240be470983627;
      (64'h1fad348dc675c675 & lut_mask_in) : lut = 64'h7ff2997bdb0e97b8;
      (64'haf39f98548884888 & lut_mask_in) : lut = 64'h2232978add280437;
      (64'h84303f20ff10ff10 & lut_mask_in) : lut = 64'hd95c8416e638910c;
      (64'h5b17628ea203a203 & lut_mask_in) : lut = 64'heecf4e989c194491;
      (64'h9daf722b99d599d5 & lut_mask_in) : lut = 64'h268927cdf15d538f;
      (64'hf7020248826d826d & lut_mask_in) : lut = 64'h8f29752b11d0e16e;
      (64'he5670a4fd589d589 & lut_mask_in) : lut = 64'hd6dca4d99bb1ce04;
      (64'h56c3198c330e330e & lut_mask_in) : lut = 64'h8a546d8a88251d96;
      (64'hc63cb5dd09360936 & lut_mask_in) : lut = 64'h769ec5fde840cc87;
      (64'h908ca8afbae1bae1 & lut_mask_in) : lut = 64'h19ad00c33e1df9ba;
      (64'h9474dcc332aa32aa & lut_mask_in) : lut = 64'hef40c1de26af5a6e;
      (64'hf5a5836f4b0e4b0e & lut_mask_in) : lut = 64'he395eb9ef62434bf;
      (64'h51f88051c535c535 & lut_mask_in) : lut = 64'hb3f2bf1f00e18b8d;
      (64'h0741e99436f936f9 & lut_mask_in) : lut = 64'h3206f5c8413c594e;
      (64'hf2f565804f294f29 & lut_mask_in) : lut = 64'h09d10f817b9fe3a1;
      (64'h4711b2330f870f87 & lut_mask_in) : lut = 64'hf9f33155c839e5db;
      (64'h0c2cd0c88ebe8ebe & lut_mask_in) : lut = 64'h7d3217eb400d5dff;
      (64'hde4a8b336abb6abb & lut_mask_in) : lut = 64'h08d490dedb68dccf;
      (64'h2880b3f71dae1dae & lut_mask_in) : lut = 64'hc88d43f917c3f34c;
      (64'hdd4aae47af7faf7f & lut_mask_in) : lut = 64'h277d0758eeb646e7;
      (64'h1913b297f5bff5bf & lut_mask_in) : lut = 64'h68cc6645d06465a3;
      (64'h26ea5bb6e4a1e4a1 & lut_mask_in) : lut = 64'h37ae5b64f31adc7a;
      (64'hb271826822d922d9 & lut_mask_in) : lut = 64'h82f35ea0a6615657;
      (64'hc08c26a3ff6fff6f & lut_mask_in) : lut = 64'h4ec96631b1695159;
      (64'hd29f737807290729 & lut_mask_in) : lut = 64'h2f36cfb7a03cc5d3;
      (64'h55bc8b3125e725e7 & lut_mask_in) : lut = 64'hc02bceb8d21ac5e7;
      (64'hc90c521885e185e1 & lut_mask_in) : lut = 64'hd0d95625f78d3f2a;
      (64'h971d56a9a42ea42e & lut_mask_in) : lut = 64'h4bfdc8453386faee;
      (64'h05570522fd38fd38 & lut_mask_in) : lut = 64'h1e07b7f0a3d4b28e;
      (64'hcd2a874c94009400 & lut_mask_in) : lut = 64'h5d86db30fd9380e4;
      (64'hdeda29cbae37ae37 & lut_mask_in) : lut = 64'h1d5660d4e758f7ba;
      (64'ha34e04deaccbaccb & lut_mask_in) : lut = 64'h201e60738c886799;
      (64'h2e32c0f55caf5caf & lut_mask_in) : lut = 64'h7d13d515b9d70d6e;
      (64'h83b071d5ea2aea2a & lut_mask_in) : lut = 64'hff1185759a46b7a0;
      (64'hb8aec52387c687c6 & lut_mask_in) : lut = 64'hd414acb5e363c830;
      (64'h0ddb8426eae8eae8 & lut_mask_in) : lut = 64'hb790c5eece63b7c0;
      (64'had038b8c48794879 & lut_mask_in) : lut = 64'hecaf46cbd1dab4d0;
      (64'h03a5efaf35803580 & lut_mask_in) : lut = 64'hef83162986f45ca5;
      (64'h1abea3a678c878c8 & lut_mask_in) : lut = 64'ha2b3f9c73012e816;
      (64'h62eba8d5ce7bce7b & lut_mask_in) : lut = 64'h130332536e533e55;
      (64'h8ce239d729642964 & lut_mask_in) : lut = 64'h8d1e2660ee4161b9;
      (64'hbcc7b9b783a983a9 & lut_mask_in) : lut = 64'h81b0e2cb03beb7d8;
      (64'h799a64d7d028d028 & lut_mask_in) : lut = 64'h104ff828f311add2;
      (64'h173bb45c106d106d & lut_mask_in) : lut = 64'h801323a63cfd4e89;
      (64'h729170fb7ac87ac8 & lut_mask_in) : lut = 64'h26e8fbfbb457a78b;
      (64'h7a13892b0b160b16 & lut_mask_in) : lut = 64'h27b683d1161b8838;
      (64'hc6b02cd2e725e725 & lut_mask_in) : lut = 64'he665c0440bd48bb8;
      (64'h266bf29d4b644b64 & lut_mask_in) : lut = 64'hb9766375d8116934;
      (64'h4243f771af8caf8c & lut_mask_in) : lut = 64'hdae24e517cff53bc;
      (64'h98604ebd10e710e7 & lut_mask_in) : lut = 64'h9448a6c42573d0bc;
      (64'h02a3323fd23bd23b & lut_mask_in) : lut = 64'h486e515331a14751;
      (64'he5983c643e263e26 & lut_mask_in) : lut = 64'h98f0e56a264a74ef;
      (64'h59d9c15f4f6d4f6d & lut_mask_in) : lut = 64'hcb57867ac3feecb6;
      (64'h9160f34a7e187e18 & lut_mask_in) : lut = 64'hf81d43b8cd023ca2;
      (64'h5e275ede5b2e5b2e & lut_mask_in) : lut = 64'h50073ca8ab257fba;
      (64'hfb8306424ed84ed8 & lut_mask_in) : lut = 64'h22cc30266aaf70cc;
      (64'hf6207f6965a065a0 & lut_mask_in) : lut = 64'h7fef8affeda3d8da;
      (64'h28da610312271227 & lut_mask_in) : lut = 64'h2de5e1f3dfdf184e;
      (64'h035241e8e2f2e2f2 & lut_mask_in) : lut = 64'h64edb8a902c03417;
      (64'hc2e72240af1caf1c & lut_mask_in) : lut = 64'hf46116485c59d257;
      (64'ha6d43ae587398739 & lut_mask_in) : lut = 64'h4147d7a77da1b626;
      (64'hac5ba1a2e71fe71f & lut_mask_in) : lut = 64'ha1e300ae697e9ae5;
      (64'h24bd5437afbeafbe & lut_mask_in) : lut = 64'hfa6dd3b4a8272534;
      (64'h210e48de10351035 & lut_mask_in) : lut = 64'hcb8c1330514b5740;
      (64'h14e185fa26f226f2 & lut_mask_in) : lut = 64'h71025ecb2168db47;
      (64'h5d673fbc06150615 & lut_mask_in) : lut = 64'h776ed9d2c74628d5;
      (64'h37e3f8ad6b3f6b3f & lut_mask_in) : lut = 64'hd6aabeed73c522f6;
      (64'h2e6b39842cbf2cbf & lut_mask_in) : lut = 64'he0b2b59f7e3893fb;
      (64'hd2aed8f5c0b4c0b4 & lut_mask_in) : lut = 64'h2fce6c584c2ead9d;
      (64'h2891b90d7d857d85 & lut_mask_in) : lut = 64'hda4881c91a6381ca;
      (64'hbfc9b13fbf6cbf6c & lut_mask_in) : lut = 64'h82603a1dcbbe439c;
      (64'h0feb97b9544b544b & lut_mask_in) : lut = 64'hbf7f755b256e395d;
      (64'h22d7412d1e191e19 & lut_mask_in) : lut = 64'h37fb1e605e877001;
      (64'heb825e191e3d1e3d & lut_mask_in) : lut = 64'ha1df864a6f2fb37b;
      (64'h081e626d5fff5fff & lut_mask_in) : lut = 64'hc3c1f1a94cdff07f;
      (64'h0e65e4b060816081 & lut_mask_in) : lut = 64'h1ba0a926a4e82bd8;
      (64'he27bcb5fba8fba8f & lut_mask_in) : lut = 64'h6aa8643761a80d8f;
      (64'hc6db43cb03b503b5 & lut_mask_in) : lut = 64'h75bc8f855c5788dc;
      (64'hed2fb47361cb61cb & lut_mask_in) : lut = 64'h74d68705dba2b8ba;
      (64'h5c15cbe97d917d91 & lut_mask_in) : lut = 64'h3e3a9c8e6d967d03;
      (64'h72f96479d3dcd3dc & lut_mask_in) : lut = 64'h09218602dc884ba3;
      (64'h6c4657d114641464 & lut_mask_in) : lut = 64'h82fd32934c4c9808;
      (64'h2f2fc7e7ec89ec89 & lut_mask_in) : lut = 64'h7a155edea613e866;
      (64'hce8622bd1e381e38 & lut_mask_in) : lut = 64'hc8d050c51680d1dd;
      (64'hcf03d094f031f031 & lut_mask_in) : lut = 64'h9e4c297427a6ce9b;
      (64'h2ef7c845322b322b & lut_mask_in) : lut = 64'hf947b1115279904b;
      (64'ha105e030b9e2b9e2 & lut_mask_in) : lut = 64'h94558acc83817e85;
      (64'h00579734db9cdb9c & lut_mask_in) : lut = 64'ha23bbb0e6cdf5a06;
      (64'hf49adcc01a881a88 & lut_mask_in) : lut = 64'ha220d0afefa3be0b;
      (64'h8d4812ddd6c2d6c2 & lut_mask_in) : lut = 64'h8f2b61e3fa20a9d9;
      (64'h94bd62aa90ab90ab & lut_mask_in) : lut = 64'hb86f25779ece3e6d;
      (64'h9814b867cf76cf76 & lut_mask_in) : lut = 64'h486f7c6a8dc86864;
      (64'h5eaf7382682f682f & lut_mask_in) : lut = 64'hf217ca4227f36751;
      (64'h3d8fe7dcef5aef5a & lut_mask_in) : lut = 64'h6b5648b13b83b082;
      (64'h9cb0f9de292f292f & lut_mask_in) : lut = 64'hbd15e9b652cce9b8;
      (64'h2182c070d0e8d0e8 & lut_mask_in) : lut = 64'hb0ad6539195d1ee0;
      (64'h44263abc6e866e86 & lut_mask_in) : lut = 64'h301fea1512cf4d83;
      (64'h446e83703f833f83 & lut_mask_in) : lut = 64'he5246b65a12caa9e;
      (64'h4171a221d49dd49d & lut_mask_in) : lut = 64'h27b5ace1f9db8ada;
      (64'h1422ec2398a198a1 & lut_mask_in) : lut = 64'hcd7a5c5c86d6d3f5;
      (64'h00b01cbea551a551 & lut_mask_in) : lut = 64'h5dec062048ab5394;
      (64'h192740189bb09bb0 & lut_mask_in) : lut = 64'h51af3f811e165176;
      (64'h97f4bbb97ed67ed6 & lut_mask_in) : lut = 64'h6fdf8a5fb07347db;
      (64'h1d5eb2bf4dec4dec & lut_mask_in) : lut = 64'h5837c7486b90312c;
      (64'h55488724c170c170 & lut_mask_in) : lut = 64'h8e307e14c1fb2971;
      (64'ha37004ead41fd41f & lut_mask_in) : lut = 64'h2887dff8ce7e485c;
      (64'h7988dbfb749e749e & lut_mask_in) : lut = 64'h3316f00a2317f5ac;
      (64'hd358ede6702a702a & lut_mask_in) : lut = 64'hf1fdb0791938370c;
      (64'h4c292793e5bee5be & lut_mask_in) : lut = 64'hd10d678e95623a16;
      (64'h7095c5ca1e731e73 & lut_mask_in) : lut = 64'h7665cd68f3245c6c;
      (64'hd91be74e19571957 & lut_mask_in) : lut = 64'h26688dd7e2b786b1;
      (64'h6ab7abe9c7dec7de & lut_mask_in) : lut = 64'h6ece2efb60964f12;
      (64'hb521a556ff5eff5e & lut_mask_in) : lut = 64'h2cdbcc5df089bd77;
      (64'hd7a9df148a318a31 & lut_mask_in) : lut = 64'hb3795843907ab3fc;
      (64'h12acef4ab2e7b2e7 & lut_mask_in) : lut = 64'h1e22e6905ee013e9;
      (64'hf8f74d228faf8faf & lut_mask_in) : lut = 64'h4418f7d6a4463cb9;
      (64'hd1b7a21b62816281 & lut_mask_in) : lut = 64'ha79767f371257dca;
      (64'ha6a2cf6b17b317b3 & lut_mask_in) : lut = 64'hfb5aa178809408cf;
      (64'h1db0fd56edecedec & lut_mask_in) : lut = 64'h9f547086188310a6;
      (64'h23d4592f31513151 & lut_mask_in) : lut = 64'h501f0b75fe854b61;
      (64'ha93735dad75cd75c & lut_mask_in) : lut = 64'h29bd3747baa75a88;
      (64'h8f7a47b4f829f829 & lut_mask_in) : lut = 64'h156f48b395c7a685;
      (64'hbf91671951855185 & lut_mask_in) : lut = 64'hc78b5432baa7d9bb;
      (64'hb76aaff320c420c4 & lut_mask_in) : lut = 64'hd12a53730abe9cdf;
      (64'h1b065df749d349d3 & lut_mask_in) : lut = 64'hcb177b92fc2b51cb;
      (64'h68b75a41e8f1e8f1 & lut_mask_in) : lut = 64'h9e2f8c282857fba5;
      (64'hfb9f5c0f47704770 & lut_mask_in) : lut = 64'h7bb90e3be7c89bbe;
      (64'h134ac6170ab40ab4 & lut_mask_in) : lut = 64'h2f361e4c24838488;
      (64'h15ef9b2ac168c168 & lut_mask_in) : lut = 64'h83228f89a36236db;
      (64'h5fac684ccf1acf1a & lut_mask_in) : lut = 64'h1f5fffa2460146e8;
      (64'h3bd5a00fddc2ddc2 & lut_mask_in) : lut = 64'hacaadb39803b3ad5;
      (64'hf43bfe37f93af93a & lut_mask_in) : lut = 64'h7ccba119475e502b;
      (64'h012b046350475047 & lut_mask_in) : lut = 64'hf53b9e7cafb9bd53;
      (64'he02026b777c177c1 & lut_mask_in) : lut = 64'h204628bb56988162;
      (64'h7fab0bdb3e383e38 & lut_mask_in) : lut = 64'hffb7048d64e9f21d;
      (64'hafc0866ed2cdd2cd & lut_mask_in) : lut = 64'h422ddb20401f9c2c;
      (64'h05c5c2e099809980 & lut_mask_in) : lut = 64'hd41e4c008ed9faeb;
      (64'h48873094be62be62 & lut_mask_in) : lut = 64'hb533ca74e6ddc8fb;
      (64'h9d7b50b853e153e1 & lut_mask_in) : lut = 64'h3173454e74b11d15;
      (64'h16d583e8154b154b & lut_mask_in) : lut = 64'hb09d6a09d2343b0c;
      (64'he1751c06f37df37d & lut_mask_in) : lut = 64'h4154850d8dc109b2;
      (64'hf2003146d2b5d2b5 & lut_mask_in) : lut = 64'hb08d7d27b9d5180b;
      (64'hbc6f31a286f186f1 & lut_mask_in) : lut = 64'ha918dfcf240d295b;
      (64'hdab27d1c4f904f90 & lut_mask_in) : lut = 64'h8fed1937430d06bc;
      (64'h1a0b3ed5a59fa59f & lut_mask_in) : lut = 64'h3637cf7df4b5fc19;
      (64'h48245690874c874c & lut_mask_in) : lut = 64'h99ee8cdbc0d749d3;
      (64'h7905df84c93dc93d & lut_mask_in) : lut = 64'h59a8d616602365eb;
      (64'h07845d5ef3d6f3d6 & lut_mask_in) : lut = 64'h0c6d5debf8e87b1e;
      (64'hc4a6007483eb83eb & lut_mask_in) : lut = 64'h8bf7ccb13f1e72ab;
      (64'h95c107bfd1bad1ba & lut_mask_in) : lut = 64'hc38dba43c9f8d430;
      (64'h860091b335033503 & lut_mask_in) : lut = 64'h014dd2e22d9982f7;
      (64'h08989b0370f070f0 & lut_mask_in) : lut = 64'h11427587f67c4356;
      (64'hb12b32f9c1d5c1d5 & lut_mask_in) : lut = 64'h8177daf2155e8b5f;
      (64'hd265e964c025c025 & lut_mask_in) : lut = 64'h7227b201dba71f48;
      (64'h57ca830fd761d761 & lut_mask_in) : lut = 64'h302cf0400cf2beaf;
      (64'hddabc1da3fe23fe2 & lut_mask_in) : lut = 64'h20c4fd3acef428f4;
      (64'hfe63432f37af37af & lut_mask_in) : lut = 64'h2da22a35134533f8;
      (64'h3743f5db00730073 & lut_mask_in) : lut = 64'h7a435131e5422013;
      (64'h2bf6c7cc9b969b96 & lut_mask_in) : lut = 64'h4fb0c317a81f27e3;
      (64'hcbaee33db665b665 & lut_mask_in) : lut = 64'h7c67eae190511933;
      (64'h93c85177deffdeff & lut_mask_in) : lut = 64'h014322a35a8e6f78;
      (64'h534309c039493949 & lut_mask_in) : lut = 64'hf1bb3b7eb45172c4;
      (64'h7abb4e8e03d503d5 & lut_mask_in) : lut = 64'h00f3c408f2c6b792;
      (64'h8299644fae42ae42 & lut_mask_in) : lut = 64'h12427b70c4dc23c6;
      (64'he16fc64873de73de & lut_mask_in) : lut = 64'h5b615429a2c54e50;
      (64'hef2c66b12ce42ce4 & lut_mask_in) : lut = 64'hf4b43b6f002b42f1;
      (64'h738055ab49d449d4 & lut_mask_in) : lut = 64'h98caf98d6fbd05fa;
      (64'h44ce24ba21a221a2 & lut_mask_in) : lut = 64'hd240b46e46794b05;
      (64'h4bf97b3645b545b5 & lut_mask_in) : lut = 64'he83c418e32bdca57;
      (64'he825edb0a667a667 & lut_mask_in) : lut = 64'hd8c77d769d1b0501;
      (64'h39232909b83ab83a & lut_mask_in) : lut = 64'hff983c6801156187;
      (64'h99426684fda1fda1 & lut_mask_in) : lut = 64'he17642c69609e6f7;
      (64'hbc172230890e890e & lut_mask_in) : lut = 64'hf0b9ce02b6328ce7;
      (64'h86a442eb25e325e3 & lut_mask_in) : lut = 64'h1ee2e3ea3eb99116;
      (64'hd1c78b3b78387838 & lut_mask_in) : lut = 64'hf8e9f609c66c7f07;
      (64'h79a1aa82d6c1d6c1 & lut_mask_in) : lut = 64'h9e4a12e90b9f4832;
      (64'h2fe8389e502f502f & lut_mask_in) : lut = 64'h09bb58a606672c5a;
      (64'h62f3def065f265f2 & lut_mask_in) : lut = 64'h76e235d2e7054cef;
      (64'h40090989015a015a & lut_mask_in) : lut = 64'hb06ca982fb174265;
      (64'h8030ba1bbd37bd37 & lut_mask_in) : lut = 64'h32905e2ab4c6d53d;
      (64'hcff9999894819481 & lut_mask_in) : lut = 64'h98940f7c4b98f6f8;
      (64'h818733d7d566d566 & lut_mask_in) : lut = 64'hfba08c218277e39d;
      (64'h799cccdf590a590a & lut_mask_in) : lut = 64'h647c4abf80780262;
      (64'h43612552aa82aa82 & lut_mask_in) : lut = 64'h36c6d814b93fd327;
      (64'h6a5f25815ae15ae1 & lut_mask_in) : lut = 64'h260e5525d2058c01;
      (64'h60f9654470a770a7 & lut_mask_in) : lut = 64'h65bf82ad29ba96f2;
      (64'hd930ef2e03d103d1 & lut_mask_in) : lut = 64'h8cbe2117134504f7;
      (64'he62c3358b62eb62e & lut_mask_in) : lut = 64'hf6d93794698b8068;
      (64'h62654d71b4eeb4ee & lut_mask_in) : lut = 64'hf93e09eecaf6d67d;
      (64'h214a9570a2b5a2b5 & lut_mask_in) : lut = 64'h4973fe2d8780b295;
      (64'h131d56ed25782578 & lut_mask_in) : lut = 64'hf3bb3ad3efef00b3;
      (64'h570d8181f524f524 & lut_mask_in) : lut = 64'h2e555cbf96013c38;
      (64'h77eae21f2f0b2f0b & lut_mask_in) : lut = 64'h9460a0ac2785cef4;
      (64'hda962e41ae02ae02 & lut_mask_in) : lut = 64'h8c86a79a2ec1dda3;
      (64'h164fb6a90c520c52 & lut_mask_in) : lut = 64'h3fa739c7556cbc7f;
      (64'hc6e91559de4dde4d & lut_mask_in) : lut = 64'h2e7d379de64e2669;
      (64'h37a831acbafabafa & lut_mask_in) : lut = 64'h835de609cee8379f;
      (64'h59907fadb011b011 & lut_mask_in) : lut = 64'he5587b2d2ff815b5;
      (64'haa2b34c95f8d5f8d & lut_mask_in) : lut = 64'h1fbe41bdf7a01289;
      (64'h36c00c4f5f255f25 & lut_mask_in) : lut = 64'ha55ad6b3ae769eaa;
      (64'haf75c386a9e4a9e4 & lut_mask_in) : lut = 64'hf242d7e0d81b2ac4;
      (64'h3fa8d7bbe2b0e2b0 & lut_mask_in) : lut = 64'hcf60fdaeb1a55e91;
      (64'hd37ba9c596349634 & lut_mask_in) : lut = 64'h39b46cd5a64e647a;
      (64'h10a799375d5c5d5c & lut_mask_in) : lut = 64'h8d1fc96ac0c84bdd;
      (64'h37e9f6d967f567f5 & lut_mask_in) : lut = 64'h63a8ae0b58f2bf6c;
      (64'hfec9d1b913161316 & lut_mask_in) : lut = 64'h7efd627e4c935ef5;
      (64'hf47a1e82135d135d & lut_mask_in) : lut = 64'h63293fcf73568738;
      (64'hf019383c633e633e & lut_mask_in) : lut = 64'ha15cd6f18372fc8c;
      (64'h20b2c7ac88038803 & lut_mask_in) : lut = 64'he1ee7cbf7634909a;
      (64'hf675e25f87b487b4 & lut_mask_in) : lut = 64'hfb9114de489082f3;
      (64'hbf3004043aa03aa0 & lut_mask_in) : lut = 64'h4c7d09fb0ebaf193;
      (64'ha6eec7dd05040504 & lut_mask_in) : lut = 64'h09f7be9447a9763b;
      (64'h61493bed707b707b & lut_mask_in) : lut = 64'h89689ffcb2a91aa2;
      (64'h7a5e16deba0bba0b & lut_mask_in) : lut = 64'h38c013457b83e5a0;
      (64'he64002d435523552 & lut_mask_in) : lut = 64'hd06451fd7b908ea3;
      (64'hcb065b47bfccbfcc & lut_mask_in) : lut = 64'hbd5119a5ff541b82;
      (64'hf735452e2ab02ab0 & lut_mask_in) : lut = 64'h21b771e3f8c9e3ab;
      (64'hd953b199933b933b & lut_mask_in) : lut = 64'h75f4646ad11fdc43;
      (64'h9c7afb1e36143614 & lut_mask_in) : lut = 64'h4055a59a30091f7c;
      (64'h7401bd6676ae76ae & lut_mask_in) : lut = 64'h16d099c0ef7b063a;
      (64'h550bc994c4ecc4ec & lut_mask_in) : lut = 64'h462719fd652080e9;
      (64'h25dbae6b80408040 & lut_mask_in) : lut = 64'hee2eb99157a381e6;
      (64'h63004471115e115e & lut_mask_in) : lut = 64'h22fb8ca6441fca05;
      (64'hf6dea1b354585458 & lut_mask_in) : lut = 64'hda0212abf70789c5;
      (64'he826edb46e1a6e1a & lut_mask_in) : lut = 64'ha5d50d52540020ff;
      (64'h4d4f738d9e559e55 & lut_mask_in) : lut = 64'h97c6afa16c56a42c;
      (64'h5d644ed8154d154d & lut_mask_in) : lut = 64'h52762c5f97d151ae;
      (64'h493cc2f881038103 & lut_mask_in) : lut = 64'hd7868053908a401e;
      (64'ha77adaa5fea7fea7 & lut_mask_in) : lut = 64'h05bfbb55f78a5d47;
      (64'h273b788bb584b584 & lut_mask_in) : lut = 64'h195ab11d71a396a9;
      (64'h3c49775010181018 & lut_mask_in) : lut = 64'hc3d0db70db36e01e;
      (64'h65ad99f7a928a928 & lut_mask_in) : lut = 64'h8850b65828cd7633;
      (64'ha13b7082b5ecb5ec & lut_mask_in) : lut = 64'hdad9e8a5019554db;
      (64'hf93efbdfc856c856 & lut_mask_in) : lut = 64'hd85bcbe740bf8ce5;
      (64'ha51b45fc8fcf8fcf & lut_mask_in) : lut = 64'h681f7b9c6540bdc7;
      (64'h2921fa179def9def & lut_mask_in) : lut = 64'hf1c0465aecb04507;
      (64'h5b1d94d1da19da19 & lut_mask_in) : lut = 64'hc16aa5f273ffffbb;
      (64'h32c83b31e056e056 & lut_mask_in) : lut = 64'hdf47ba3c07902004;
      (64'hac17d55c6aa76aa7 & lut_mask_in) : lut = 64'hf1eba30213201b01;
      (64'ha86c9291fe90fe90 & lut_mask_in) : lut = 64'h18755ddc71548336;
      (64'h9651d7ebc068c068 & lut_mask_in) : lut = 64'he028245fe87bc524;
      (64'h1f389baf1a9a1a9a & lut_mask_in) : lut = 64'h239fc0457ddba9d7;
      (64'hb1709c689f699f69 & lut_mask_in) : lut = 64'h5c628ff2ad934ce2;
      (64'he0b164b9dab1dab1 & lut_mask_in) : lut = 64'h5335269eeda19b78;
      (64'h544ecbf5c35dc35d & lut_mask_in) : lut = 64'h60cbe67acce1ec70;
      (64'hf6d6d4062c182c18 & lut_mask_in) : lut = 64'h4c0486cabb295dab;
      (64'h407fa7051d2b1d2b & lut_mask_in) : lut = 64'h1777945bac8690fc;
      (64'ha6eac3e7fe2dfe2d & lut_mask_in) : lut = 64'h98a708f7b121648a;
      (64'hade919306a106a10 & lut_mask_in) : lut = 64'hbf9604cb0fe69f0d;
      (64'h1fb92bea61516151 & lut_mask_in) : lut = 64'h0e750088cb3cb4f3;
      (64'h4be0521210001000 & lut_mask_in) : lut = 64'hea1710f390cf7214;
      (64'h7236ca8e73707370 & lut_mask_in) : lut = 64'hcb2954076b2c5356;
      (64'h86941816ca20ca20 & lut_mask_in) : lut = 64'h4a0e50eeabba6c2f;
      (64'hbd9ef6c73a7c3a7c & lut_mask_in) : lut = 64'hbcaab8a21e6de6c7;
      (64'h4fdb7b23b281b281 & lut_mask_in) : lut = 64'h11a69a7fc464d254;
      (64'heba9e92a630a630a & lut_mask_in) : lut = 64'h04e35913644ec085;
      (64'hf54cd9433f653f65 & lut_mask_in) : lut = 64'hd5ace184d86d7867;
      (64'hd18837c23b433b43 & lut_mask_in) : lut = 64'hc1272d6e7f3046c2;
      (64'h3216021ed96ad96a & lut_mask_in) : lut = 64'hb7cd296dca2c6287;
      (64'h9c3f0a27e710e710 & lut_mask_in) : lut = 64'hb1b275c0d8dc0e50;
      (64'h3bfc4d8ccdcecdce & lut_mask_in) : lut = 64'h3c6ce5c64e653c10;
      (64'h8dd5dc239d109d10 & lut_mask_in) : lut = 64'h698778f6462e9c30;
      (64'hd89c5d27a9d8a9d8 & lut_mask_in) : lut = 64'h14cf161ece3df744;
      (64'hd2304822bd0cbd0c & lut_mask_in) : lut = 64'h469daf42d8605e6f;
      (64'h451ffb5773f173f1 & lut_mask_in) : lut = 64'hb04df7d0b075016d;
      (64'he0d0a392ee56ee56 & lut_mask_in) : lut = 64'h546a973210d39a38;
      (64'heebd18146fa66fa6 & lut_mask_in) : lut = 64'h0e95f97be087f67e;
      (64'h82f15c6b2bfa2bfa & lut_mask_in) : lut = 64'h6a61f46e51eed159;
      (64'h6f2407d945e745e7 & lut_mask_in) : lut = 64'haf1ccdd63b09cf0c;
      (64'h261c82ef77187718 & lut_mask_in) : lut = 64'h0360f6f7a27d2e0e;
      (64'h0beca63df498f498 & lut_mask_in) : lut = 64'hbd49494a60cdb329;
      (64'h108e30975e995e99 & lut_mask_in) : lut = 64'h86642073c258dc33;
      (64'h507e1b0e9b7e9b7e & lut_mask_in) : lut = 64'h1f81560303349297;
      (64'h83b872e288818881 & lut_mask_in) : lut = 64'he37f087329d7bcc1;
      (64'h2ea4a86bffeaffea & lut_mask_in) : lut = 64'hbd04793544173b8f;
      (64'h044f51e693449344 & lut_mask_in) : lut = 64'hfc467d0d0a700748;
      (64'h9dbe8e908e228e22 & lut_mask_in) : lut = 64'h653d7e7522ac33ed;
      (64'h5361c0af81478147 & lut_mask_in) : lut = 64'hb07aaf487ab34465;
      (64'he721273c8a728a72 & lut_mask_in) : lut = 64'h76bf67d7501443b9;
      (64'h4805130761826182 & lut_mask_in) : lut = 64'hcfd7e6a6c26a6bca;
      (64'hb1233290b971b971 & lut_mask_in) : lut = 64'h241c5a05d6a6a4fc;
      (64'h1222cdebbaddbadd & lut_mask_in) : lut = 64'h76bb0543fb01862d;
      (64'h4e162a031abe1abe & lut_mask_in) : lut = 64'ha3b989db4a5ac438;
      (64'h0be8dc92e2bfe2bf & lut_mask_in) : lut = 64'h7f60ad311eb7cb0e;
      (64'h4cc0b422a3baa3ba & lut_mask_in) : lut = 64'h2834ad10517ce1ec;
      (64'h7c688a5f499a499a & lut_mask_in) : lut = 64'hf1dcf749efeebaec;
      (64'hb3e7ce5a553b553b & lut_mask_in) : lut = 64'h548b890bb0d52f36;
      (64'he7d57b12d5b6d5b6 & lut_mask_in) : lut = 64'h30359de525dc563e;
      (64'h30a60adcdc34dc34 & lut_mask_in) : lut = 64'h5d2a18b6af3a1758;
      (64'haa71adc6de9dde9d & lut_mask_in) : lut = 64'h01a9c9363ff8ec33;
      (64'hd29c09f541a941a9 & lut_mask_in) : lut = 64'h3f75365d77443a4c;
      (64'h3c732a83df25df25 & lut_mask_in) : lut = 64'hac0d48fc5c56a20e;
      (64'h260b9e981e211e21 & lut_mask_in) : lut = 64'h0627525b6658a6a8;
      (64'h7f0d2aa431623162 & lut_mask_in) : lut = 64'h21c579fe5feb4c35;
      (64'h5a93468f4e424e42 & lut_mask_in) : lut = 64'hdacc6020d8c87b3c;
      (64'h96f1bfd2dbeddbed & lut_mask_in) : lut = 64'hfbebe46647ffabd1;
      (64'hf79e282acbc7cbc7 & lut_mask_in) : lut = 64'h4b7e86973bdea684;
      (64'hd18b7a62acb6acb6 & lut_mask_in) : lut = 64'h5a6f46549a1a0e99;
      (64'h0f8c57f6e675e675 & lut_mask_in) : lut = 64'hb9e7e70b78d8cd97;
      (64'h46e612251cc21cc2 & lut_mask_in) : lut = 64'h1c37eff2352cdd07;
      (64'h150b6d5538c438c4 & lut_mask_in) : lut = 64'hb1859e5c6b1aa531;
      (64'h0302bf05ea5aea5a & lut_mask_in) : lut = 64'he7bb6b274214ae31;
      (64'h6699cdc1e14ce14c & lut_mask_in) : lut = 64'h61ba32a27ca401be;
      (64'h3738088449294929 & lut_mask_in) : lut = 64'h9dbfb7b440b3452b;
      (64'hc408a0df41df41df & lut_mask_in) : lut = 64'hab5d096869e80b6a;
      (64'h1b23698ac56ac56a & lut_mask_in) : lut = 64'h34f8d8817c26c90d;
      (64'h3d8faaccdc9cdc9c & lut_mask_in) : lut = 64'he2b72a15f8a57d2c;
      (64'h709669f5a4eca4ec & lut_mask_in) : lut = 64'h0987fafd739f892b;
      (64'ha505a957af2daf2d & lut_mask_in) : lut = 64'hb63799f54adf2063;
      (64'h05f60a38e207e207 & lut_mask_in) : lut = 64'hb29216b871116d4f;
      (64'h9f99c0fe5ea25ea2 & lut_mask_in) : lut = 64'h2ef51857a9122dac;
      (64'h59a8e5d610f510f5 & lut_mask_in) : lut = 64'h04f31acef0154d54;
      (64'h0fb108496af66af6 & lut_mask_in) : lut = 64'h1860003ac6f85cd1;
      (64'h19697b604d414d41 & lut_mask_in) : lut = 64'h025ad0a5ccf8525a;
      (64'h21d88171fafffaff & lut_mask_in) : lut = 64'he0341e6e626df185;
      (64'hee367a0db3b8b3b8 & lut_mask_in) : lut = 64'hb008fdfc71183182;
      (64'h55e4f7df01e201e2 & lut_mask_in) : lut = 64'h1523588388d82ba9;
      (64'ha99bc8a0c879c879 & lut_mask_in) : lut = 64'hf4e5e07cffe001df;
      (64'h25f8e6eab40cb40c & lut_mask_in) : lut = 64'h209cafe9f9e3e48d;
      (64'h39101228ac35ac35 & lut_mask_in) : lut = 64'h16809a50f4c870f5;
      (64'h394d5df7dedadeda & lut_mask_in) : lut = 64'h70652514efe3fcad;
      (64'h4cdd0b79dea2dea2 & lut_mask_in) : lut = 64'hb7c2b11c016d4ec7;
      (64'hb34342aa86418641 & lut_mask_in) : lut = 64'h38bd5aefc3a0070c;
      (64'hde8719e02d5c2d5c & lut_mask_in) : lut = 64'h35e1f0d8c5ef921d;
      (64'h83796e97faf7faf7 & lut_mask_in) : lut = 64'hadb4ee1c51d6a292;
      (64'h3b571936a463a463 & lut_mask_in) : lut = 64'h0e4f3c1e335dd9ff;
      (64'h08fd9297649f649f & lut_mask_in) : lut = 64'hadd87d2f111c5942;
      (64'h13494f7737c937c9 & lut_mask_in) : lut = 64'h1ea4fc54603f45ef;
      (64'hecc4d399727e727e & lut_mask_in) : lut = 64'hf7a89fb030625a30;
      (64'hba8544bcde5ade5a & lut_mask_in) : lut = 64'h2b71a4ac1a399880;
      (64'hb62b3bdf08190819 & lut_mask_in) : lut = 64'h25d9ecb01500ca8d;
      (64'h656c01bec612c612 & lut_mask_in) : lut = 64'h7183473aea83acc1;
      (64'h0171888102830283 & lut_mask_in) : lut = 64'hfa0789aa9224acef;
      (64'h867c02430adf0adf & lut_mask_in) : lut = 64'h7c122fe10c8d5892;
      (64'hb2949039beacbeac & lut_mask_in) : lut = 64'h004cf8b08b6224ea;
      (64'he5a2bae047624762 & lut_mask_in) : lut = 64'h01da7e3d03340f52;
      (64'hd54ebca085fa85fa & lut_mask_in) : lut = 64'h74a08c3a34ff1aea;
      (64'h02efe44ff843f843 & lut_mask_in) : lut = 64'hd7b4c3c596a7cdca;
      (64'hcec0ab4e1a321a32 & lut_mask_in) : lut = 64'hfa20531298e6b1d3;
      (64'hf3b16c3cd1d6d1d6 & lut_mask_in) : lut = 64'h8b67fc94824a163f;
      (64'h0e8521bd786f786f & lut_mask_in) : lut = 64'h56e3322d486a4948;
      (64'hd90f6c09ed4eed4e & lut_mask_in) : lut = 64'heacce3e14578949e;
      (64'h2f9221c5dadbdadb & lut_mask_in) : lut = 64'hefddc0fc6be93884;
      (64'h01a5bc666d356d35 & lut_mask_in) : lut = 64'hf90c8cb51a7ff987;
      (64'h7dd1b853ef4bef4b & lut_mask_in) : lut = 64'h6dcafbc948fd5249;
      (64'h8ce0f93e634a634a & lut_mask_in) : lut = 64'hf21942363d8ef002;
      (64'h45587492a1d9a1d9 & lut_mask_in) : lut = 64'h24530f4fb09c9b5b;
      (64'hf5c2f76ce807e807 & lut_mask_in) : lut = 64'hdeada5b8bd7e942f;
      (64'h2a30476825b825b8 & lut_mask_in) : lut = 64'h5769e347792ec8e2;
      (64'ha9d4e4dd8a4f8a4f & lut_mask_in) : lut = 64'hac67553fcecec2a0;
      (64'h0095a90a57d657d6 & lut_mask_in) : lut = 64'h36337869032173e6;
      (64'h2fa86025dc15dc15 & lut_mask_in) : lut = 64'h5f7f713174cde0eb;
      (64'h8b21c2fd09b709b7 & lut_mask_in) : lut = 64'h4ab32615a07b5fe4;
      (64'hefb4465ecfd7cfd7 & lut_mask_in) : lut = 64'h3bb55ca0160b20a4;
      (64'hb52af1ad45804580 & lut_mask_in) : lut = 64'h4d276262b2760350;
      (64'h8f8e45a5db07db07 & lut_mask_in) : lut = 64'hee27227bfce8e20d;
      (64'h431c63b9ded1ded1 & lut_mask_in) : lut = 64'hd237a3ff6c33e49a;
      (64'h98571f6e8a768a76 & lut_mask_in) : lut = 64'h3e1ca7083aa397c9;
      (64'hf382c04888e988e9 & lut_mask_in) : lut = 64'h9b48d6884d25f8cc;
      (64'hb5d3c478863a863a & lut_mask_in) : lut = 64'h1a935799ac3b657f;
      (64'h4a12cb2a6c4c6c4c & lut_mask_in) : lut = 64'h42aa9d9b8231ffb7;
      (64'h9605aa0205720572 & lut_mask_in) : lut = 64'hf293e70c4f1460f8;
      (64'h92d09e018df08df0 & lut_mask_in) : lut = 64'hc46632a8876dc84a;
      (64'hfb251d98c356c356 & lut_mask_in) : lut = 64'h8c5a4f88c64e6f11;
      (64'h2c929e4a7faa7faa & lut_mask_in) : lut = 64'hd11f2969b7ed401b;
      (64'hfdd76fb977ca77ca & lut_mask_in) : lut = 64'h36559813b0f45f7b;
      (64'h715036b89e1b9e1b & lut_mask_in) : lut = 64'h0a78e4c0cb675e38;
      (64'h3fa966640bca0bca & lut_mask_in) : lut = 64'hd9ed244f7d63940f;
      (64'h99347b9d084b084b & lut_mask_in) : lut = 64'ha80647d3fad763c0;
      (64'h717f56437caa7caa & lut_mask_in) : lut = 64'h7cad1b03c25f68be;
      (64'hbe9c4f7d92429242 & lut_mask_in) : lut = 64'hd8dfb86ce6c92dc5;
      (64'hc9ee515165256525 & lut_mask_in) : lut = 64'hd312a9d43e5e55a6;
      (64'h576b785285de85de & lut_mask_in) : lut = 64'h984d38239d224613;
      (64'h229f2242c5c2c5c2 & lut_mask_in) : lut = 64'h71308e45291e2bc7;
      (64'h4158396174007400 & lut_mask_in) : lut = 64'h7343baee8e4a26f8;
      (64'hdfa7449acf13cf13 & lut_mask_in) : lut = 64'h7721f587985c527d;
      (64'h35ab1e1518431843 & lut_mask_in) : lut = 64'hed231480777e999e;
      (64'h9936d1910d890d89 & lut_mask_in) : lut = 64'h9494b511083ce3de;
      (64'h91ce9aeed3b2d3b2 & lut_mask_in) : lut = 64'h7d5308ee15b0a14e;
      (64'h4e19f7a44dbe4dbe & lut_mask_in) : lut = 64'hff0f456d949e6d48;
      (64'h0aa74b3a0aed0aed & lut_mask_in) : lut = 64'hd19e62f567567706;
      (64'h2c36fe1181a481a4 & lut_mask_in) : lut = 64'hca00d27f8c2c91c2;
      (64'h110ecbf449344934 & lut_mask_in) : lut = 64'h8354d99726eeb9e7;
      (64'hdd573e821bfe1bfe & lut_mask_in) : lut = 64'haa8c9ff177ca97c2;
      (64'h11b3ec27fb91fb91 & lut_mask_in) : lut = 64'h4a9ca9af2e401e6f;
      (64'hec1a5e3105070507 & lut_mask_in) : lut = 64'h019dd2785b92c425;
      (64'h3dd211272c642c64 & lut_mask_in) : lut = 64'h506093282b29badd;
      (64'h4b80020f863b863b & lut_mask_in) : lut = 64'hbb60cee74bf5c476;
      (64'h2674cf81ad04ad04 & lut_mask_in) : lut = 64'hcea41bbf679fc570;
      (64'ha08b822216211621 & lut_mask_in) : lut = 64'h57b88dcc8bd22eff;
      (64'hbe3203bedf88df88 & lut_mask_in) : lut = 64'h2713c58e81d1d65d;
      (64'ha70370e489cb89cb & lut_mask_in) : lut = 64'h4202fd85ad27ebb8;
      (64'hb9eb942b7a8f7a8f & lut_mask_in) : lut = 64'h7098f19ce93e0191;
      (64'h839716e281ac81ac & lut_mask_in) : lut = 64'h48e5e2f1bcac3630;
      (64'h6e34bbbc4cc24cc2 & lut_mask_in) : lut = 64'he6ca4ad8582a4629;
      (64'hd4ac194c69ba69ba & lut_mask_in) : lut = 64'h23a529ccfb389730;
      (64'h9cc85150581d581d & lut_mask_in) : lut = 64'hea31fb90ad7d2169;
      (64'h30e83988df20df20 & lut_mask_in) : lut = 64'h6028ea35ab570ead;
      (64'h54c815fcd6c4d6c4 & lut_mask_in) : lut = 64'h173dc30b671516a7;
      (64'hfbcbbeda1a271a27 & lut_mask_in) : lut = 64'hdc914e9f8267dcc6;
      (64'h80b5e1ae324d324d & lut_mask_in) : lut = 64'heb7ae5302a96fb72;
      (64'h2136c9988e2d8e2d & lut_mask_in) : lut = 64'h5231779e16ac779d;
      (64'h169f0f726ca06ca0 & lut_mask_in) : lut = 64'h8f21cce401332e07;
      (64'h6adcd5a1b6d8b6d8 & lut_mask_in) : lut = 64'h99e70efb1d17c1a0;
      (64'hc935179b3bbc3bbc & lut_mask_in) : lut = 64'hbfdc95fb9ee8e556;
      (64'h015b44aaba36ba36 & lut_mask_in) : lut = 64'hd072b3bfbc0439a5;
      (64'hd0b52ce24d7d4d7d & lut_mask_in) : lut = 64'hcf1f6a39e87d255c;
      (64'h80090837822c822c & lut_mask_in) : lut = 64'h1421ea2048e10f76;
      (64'hd38499d217951795 & lut_mask_in) : lut = 64'haed5568e9c44b77d;
      (64'h586247a753495349 & lut_mask_in) : lut = 64'hb67a8dd9515c8f36;
      (64'hf9210718ff9aff9a & lut_mask_in) : lut = 64'h3917a9ab89cb0159;
      (64'h31e51798ffdbffdb & lut_mask_in) : lut = 64'h91c3f3b30a3cc479;
      (64'h0e04d047b635b635 & lut_mask_in) : lut = 64'h963ce3fb3b63533e;
      (64'hd1c64aec66626662 & lut_mask_in) : lut = 64'h9819de035339280c;
      (64'hcccaa458ea4fea4f & lut_mask_in) : lut = 64'hcbaec76d7dcfef21;
      (64'hc3a03ed7118e118e & lut_mask_in) : lut = 64'h29dc6a94255e7985;
      (64'h2f67433cb3fcb3fc & lut_mask_in) : lut = 64'h99c2e441149313ae;
      (64'h35eacb54a56ea56e & lut_mask_in) : lut = 64'h1af130ba6bfb9dbb;
      (64'hb6a5f268f78bf78b & lut_mask_in) : lut = 64'h9ede7efb67141323;
      (64'h2e1013bed24fd24f & lut_mask_in) : lut = 64'h25f7278b3f323a01;
      (64'h0ce680dc7f707f70 & lut_mask_in) : lut = 64'h787e2be712a1087c;
      (64'haf39a46cc0b2c0b2 & lut_mask_in) : lut = 64'h9f97744592cfd9fd;
      (64'hbb88a4f0f3f5f3f5 & lut_mask_in) : lut = 64'h42f8aa3825820de4;
      (64'h22e8b1f85cfb5cfb & lut_mask_in) : lut = 64'hf8b98cb1f7ccd79a;
      (64'h5e754d3377c577c5 & lut_mask_in) : lut = 64'hba9538982d037549;
      (64'h15d7bcb933133313 & lut_mask_in) : lut = 64'h902c34a684c71134;
      (64'h9a67701551d151d1 & lut_mask_in) : lut = 64'h7a2a2f4585b5e208;
      (64'h796f7020a322a322 & lut_mask_in) : lut = 64'ha99b52ee6ca7a007;
      (64'h8b661e6d4b2a4b2a & lut_mask_in) : lut = 64'h89225e2f2dfd0222;
      (64'h7a29535ae095e095 & lut_mask_in) : lut = 64'h6cf55bea6f93571a;
      (64'ha4b1874485f485f4 & lut_mask_in) : lut = 64'hee41eabcd8697c0b;
      (64'h817b0b205e265e26 & lut_mask_in) : lut = 64'hf3638d0ba310bcca;
      (64'h448008363ce43ce4 & lut_mask_in) : lut = 64'h5e0eaad0b7894893;
      (64'hd932027ab310b310 & lut_mask_in) : lut = 64'h89030107a36f92a5;
      (64'h61074d90ffbeffbe & lut_mask_in) : lut = 64'hd673fbafa6e036ef;
      (64'h64c844b733ee33ee & lut_mask_in) : lut = 64'h316e865c8669b8a9;
      (64'h7fe43dc571327132 & lut_mask_in) : lut = 64'hbb85189836168d4a;
      (64'hf6013be0b915b915 & lut_mask_in) : lut = 64'h2d756f602dc7d925;
      (64'h54ed7c01144a144a & lut_mask_in) : lut = 64'h962c769aa87ca995;
      (64'h39362d7c2b2c2b2c & lut_mask_in) : lut = 64'h236bd866f729364c;
      (64'hea3049d78a0e8a0e & lut_mask_in) : lut = 64'h755c23a2fcb612c7;
      (64'h445c2187b732b732 & lut_mask_in) : lut = 64'h929b232dbad5261e;
      (64'h8a101090407c407c & lut_mask_in) : lut = 64'h0c5aceb54a3036bb;
      (64'hf699ef8cc02cc02c & lut_mask_in) : lut = 64'h9bc9f7efa3e4db26;
      (64'h6acbe8b7ac91ac91 & lut_mask_in) : lut = 64'hfcedaead45f83a3c;
      (64'he480352c1dc41dc4 & lut_mask_in) : lut = 64'hf231d062a764a284;
      (64'hda4a81293b233b23 & lut_mask_in) : lut = 64'hbbaa1c7aed0156dd;
      (64'h1d11d51881b481b4 & lut_mask_in) : lut = 64'hbafa393c609e650d;
      (64'hbe8281d45b145b14 & lut_mask_in) : lut = 64'h7256aee5ef978315;
      (64'h90efab46bb75bb75 & lut_mask_in) : lut = 64'h70b5ed3d3ba545a8;
      (64'h5fb4830715951595 & lut_mask_in) : lut = 64'h8caff0f504b03b63;
      (64'h94e34867f7cef7ce & lut_mask_in) : lut = 64'h27e30f86dedfd574;
      (64'h9b03a95720dd20dd & lut_mask_in) : lut = 64'h01b52f7249ccf6b6;
      (64'hfd061ead95eb95eb & lut_mask_in) : lut = 64'hb89e5cf0ad44d1a1;
      (64'h1eddbfeb94fb94fb & lut_mask_in) : lut = 64'h1f00b68290ec74c6;
      (64'hce3e700aec14ec14 & lut_mask_in) : lut = 64'h7df5fcfd2d8a5bb6;
      (64'h9c8c925731933193 & lut_mask_in) : lut = 64'hc32f05925215d38f;
      (64'h22ea556fdd52dd52 & lut_mask_in) : lut = 64'h8b49aeab95e4615a;
      (64'h784ca5be4fc44fc4 & lut_mask_in) : lut = 64'hab65e30a2965eaa9;
      (64'h84e7a7d0cfaecfae & lut_mask_in) : lut = 64'h0a63da7c74796d7a;
      (64'he064f8afbe8abe8a & lut_mask_in) : lut = 64'h2958990d206cdbf2;
      (64'hc65159606dd66dd6 & lut_mask_in) : lut = 64'h8d8d2fa35bd12329;
      (64'h8060529832433243 & lut_mask_in) : lut = 64'hdd07cc7094db4be0;
      (64'h90a029d5eae9eae9 & lut_mask_in) : lut = 64'h8e252704ed0d23c3;
      (64'hec54316195fd95fd & lut_mask_in) : lut = 64'h4d9ec60451af8e1a;
      (64'hc666d34246434643 & lut_mask_in) : lut = 64'h71595dcd3af75da5;
      (64'hf004bcdb160c160c & lut_mask_in) : lut = 64'hee1932669624d420;
      (64'hd3e0cb5785838583 & lut_mask_in) : lut = 64'h01cba01919db2fd8;
      (64'hc20fe87a64b164b1 & lut_mask_in) : lut = 64'h4ed09e5ecf8272a9;
      (64'h519c6220d385d385 & lut_mask_in) : lut = 64'h3ca43f563734ed25;
      (64'hec786fa1ec1aec1a & lut_mask_in) : lut = 64'hfa6904d715a1f126;
      (64'h540a2f9aa944a944 & lut_mask_in) : lut = 64'h6dbf143f2d6c717a;
      (64'h564f3642c73cc73c & lut_mask_in) : lut = 64'hb186d08c33f7828a;
      (64'hfe62028360736073 & lut_mask_in) : lut = 64'hc3ac373a58b20057;
      (64'ha33c8c7636fc36fc & lut_mask_in) : lut = 64'h7110d9498d41c919;
      (64'hcfd3ee92fe98fe98 & lut_mask_in) : lut = 64'heff30e45bbc32dc8;
      (64'h69d25e36e76ce76c & lut_mask_in) : lut = 64'h5a684dcf0a0e7a24;
      (64'h3a9363e0a05ca05c & lut_mask_in) : lut = 64'h83663337662db6f4;
      (64'ha4c4bc1332cb32cb & lut_mask_in) : lut = 64'hc8a3d199dc627b02;
      (64'he2277a08d045d045 & lut_mask_in) : lut = 64'h39e6bb7940079f05;
      (64'h3074332268a568a5 & lut_mask_in) : lut = 64'hf4c4d938ca042e64;
      (64'hfa578c4053e253e2 & lut_mask_in) : lut = 64'h3599c221505b91f0;
      (64'h95c2f43853045304 & lut_mask_in) : lut = 64'h5a76ade01c3000c3;
      (64'hb55d0ab75e085e08 & lut_mask_in) : lut = 64'h1e312182e1a91cf8;
      (64'h7d56605183088308 & lut_mask_in) : lut = 64'h4ec0d1f116adbfc4;
      (64'hf420426c9ed19ed1 & lut_mask_in) : lut = 64'h2365aa6e1f6b6474;
      (64'h3e18e004cdc9cdc9 & lut_mask_in) : lut = 64'h2e5aa3647149cc09;
      (64'hbae73fe857715771 & lut_mask_in) : lut = 64'h2197baf0ab9ca702;
      (64'h17bc5ef4e109e109 & lut_mask_in) : lut = 64'hd141990fac28785f;
      (64'hca3822f440134013 & lut_mask_in) : lut = 64'h38997fa5fb873a9c;
      (64'h4b9cf01eb756b756 & lut_mask_in) : lut = 64'h937f86c7bd751a9b;
      (64'h06318c5c88b788b7 & lut_mask_in) : lut = 64'h787f5076f142b94b;
      (64'h2b930a50c052c052 & lut_mask_in) : lut = 64'h0304dd64af41ea71;
      (64'h139b253262fd62fd & lut_mask_in) : lut = 64'hb35b0bece3705a2f;
      (64'h55ea44d2d251d251 & lut_mask_in) : lut = 64'h787585cd66a7afe6;
      (64'hb2a349b3dad0dad0 & lut_mask_in) : lut = 64'h01d9379cb05b1ff7;
      (64'h9342668ccbefcbef & lut_mask_in) : lut = 64'h4fe244da38ae089f;
      (64'hf257b6c7d84ad84a & lut_mask_in) : lut = 64'h28315d6f60aa313f;
      (64'h7c6ce7ae05100510 & lut_mask_in) : lut = 64'h3d69bbc7167ed288;
      (64'h3579bc77621c621c & lut_mask_in) : lut = 64'h3390c87bb162a311;
      (64'h9d9b438045684568 & lut_mask_in) : lut = 64'h16809d9af66532db;
      (64'h88944ee4e227e227 & lut_mask_in) : lut = 64'hfd799aa90dafd005;
      (64'h85a914c49ed29ed2 & lut_mask_in) : lut = 64'ha10738e260504815;
      (64'h946613bff6fdf6fd & lut_mask_in) : lut = 64'h4ceca0934cc7c83d;
      (64'hf2c1481f6a8b6a8b & lut_mask_in) : lut = 64'h9b357b057ecb6802;
      (64'he6c5df4fe70ae70a & lut_mask_in) : lut = 64'heba5f3723bc0b0f3;
      (64'h7428d83463e763e7 & lut_mask_in) : lut = 64'h6bedf46a13e027bd;
      (64'hcd79999b130b130b & lut_mask_in) : lut = 64'hf881c4b74239c88b;
      (64'hd37703786e016e01 & lut_mask_in) : lut = 64'h955090e87cc53f57;
      (64'h5d8ef4ee394a394a & lut_mask_in) : lut = 64'h917e9be3bc363edf;
      (64'hedad28a73d543d54 & lut_mask_in) : lut = 64'h7bd4c2f122f409f6;
      (64'hae6c9fbe8d598d59 & lut_mask_in) : lut = 64'h779f6de7ad9e35e2;
      (64'hb8cd8918d06cd06c & lut_mask_in) : lut = 64'h286bf543072cb255;
      (64'h7175c50f84508450 & lut_mask_in) : lut = 64'h25109ac5149adb2b;
      (64'h819e6022a480a480 & lut_mask_in) : lut = 64'h8c06cc67ccc9d93f;
      (64'h034ddf38d276d276 & lut_mask_in) : lut = 64'h62430ce48b6aca7b;
      (64'h21ad2bf55bd35bd3 & lut_mask_in) : lut = 64'hd78cf45c24240568;
      (64'h4ea33db9b5abb5ab & lut_mask_in) : lut = 64'hd865df66c727c311;
      (64'h4619e7ec2afb2afb & lut_mask_in) : lut = 64'h256a76cb752b36fa;
      (64'h3e4277f4ceb6ceb6 & lut_mask_in) : lut = 64'h1178a2b871808f6d;
      (64'h72250e85472b472b & lut_mask_in) : lut = 64'h35b78243c43dfefd;
      (64'h0e34853f5bea5bea & lut_mask_in) : lut = 64'ha823fa9223eeb79e;
      (64'hc24daec7835b835b & lut_mask_in) : lut = 64'hd3df2c231a98850d;
      (64'hbca602ccfd44fd44 & lut_mask_in) : lut = 64'he60eb3cb2d1459d6;
      (64'he529be698e238e23 & lut_mask_in) : lut = 64'h47ce1b299b84ff5e;
      (64'hee4e551dbc00bc00 & lut_mask_in) : lut = 64'hd86cfc05fcc944fc;
      (64'h453d9ba0a67aa67a & lut_mask_in) : lut = 64'h5317395e446cae87;
      (64'h3cdb12b5a963a963 & lut_mask_in) : lut = 64'h78114c645e616eb5;
      (64'hb458c445d7aad7aa & lut_mask_in) : lut = 64'h4db7ae498c7e1580;
      (64'hf832636e12771277 & lut_mask_in) : lut = 64'hf5a55f98dae2b8e1;
      (64'hda4036355c3d5c3d & lut_mask_in) : lut = 64'hf102e3783eb5c1b4;
      (64'he554d735ab5aab5a & lut_mask_in) : lut = 64'haed17c451812f422;
      (64'h75381f62ce83ce83 & lut_mask_in) : lut = 64'h8fa0aa1658cbef01;
      (64'h35fc66311b481b48 & lut_mask_in) : lut = 64'h90d90f60b2176868;
      (64'he9c7c0e84ff54ff5 & lut_mask_in) : lut = 64'h372b143faeec3c30;
      (64'he47ffdb683828382 & lut_mask_in) : lut = 64'h26ac25bf17376bf2;
      (64'h47c10e5aea4aea4a & lut_mask_in) : lut = 64'h6ff7cb595dcb083b;
      (64'h4a0bc512cd4dcd4d & lut_mask_in) : lut = 64'hd0df247ac57b38fa;
      (64'h138d15207ef37ef3 & lut_mask_in) : lut = 64'h814a09026bb4cdaa;
      (64'h32a14d1bb9abb9ab & lut_mask_in) : lut = 64'h4dac2bc3cd011217;
      (64'hbf2f5a75922a922a & lut_mask_in) : lut = 64'hce59c581cae2bbdd;
      (64'hcb515b4b3d333d33 & lut_mask_in) : lut = 64'hcab12a99464c4a2e;
      (64'hddad4f76ec94ec94 & lut_mask_in) : lut = 64'h557e6ce9e38595c5;
      (64'h1ae3eaa901460146 & lut_mask_in) : lut = 64'h38041c7c93664a4b;
      (64'hc203b9a7ceedceed & lut_mask_in) : lut = 64'h8df2ecec937583e2;
      (64'h468e3eed5a855a85 & lut_mask_in) : lut = 64'h4f9342a4fe0a3a04;
      (64'ha99b6317d5bad5ba & lut_mask_in) : lut = 64'h21f3b6f31e981d56;
      (64'ha40e1347d6fcd6fc & lut_mask_in) : lut = 64'he5c97b77da89c7c7;
      (64'h61ee1e0e745c745c & lut_mask_in) : lut = 64'h37d87473dee4506f;
      (64'hc0257b9a5fea5fea & lut_mask_in) : lut = 64'hb8290ae635e0d948;
      (64'hb945bc941bd21bd2 & lut_mask_in) : lut = 64'ha39258b8252f903f;
      (64'h9ef4c79397c297c2 & lut_mask_in) : lut = 64'hdd7d0f94f992b49a;
      (64'h4dd44fc250735073 & lut_mask_in) : lut = 64'h45e114cfa5ebc7be;
      (64'h501ad74ee15be15b & lut_mask_in) : lut = 64'h0e7ef25e524bdd23;
      (64'hcc0f8c155b0f5b0f & lut_mask_in) : lut = 64'hcd8d5863873728e7;
      (64'h7545fc0b53bf53bf & lut_mask_in) : lut = 64'hc05fab568c2c272b;
      (64'h4a88bc2d2f372f37 & lut_mask_in) : lut = 64'h6c5a50df603541fd;
      (64'h5b76b774daf2daf2 & lut_mask_in) : lut = 64'heb73937cf49da945;
      (64'h8c96f61b75aa75aa & lut_mask_in) : lut = 64'hcb066ba7b641d541;
      (64'h43492fe427742774 & lut_mask_in) : lut = 64'ha80ba4e40bc4a0f4;
      (64'hbdcf85714e784e78 & lut_mask_in) : lut = 64'h641e71a2b27e9b44;
      (64'h8db41a11ac44ac44 & lut_mask_in) : lut = 64'heebe4138a16a4f98;
      (64'h3d95fe6bdbe6dbe6 & lut_mask_in) : lut = 64'hb6cbfcfa7a152631;
      (64'he8abed2006950695 & lut_mask_in) : lut = 64'h3ecd2a350f86405a;
      (64'hff741b915a665a66 & lut_mask_in) : lut = 64'h9a5794132d914c5c;
      (64'h1008f8e3ffafffaf & lut_mask_in) : lut = 64'hda74a416e2d38a0b;
      (64'he88b22d5497f497f & lut_mask_in) : lut = 64'hf983e21da48f1972;
      (64'h03bc16e067596759 & lut_mask_in) : lut = 64'hcf1c0bae4b69640b;
      (64'h5f554a71392c392c & lut_mask_in) : lut = 64'h7bc4bc0e6721e140;
      (64'h706a94f593789378 & lut_mask_in) : lut = 64'h156667a36f1b70c4;
      (64'hb5a212c2cd63cd63 & lut_mask_in) : lut = 64'h8c5df4a1a52cba10;
      (64'hbe4647dc20a420a4 & lut_mask_in) : lut = 64'h356a62561d1d26b8;
      (64'h072c02aefa14fa14 & lut_mask_in) : lut = 64'h7f5ae8ac7d62f1eb;
      (64'h6b2b228539d039d0 & lut_mask_in) : lut = 64'h91b6f35570d20a41;
      (64'h5fe66670bd10bd10 & lut_mask_in) : lut = 64'h69e0974dcfc11619;
      (64'hb049f8b3a598a598 & lut_mask_in) : lut = 64'h389bf85bc1debf08;
      (64'h4fef6e1dcf50cf50 & lut_mask_in) : lut = 64'h4334a8e4def5db17;
      (64'hca260b068fc98fc9 & lut_mask_in) : lut = 64'h02129c04f97da30a;
      (64'h4e79f54000560056 & lut_mask_in) : lut = 64'h20ac6fa6f0cef527;
      (64'h959a015d1c9a1c9a & lut_mask_in) : lut = 64'h0f7a054df6c8caf2;
      (64'h4e3f2a8400ba00ba & lut_mask_in) : lut = 64'h3e527966671c154c;
      (64'h0bc2a24be4d8e4d8 & lut_mask_in) : lut = 64'hac4932de96fa019b;
      (64'hf622246741594159 & lut_mask_in) : lut = 64'hf3b0cda8463e66d9;
      (64'h3c2ba89a59925992 & lut_mask_in) : lut = 64'hbbf4fa3d5fed3db1;
      (64'h1711d1128aeb8aeb & lut_mask_in) : lut = 64'h4e6ca78234936126;
      (64'h58e1d53c8ae88ae8 & lut_mask_in) : lut = 64'he908272c9a924171;
      (64'h8c032ec5a8c9a8c9 & lut_mask_in) : lut = 64'hccb89400fcb0405a;
      (64'h73fc567a4df74df7 & lut_mask_in) : lut = 64'h8992923be95bdceb;
      (64'hc274ec9fb019b019 & lut_mask_in) : lut = 64'h42b0a0e9fb168183;
      (64'h6eda6caf6f1a6f1a & lut_mask_in) : lut = 64'h30637fd726fcba8f;
      (64'h0b90bd3552d652d6 & lut_mask_in) : lut = 64'h3f4163607ac95b79;
      (64'h8ffccc7296fe96fe & lut_mask_in) : lut = 64'h29b14f927a0afcb3;
      (64'h88885e33226a226a & lut_mask_in) : lut = 64'h575463cdffb3b5e5;
      (64'h4c04864176657665 & lut_mask_in) : lut = 64'h9f47a84aea2ec586;
      (64'hbecbf5f111f311f3 & lut_mask_in) : lut = 64'h6429ae365e090500;
      (64'hb5e7daa9a140a140 & lut_mask_in) : lut = 64'hbf60931e0a2b8bb8;
      (64'hf40944a295de95de & lut_mask_in) : lut = 64'he88fee48cc07acc1;
      (64'hf3bd2be540f040f0 & lut_mask_in) : lut = 64'h7b5b9c6fc97a3625;
      (64'h8a8da80b81348134 & lut_mask_in) : lut = 64'h10dd2c20e94a6d07;
      (64'h28e12cc8b241b241 & lut_mask_in) : lut = 64'hf3bbf77fe016042b;
      (64'h9e0d7bb004240424 & lut_mask_in) : lut = 64'hc2ed4593955277f5;
      (64'h672c5c1c0d670d67 & lut_mask_in) : lut = 64'h3bb8b460acf37d81;
      (64'h868db82122042204 & lut_mask_in) : lut = 64'h3572faacfe20b859;
      (64'h1c680a9250ca50ca & lut_mask_in) : lut = 64'h1f3703f651bb3128;
      (64'ha13381d006760676 & lut_mask_in) : lut = 64'h5395fcb33a104497;
      (64'h5197716735d735d7 & lut_mask_in) : lut = 64'hfa38c9f810f39425;
      (64'h3f2394e4be44be44 & lut_mask_in) : lut = 64'h88f39306f97d1824;
      (64'h6d140bb4932d932d & lut_mask_in) : lut = 64'hb43340ba08695d91;
      (64'hbf7ba4cdabc7abc7 & lut_mask_in) : lut = 64'hddc3d1384dcd407e;
      (64'h7b422d429bb39bb3 & lut_mask_in) : lut = 64'h304a5245d87a4b2a;
      (64'h1f8b8a1736833683 & lut_mask_in) : lut = 64'h4a2bc16adc3f1712;
      (64'h84ed4fd207f607f6 & lut_mask_in) : lut = 64'h71e55f86a13bfb0b;
      (64'h2ab581d2dfa0dfa0 & lut_mask_in) : lut = 64'h3521101eee68f82b;
      (64'h15b60cc394579457 & lut_mask_in) : lut = 64'h7df4a1bc89816c04;
      (64'h0f6d2a83e45ce45c & lut_mask_in) : lut = 64'hdc07f53e274cd8ee;
      (64'h0250633c85848584 & lut_mask_in) : lut = 64'h594fd670ee25e1c7;
      (64'hdfbe5c7cb66eb66e & lut_mask_in) : lut = 64'hbbef955f09cd6d84;
      (64'h9ee74a280ab70ab7 & lut_mask_in) : lut = 64'hf5e6e7e784fc782f;
      (64'h5f98e92c98d498d4 & lut_mask_in) : lut = 64'h1001addfbcf90dfa;
      (64'h25dab3fbc081c081 & lut_mask_in) : lut = 64'hcc83f35ea7134c5d;
      (64'hcc1aba0d8cec8cec & lut_mask_in) : lut = 64'h2478bfdc0039c1cb;
      (64'h28ab74c409250925 & lut_mask_in) : lut = 64'h432f93fa32bb24e4;
      (64'h3617d126726b726b & lut_mask_in) : lut = 64'h14b7d3a94db54340;
      (64'h09f2fed7f5a2f5a2 & lut_mask_in) : lut = 64'he0d16259e2e10fde;
      (64'h8d57ce1f7aec7aec & lut_mask_in) : lut = 64'h11ff6de9a9528be6;
      (64'hde18a7555b985b98 & lut_mask_in) : lut = 64'hfe1cfb7946c425de;
      (64'he91af99d8c968c96 & lut_mask_in) : lut = 64'hdb0c27cc4c8ee0e2;
      (64'hc75d30f3ec82ec82 & lut_mask_in) : lut = 64'h1b34f38e87f9c739;
      (64'hb987221978957895 & lut_mask_in) : lut = 64'h63901cdac8ae50b1;
      (64'h1e4c8f9bbb43bb43 & lut_mask_in) : lut = 64'hf8e8641a4ec1218f;
      (64'h92a25cbd585c585c & lut_mask_in) : lut = 64'h4793a5e49f8cf342;
      (64'hb207171d04330433 & lut_mask_in) : lut = 64'hda4af2360d05ecb7;
      (64'h66a149fcb8dcb8dc & lut_mask_in) : lut = 64'ha4d6346087b0148a;
      (64'ha290fdf0acf3acf3 & lut_mask_in) : lut = 64'hef8c5b158642b4cf;
      (64'hb4d41119a0f5a0f5 & lut_mask_in) : lut = 64'h150b855388a60824;
      (64'h9233ad213ccc3ccc & lut_mask_in) : lut = 64'h872e91e9dd8253ae;
      (64'heb8e123ba309a309 & lut_mask_in) : lut = 64'h54153d2c2890ca7a;
      (64'h762b4aa0d472d472 & lut_mask_in) : lut = 64'hb746208b0dcd0346;
      (64'h14e85cee9b769b76 & lut_mask_in) : lut = 64'h27b727649c15cc09;
      (64'h1b038ecc9f0c9f0c & lut_mask_in) : lut = 64'h39209a0a7f0e66d2;
      (64'h504879fbf9c8f9c8 & lut_mask_in) : lut = 64'hb458060a42e5af3a;
      (64'hde9f00c2f91cf91c & lut_mask_in) : lut = 64'h4dd42e955b7fa78d;
      (64'h3f5ab7609f099f09 & lut_mask_in) : lut = 64'hdab132bf04c94c09;
      (64'h5abe9a7821fb21fb & lut_mask_in) : lut = 64'h34451a2b7c2b7426;
      (64'h24a8d5b8e808e808 & lut_mask_in) : lut = 64'h944d09503635abae;
      (64'h948469f99dca9dca & lut_mask_in) : lut = 64'h7c60f94e3123a4d3;
      (64'h6bebc44077e777e7 & lut_mask_in) : lut = 64'h0851d5793692258c;
      (64'h526a292103b403b4 & lut_mask_in) : lut = 64'h8831a4ff3ac6dc2d;
      (64'h59e070f24daf4daf & lut_mask_in) : lut = 64'hcac75f9bb4f1a08d;
      (64'ha2b0f0463ee73ee7 & lut_mask_in) : lut = 64'h74205431f5480a57;
      (64'h16c01c8bd124d124 & lut_mask_in) : lut = 64'h1d4df5d3472db6ec;
      (64'h9986d5a69bb89bb8 & lut_mask_in) : lut = 64'h8d179501e044617b;
      (64'h88acf1578a098a09 & lut_mask_in) : lut = 64'h1b770893da5cea5a;
      (64'hf450620f6cb86cb8 & lut_mask_in) : lut = 64'h53265507dce5d395;
      (64'h1dfc1819c05ec05e & lut_mask_in) : lut = 64'hfa050c4602689a09;
      (64'hdaf47da16e496e49 & lut_mask_in) : lut = 64'h9b008757de73077d;
      (64'h883d41bfa0caa0ca & lut_mask_in) : lut = 64'h28218475cf3866c4;
      (64'h4203a7b058635863 & lut_mask_in) : lut = 64'h651f133663b1f3fc;
      (64'hf1a60110e4aee4ae & lut_mask_in) : lut = 64'h7d74e20b8a4df37c;
      (64'hda737d6674ef74ef & lut_mask_in) : lut = 64'hb9f805f7ce9ed1ef;
      (64'h0f41572c2a7a2a7a & lut_mask_in) : lut = 64'h331370987e7291a3;
      (64'h558c61dacf64cf64 & lut_mask_in) : lut = 64'hb2b9426b744c672b;
      (64'ha75fbc65d002d002 & lut_mask_in) : lut = 64'h9cb99bfb8cd3687b;
      (64'hd9684b8055895589 & lut_mask_in) : lut = 64'h5bf875dee800648b;
      (64'h935e2649d5a2d5a2 & lut_mask_in) : lut = 64'ha3991633791741ab;
      (64'h18669b1b8ca28ca2 & lut_mask_in) : lut = 64'h35d5d417711bf688;
      (64'h1087384416bf16bf & lut_mask_in) : lut = 64'h9a51acb12b8a469d;
      (64'hbfdc6f7e5a415a41 & lut_mask_in) : lut = 64'h6fa253a1642b3098;
      (64'h8005f90486178617 & lut_mask_in) : lut = 64'h16e4a243a09ceded;
      (64'hd0b5dfe775607560 & lut_mask_in) : lut = 64'h4721890330fa4091;
      (64'hf74502dc16531653 & lut_mask_in) : lut = 64'h354ac27f447eed21;
      (64'h80258f20d12bd12b & lut_mask_in) : lut = 64'h02f658dc198439e5;
      (64'he2f97d1084b484b4 & lut_mask_in) : lut = 64'h1613037d0910580e;
      (64'h4cfe549d852e852e & lut_mask_in) : lut = 64'h71488bc53b27f39e;
      (64'h5cf95d0ab43ab43a & lut_mask_in) : lut = 64'h23321048b079eca2;
      (64'h79bdce3a71a971a9 & lut_mask_in) : lut = 64'he2d12da149508e92;
      (64'hda3114aa11eb11eb & lut_mask_in) : lut = 64'hab1d7d4ee5b7e27a;
      (64'h1f6d3dcf96909690 & lut_mask_in) : lut = 64'h649bc731f55555e0;
      (64'hffc238e701db01db & lut_mask_in) : lut = 64'h55fc528750524b09;
      (64'ha6134f04efedefed & lut_mask_in) : lut = 64'h116622f180544410;
      (64'h69fa64e6dbb9dbb9 & lut_mask_in) : lut = 64'h9e21d4309313dbc9;
      (64'h5d238c9c61216121 & lut_mask_in) : lut = 64'hcb7d77330b24d879;
      (64'h520895bbf193f193 & lut_mask_in) : lut = 64'h9c2fe9d49fe6971b;
      (64'h45fcfc9b0d8a0d8a & lut_mask_in) : lut = 64'h90cc19b445bbd446;
      (64'h7ec047bfe7d1e7d1 & lut_mask_in) : lut = 64'he15a3dc36c87a352;
      (64'h2982f77c781f781f & lut_mask_in) : lut = 64'h520afe54dc6b1c73;
      (64'h7448487e57b157b1 & lut_mask_in) : lut = 64'h0b3d111fa87e2fab;
      (64'h3d2cf8a930363036 & lut_mask_in) : lut = 64'h8b05052b892d4978;
      (64'h4ce1fc61666c666c & lut_mask_in) : lut = 64'hba8fd93f6aa68544;
      (64'hce2b32fe55de55de & lut_mask_in) : lut = 64'h9468eb526de9881e;
      (64'hd30e6b037fb27fb2 & lut_mask_in) : lut = 64'hd974e3f069c4453c;
      (64'h806173b906c906c9 & lut_mask_in) : lut = 64'hd884bb49dc798ef6;
      (64'hf9b2cf0f946d946d & lut_mask_in) : lut = 64'he0a308b25a7255a7;
      (64'h8aa2fe32921a921a & lut_mask_in) : lut = 64'h4138d455e5a5c48c;
      (64'h888aeb891abf1abf & lut_mask_in) : lut = 64'ha74c0c9f4f1945a4;
      (64'hbe23715116d016d0 & lut_mask_in) : lut = 64'h19437512be2508dc;
      (64'hcad5b365c7d1c7d1 & lut_mask_in) : lut = 64'h42e656c7c7297592;
      (64'h064e234a728a728a & lut_mask_in) : lut = 64'hf14d85feb3f015c6;
      (64'h0ccefc7fd0b5d0b5 & lut_mask_in) : lut = 64'hfa720b39d43dc3b9;
      (64'h928f761953025302 & lut_mask_in) : lut = 64'hdef09045729416fd;
      (64'h08b5965abbccbbcc & lut_mask_in) : lut = 64'ha77624005688b66b;
      (64'h36683a115ef95ef9 & lut_mask_in) : lut = 64'hdf99d18624a10268;
      (64'hd0a6bf663c2a3c2a & lut_mask_in) : lut = 64'h1ac934c35b22515f;
      (64'hde82b96d116d116d & lut_mask_in) : lut = 64'h7b306179e6b450c1;
      (64'hc61ac3820c1b0c1b & lut_mask_in) : lut = 64'h8bd2dcc67e06f5fc;
      (64'hf653aa90e0bee0be & lut_mask_in) : lut = 64'h52b64f310aa2feef;
      (64'h4ad03d01dc0adc0a & lut_mask_in) : lut = 64'h74e73e5df916c75e;
      (64'ha4eafda253175317 & lut_mask_in) : lut = 64'h71105e7529602e52;
      (64'h292106952fd72fd7 & lut_mask_in) : lut = 64'hf1b7bd0232565a5f;
      (64'hed9a2694edbfedbf & lut_mask_in) : lut = 64'h09f8315d66212a4d;
      (64'h8a7eadc9b07fb07f & lut_mask_in) : lut = 64'hc4b241185385661e;
      (64'hae56967c99a999a9 & lut_mask_in) : lut = 64'h227b1d662523a1e6;
      (64'h990ff0d2444d444d & lut_mask_in) : lut = 64'h4b541191d0a1ba7a;
      (64'h5ede7c0d5ac35ac3 & lut_mask_in) : lut = 64'h83dc0dc79a966afb;
      (64'hcd1916a513891389 & lut_mask_in) : lut = 64'h178d45b78854297f;
      (64'hcd2350f4bba7bba7 & lut_mask_in) : lut = 64'haf00308d2d80cd34;
      (64'ha9a932b7eb0feb0f & lut_mask_in) : lut = 64'h99fd9ea504dac95d;
      (64'he971cec82f3c2f3c & lut_mask_in) : lut = 64'h1c4bc51d99fd2c64;
      (64'h27ee9f4323152315 & lut_mask_in) : lut = 64'hf47195b669daa2a2;
      (64'h95e859d0749c749c & lut_mask_in) : lut = 64'hbd961cb1405ecdc4;
      (64'heb16cc45aebdaebd & lut_mask_in) : lut = 64'h56726f1b96d02528;
      (64'h39595b9b1b9a1b9a & lut_mask_in) : lut = 64'h4407c1a50d180860;
      (64'h3cfd35cd39bc39bc & lut_mask_in) : lut = 64'hded9007851e624be;
      (64'h41958b9e8e7d8e7d & lut_mask_in) : lut = 64'hd1b56e80cfe7abb0;
      (64'hb00dec9ae61ce61c & lut_mask_in) : lut = 64'hfe105d7a081038d4;
      (64'h3fdafe4c756f756f & lut_mask_in) : lut = 64'h20c3e52265551893;
      (64'hdcc2fe00ce36ce36 & lut_mask_in) : lut = 64'h4c702ded6d756548;
      (64'h569c76766b936b93 & lut_mask_in) : lut = 64'h82c69b5f03e05752;
      (64'h5cb7b7519b619b61 & lut_mask_in) : lut = 64'h7c374d7d94501274;
      (64'haa94296c6b236b23 & lut_mask_in) : lut = 64'h9556f70d9d7ee3e8;
      (64'h331d544ff412f412 & lut_mask_in) : lut = 64'h314942f2e0c7cbb9;
      (64'hdd5fbfdff798f798 & lut_mask_in) : lut = 64'hb02e96beb50daf19;
      (64'hde72aa1b37123712 & lut_mask_in) : lut = 64'h8f4d4418704e3482;
      (64'h613b349dbacbbacb & lut_mask_in) : lut = 64'h3fdd80f4da4f8d45;
      (64'h2889d3a188368836 & lut_mask_in) : lut = 64'h8c81bd62148b7989;
      (64'h462d9f44b1ffb1ff & lut_mask_in) : lut = 64'h9bec5e01080c546a;
      (64'hc567c23b19081908 & lut_mask_in) : lut = 64'h16823c6ce8f5f20f;
      (64'h2bd2e85194609460 & lut_mask_in) : lut = 64'h023fc9c2a55e0bb5;
      (64'h444591d543394339 & lut_mask_in) : lut = 64'h750646fc6b5f1548;
      (64'hf93f145987428742 & lut_mask_in) : lut = 64'hcbfa8fff9f35a90d;
      (64'h759db7f507f507f5 & lut_mask_in) : lut = 64'hb618f4b9cd71cff0;
      (64'hffe0f2b76a386a38 & lut_mask_in) : lut = 64'h4a9d8489bb5bfea3;
      (64'h87e4928d98bb98bb & lut_mask_in) : lut = 64'h49222940b861c174;
      (64'hb12687f02cfe2cfe & lut_mask_in) : lut = 64'hbdcf04a46ec77653;
      (64'hcd6d74d6151c151c & lut_mask_in) : lut = 64'hea95a0507b47ef0d;
      (64'h0158fec415d415d4 & lut_mask_in) : lut = 64'hd5a46c8985d95986;
      (64'h62403bdd40a440a4 & lut_mask_in) : lut = 64'h41f547f510789813;
      (64'h06ca56d6d45cd45c & lut_mask_in) : lut = 64'h39d58922f1d7c8ad;
      (64'haf1dd13bf55cf55c & lut_mask_in) : lut = 64'h3a1e1ac46fecb11b;
      (64'hed7995f075dc75dc & lut_mask_in) : lut = 64'h603c15e47be5cae4;
      (64'hb0901777f77af77a & lut_mask_in) : lut = 64'hb33ae22fc769c944;
      (64'hedfec3aa9bd49bd4 & lut_mask_in) : lut = 64'hb08e8972b19ceb5b;
      (64'h08374d7fadf5adf5 & lut_mask_in) : lut = 64'hb9d6117796955d61;
      (64'hd36ebcfabdeabdea & lut_mask_in) : lut = 64'h15f0763e0938005d;
      (64'he5657b0277797779 & lut_mask_in) : lut = 64'h453c7c287f1979c9;
      (64'hdb577fe6c035c035 & lut_mask_in) : lut = 64'h2e7e72cab38f440d;
      (64'h78a4841c05b105b1 & lut_mask_in) : lut = 64'hcecd23ab6d325a96;
      (64'heae1324fc9ccc9cc & lut_mask_in) : lut = 64'hcd4b0ec10fb06a2a;
      (64'h2b351b38a01fa01f & lut_mask_in) : lut = 64'hdfa25e8e02eece0a;
      (64'h812c118692499249 & lut_mask_in) : lut = 64'h62cbdf22a1aa7f68;
      (64'hb265258a20cd20cd & lut_mask_in) : lut = 64'h22708d85fe68278a;
      (64'ha632e75176257625 & lut_mask_in) : lut = 64'h55e5d0f0ab3742a2;
      (64'h178a35ad7b3e7b3e & lut_mask_in) : lut = 64'h3d4f164ddfe49de3;
      (64'ha4ec2ef02fba2fba & lut_mask_in) : lut = 64'hb5f407657c85adfc;
      (64'hcd56e37796df96df & lut_mask_in) : lut = 64'hb4c5258e1941f11e;
      (64'h19bc22d61a6e1a6e & lut_mask_in) : lut = 64'h79d2a94a43c29d7c;
      (64'h0dd4f9ad54975497 & lut_mask_in) : lut = 64'h8d51a0276143e099;
      (64'h3bcb00668e808e80 & lut_mask_in) : lut = 64'h8b0bef0afe2fb1c1;
      (64'h0f6896759fbf9fbf & lut_mask_in) : lut = 64'ha35c0c688cb68d15;
      (64'hcc8b266dd454d454 & lut_mask_in) : lut = 64'h2a1df9549134e1d5;
      (64'hf0b7e984e7cae7ca & lut_mask_in) : lut = 64'h7db8bb9ddc10a334;
      (64'h91f4d133bb1bbb1b & lut_mask_in) : lut = 64'hcbd3b434708e55d2;
      (64'h2d42b5a016fd16fd & lut_mask_in) : lut = 64'h76fc88c986566eba;
      (64'hf320bac56c646c64 & lut_mask_in) : lut = 64'h4060dc7fca94dbf1;
      (64'h5cc67bf63e4b3e4b & lut_mask_in) : lut = 64'h19333a2fbb6ad4bc;
      (64'h5adf67cfce57ce57 & lut_mask_in) : lut = 64'h4cb58e77df08e6e5;
      (64'h2b6a289cd12ad12a & lut_mask_in) : lut = 64'h5e614bf77b804f97;
      (64'h38096a8050e650e6 & lut_mask_in) : lut = 64'h114482914c7400e3;
      (64'h4855aad458ff58ff & lut_mask_in) : lut = 64'ha4eefdcd88cbdad3;
      (64'h825c1ee104670467 & lut_mask_in) : lut = 64'heeecca232fe2a219;
      (64'h7253dbe420a520a5 & lut_mask_in) : lut = 64'hb195183ab754d1e3;
      (64'h5e59ae744ebb4ebb & lut_mask_in) : lut = 64'hd6d0926b8d542bc4;
      (64'hdf88f741f5e1f5e1 & lut_mask_in) : lut = 64'h664d3f1481f28af3;
      (64'he7115a3b93199319 & lut_mask_in) : lut = 64'h72f1bc4939061039;
      (64'ha5a1383788408840 & lut_mask_in) : lut = 64'h782ba0d2374d0320;
      (64'h8aab6ecd4a874a87 & lut_mask_in) : lut = 64'haa974e6ca21df088;
      (64'hb523d41506740674 & lut_mask_in) : lut = 64'hee9fcd4a4495272e;
      (64'hc93544e7bafebafe & lut_mask_in) : lut = 64'he6ff0fa080e0eb0c;
      (64'h09fba7a480f680f6 & lut_mask_in) : lut = 64'hb062b2677fb64d66;
      (64'h26e42800a274a274 & lut_mask_in) : lut = 64'h7462c7d5704c65ad;
      (64'h70a2cece89c589c5 & lut_mask_in) : lut = 64'h6180bfe5c8facb85;
      (64'h91fc2f2efc2cfc2c & lut_mask_in) : lut = 64'h5a1b70245b804ada;
      (64'hbd0ae0c97d8f7d8f & lut_mask_in) : lut = 64'hfc968b8d950df94a;
      (64'h70d2dc70488e488e & lut_mask_in) : lut = 64'h702f1e8b4ee30672;
      (64'h7695272a85348534 & lut_mask_in) : lut = 64'hb962c7a71aa65980;
      (64'h7856f8f832763276 & lut_mask_in) : lut = 64'h1f54669201268c6f;
      (64'h4dcef32617771777 & lut_mask_in) : lut = 64'hea207118dee00fc7;
      (64'h6885e294b2a0b2a0 & lut_mask_in) : lut = 64'h0a1d360a61b73206;
      (64'h99042ced66d366d3 & lut_mask_in) : lut = 64'h592f8b60bc17fc8d;
      (64'hfd834721cedbcedb & lut_mask_in) : lut = 64'h456fabf475c8c28f;
      (64'hf330964ec077c077 & lut_mask_in) : lut = 64'h6585783a8137ee89;
      (64'hcfa12b7bfbaefbae & lut_mask_in) : lut = 64'h0b76bc6399f5943e;
      (64'h9c59883682e082e0 & lut_mask_in) : lut = 64'hfa758c44439bd4fd;
      (64'h190c2d546ec36ec3 & lut_mask_in) : lut = 64'h5867b9c960cb769d;
      (64'h3fbcf567d431d431 & lut_mask_in) : lut = 64'hd6f18e5eceb46822;
      (64'hef8d80280c620c62 & lut_mask_in) : lut = 64'he549716dd09b3c7f;
      (64'hbcf94258348c348c & lut_mask_in) : lut = 64'h503ae314c7e6a9a5;
      (64'h16303997148f148f & lut_mask_in) : lut = 64'h76f3c51bc086c7d6;
      (64'h123755aad22dd22d & lut_mask_in) : lut = 64'h8d05c24d43b31312;
      (64'hf86b5c78c1e2c1e2 & lut_mask_in) : lut = 64'h7e92c1ad5be7567d;
      (64'hf184b32f02340234 & lut_mask_in) : lut = 64'h93e3222c50a71b64;
      (64'hc6c722a6b508b508 & lut_mask_in) : lut = 64'h7f368de42a2b6d88;
      (64'hbe61e2c8306a306a & lut_mask_in) : lut = 64'hbbd08bfd8e97d3c6;
      (64'h0f7863d4ae52ae52 & lut_mask_in) : lut = 64'hb05092ebeb249d3c;
      (64'h561f6479acceacce & lut_mask_in) : lut = 64'hb85f6b93e6824869;
      (64'h070b8cb920a020a0 & lut_mask_in) : lut = 64'h771b8df71bed9eee;
      (64'h1d43b45cea70ea70 & lut_mask_in) : lut = 64'h98cf37aedaca1a9f;
      (64'h01394a1e76cc76cc & lut_mask_in) : lut = 64'h1c1879a8b5155bc0;
      (64'hda0175ad86498649 & lut_mask_in) : lut = 64'ha4c461fef3d28f40;
      (64'h794c56c452145214 & lut_mask_in) : lut = 64'h2175400942f2ac90;
      (64'h4429a191c2b2c2b2 & lut_mask_in) : lut = 64'h776e07d990fdf08c;
      (64'h6a0ad95d4b4d4b4d & lut_mask_in) : lut = 64'hb9b4206c3596c7ef;
      (64'h3465f6e1bd42bd42 & lut_mask_in) : lut = 64'heb53f49a2d83dac2;
      (64'h7ed6b0aa4ff24ff2 & lut_mask_in) : lut = 64'hdf2e078d9cfe2054;
      (64'h7b2c51d5ace9ace9 & lut_mask_in) : lut = 64'h0f89641a88489e63;
      (64'h6119f3362a712a71 & lut_mask_in) : lut = 64'h99fb92b4b247f1e0;
      (64'hab45303b6d566d56 & lut_mask_in) : lut = 64'hc67b3c1252c558a3;
      (64'h3255bf1565c765c7 & lut_mask_in) : lut = 64'hf0b425dd7dbd83a3;
      (64'hb8bbe87e178d178d & lut_mask_in) : lut = 64'h8b6bb4a06d381e07;
      (64'h5b9c334e4a5a4a5a & lut_mask_in) : lut = 64'h3ee4c472d49d647f;
      (64'hb717f0e262626262 & lut_mask_in) : lut = 64'h8c4ca5b62c90641e;
      (64'hb245f8a315001500 & lut_mask_in) : lut = 64'h0e1529723733ed06;
      (64'hb65eb13becf0ecf0 & lut_mask_in) : lut = 64'hb3c8026abc86ed5a;
      (64'hdfaa3184b8bbb8bb & lut_mask_in) : lut = 64'hb19ef3a408be4cb1;
      (64'hd5341712368c368c & lut_mask_in) : lut = 64'h600b9d8017b58820;
      (64'h50a68edd2fa42fa4 & lut_mask_in) : lut = 64'h8a60ff0c65b7d7b0;
      (64'heb47bd83cdb2cdb2 & lut_mask_in) : lut = 64'haa76aef257e59399;
      (64'h36eb5ed981428142 & lut_mask_in) : lut = 64'h6576d8c47240bf87;
      (64'hb9194b2634b334b3 & lut_mask_in) : lut = 64'h2ff28432b1e2548b;
      (64'h1017e5f0faf9faf9 & lut_mask_in) : lut = 64'h4842922b16cb7946;
      (64'hf24403421fe41fe4 & lut_mask_in) : lut = 64'h86ad7d553a8e8e9a;
      (64'h1740c9abc6e5c6e5 & lut_mask_in) : lut = 64'hcf1b7e1d86369d0c;
      (64'h6f733199ff2dff2d & lut_mask_in) : lut = 64'h9bc7f42099902127;
      (64'h320c4692046f046f & lut_mask_in) : lut = 64'hd70a5cd12d42d828;
      (64'h0cc6ef173d483d48 & lut_mask_in) : lut = 64'h19365fd6e47bdb23;
      (64'hf7634f5f552f552f & lut_mask_in) : lut = 64'hba00a9a9d1a1be1e;
      (64'ha35b631fbeb8beb8 & lut_mask_in) : lut = 64'h6f6feecf8c6fac1c;
      (64'hecd6111e447e447e & lut_mask_in) : lut = 64'hcb034570ed9ee2a9;
      (64'ha4185086e92ae92a & lut_mask_in) : lut = 64'hc5c78e4efa3436ba;
      (64'hd462b48604dd04dd & lut_mask_in) : lut = 64'hbcc854ce86689142;
      (64'h3f4a19697f567f56 & lut_mask_in) : lut = 64'hb14e7e9a798a164a;
      (64'h4451843fe822e822 & lut_mask_in) : lut = 64'h122c5694ef2c4ece;
      (64'hba272a102aa72aa7 & lut_mask_in) : lut = 64'h4f8a0f82404f741d;
      (64'h9654145f3b1e3b1e & lut_mask_in) : lut = 64'h14fbc0e18c9976bd;
      (64'he218a0fb5af25af2 & lut_mask_in) : lut = 64'h408b4386bd2ebec9;
      (64'h479e9e5ec78bc78b & lut_mask_in) : lut = 64'h840674802f39e64a;
      (64'h40acbefa96a596a5 & lut_mask_in) : lut = 64'h8b86866de41af439;
      (64'h2691467a64ea64ea & lut_mask_in) : lut = 64'h68a9c29b4b4900c0;
      (64'h331e6d5d514b514b & lut_mask_in) : lut = 64'h99519f51ba3f1d58;
      (64'h4311afcf4a714a71 & lut_mask_in) : lut = 64'h13a81fd9a7e2481a;
      (64'he4558a0379cc79cc & lut_mask_in) : lut = 64'h8bb04b02e80fbbba;
      (64'h0100d4d95ccf5ccf & lut_mask_in) : lut = 64'h5ea9e1e0016ae7cb;
      (64'h2422bc30318c318c & lut_mask_in) : lut = 64'h351663b1289d5059;
      (64'hc7696f990b500b50 & lut_mask_in) : lut = 64'h5038b3c1fac5cce5;
      (64'h0891bc15ce4fce4f & lut_mask_in) : lut = 64'hfc41196012bca40c;
      (64'h4514458dd052d052 & lut_mask_in) : lut = 64'h3b4da7a45cd83aff;
      (64'h3c2f5e3ad9f9d9f9 & lut_mask_in) : lut = 64'h3fce4648d1f14985;
      (64'hada4028990859085 & lut_mask_in) : lut = 64'h505c47da20111d98;
      (64'hd9a3db4d429e429e & lut_mask_in) : lut = 64'h1d03b0c810b46116;
      (64'h9c13bf6dc367c367 & lut_mask_in) : lut = 64'hd42b6eea30a4b8cf;
      (64'h7b606127c335c335 & lut_mask_in) : lut = 64'hcf0011e8a4901177;
      (64'h1d0e0de80b4d0b4d & lut_mask_in) : lut = 64'h20794b8190e38da2;
      (64'h78afe813ee46ee46 & lut_mask_in) : lut = 64'h337f69b61495526b;
      (64'h6fefe8bf63cb63cb & lut_mask_in) : lut = 64'h9aecc9011301b584;
      (64'hac2d3382d1e7d1e7 & lut_mask_in) : lut = 64'h6f2d444a3531c3bf;
      (64'hfae81a69c3f3c3f3 & lut_mask_in) : lut = 64'h7161166903eed0df;
      (64'h4b43d39ec2b1c2b1 & lut_mask_in) : lut = 64'hab6c807d846a2da8;
      (64'h929754e9f74ef74e & lut_mask_in) : lut = 64'hdf6503af2d832716;
      (64'h4bdd603147d547d5 & lut_mask_in) : lut = 64'h01f516588006bb86;
      (64'hfad9b45412031203 & lut_mask_in) : lut = 64'h40193c79a8f4daf7;
      (64'he7284d64af9baf9b & lut_mask_in) : lut = 64'ha7fa28c5a20903dc;
      (64'h52093017f703f703 & lut_mask_in) : lut = 64'h70f87c96c9d3fc05;
      (64'h9739dfcb004a004a & lut_mask_in) : lut = 64'h3e2138f4a6ce534c;
      (64'hf085212025682568 & lut_mask_in) : lut = 64'h4a38f184b7a9de9b;
      (64'he58dbf6e0be50be5 & lut_mask_in) : lut = 64'h006e827181059b72;
      (64'hbfc8450e25af25af & lut_mask_in) : lut = 64'hfaf310027adc12f0;
      (64'h1b0a9c6641084108 & lut_mask_in) : lut = 64'h302efd792a1d6a90;
      (64'h793d38de86428642 & lut_mask_in) : lut = 64'hbdd86db98b26a098;
      (64'hea65ce866ed86ed8 & lut_mask_in) : lut = 64'h8cb1f48db3e2c4a3;
      (64'hde4ef6c029522952 & lut_mask_in) : lut = 64'hc3e6eed0257bda74;
      (64'hbbfc6fdbd8b3d8b3 & lut_mask_in) : lut = 64'h199627125453a85c;
      (64'h6b3be4aee9fae9fa & lut_mask_in) : lut = 64'h9c111c7ea86fff33;
      (64'haa4d323a2eab2eab & lut_mask_in) : lut = 64'hc641df14d73cab0c;
      (64'h9ef508c8e8c7e8c7 & lut_mask_in) : lut = 64'h6578d6168d550d13;
      (64'h529ec7ad798c798c & lut_mask_in) : lut = 64'h6066219ba2993934;
      (64'h3870e8c60bc90bc9 & lut_mask_in) : lut = 64'h1663c253fdc57669;
      (64'hbdc7d535e5bfe5bf & lut_mask_in) : lut = 64'hffc71bc036ed6958;
      (64'h9a6f9aa8832e832e & lut_mask_in) : lut = 64'h28aebf3432080966;
      (64'h2aa6d9c56ca36ca3 & lut_mask_in) : lut = 64'h68a1fa47476f1d85;
      (64'hda3b5b48597a597a & lut_mask_in) : lut = 64'he8fbcbc849425904;
      (64'hfcbcf3958cda8cda & lut_mask_in) : lut = 64'h876bd44a26f9cb2d;
      (64'h0b808b6a7a6c7a6c & lut_mask_in) : lut = 64'hd03d497989883a68;
      (64'h5a4467084f534f53 & lut_mask_in) : lut = 64'hfebb90a37d1b6384;
      (64'h0380d288aa89aa89 & lut_mask_in) : lut = 64'h1bb5310cdb66e306;
      (64'hc1ca1f7313f613f6 & lut_mask_in) : lut = 64'h66424f49269ad311;
      (64'h3df2a69f7bee7bee & lut_mask_in) : lut = 64'hb56047b05337e817;
      (64'ha811d76a86cf86cf & lut_mask_in) : lut = 64'h9cce299fa3fc01af;
      (64'h8f6dac8d89c789c7 & lut_mask_in) : lut = 64'h5260944de4d176dd;
      (64'h5e6732506a016a01 & lut_mask_in) : lut = 64'ha0c95d978230c085;
      (64'hb6dd12f5801d801d & lut_mask_in) : lut = 64'h3848d3b9901a772e;
      (64'h22ae18d804c404c4 & lut_mask_in) : lut = 64'h3031dae52d09e419;
      (64'h0f53043006660666 & lut_mask_in) : lut = 64'hf0532e3ed14d3606;
      (64'hc933f102521d521d & lut_mask_in) : lut = 64'h7144212e45bf7259;
      (64'h47dd287d07cd07cd & lut_mask_in) : lut = 64'hfc20d7f0a6d8318b;
      (64'hf390d73161f761f7 & lut_mask_in) : lut = 64'hb9d21760b6058d45;
      (64'had9bc168c057c057 & lut_mask_in) : lut = 64'h21e1245c0216af9b;
      (64'h48d576e3bce7bce7 & lut_mask_in) : lut = 64'h4fdb3277964ba910;
      (64'he9d8d42df3c4f3c4 & lut_mask_in) : lut = 64'h94fb96e57c588418;
      (64'ha0501482de86de86 & lut_mask_in) : lut = 64'h57360dd9df0afadd;
      (64'hafb3ca1733573357 & lut_mask_in) : lut = 64'he89458adb0441e7d;
      (64'h0efb66f7a425a425 & lut_mask_in) : lut = 64'h20ae74ad45adae9b;
      (64'h1755b4608ad18ad1 & lut_mask_in) : lut = 64'h68292cd1fa33dc8a;
      (64'hd4dd761eaeebaeeb & lut_mask_in) : lut = 64'h89bd3bfd68b02dde;
      (64'hf5d5e50df180f180 & lut_mask_in) : lut = 64'h7b9b61fab683a49a;
      (64'h1d672e2b16511651 & lut_mask_in) : lut = 64'ha95119765b1e8567;
      (64'hbd9321bb48984898 & lut_mask_in) : lut = 64'h029f45a3127e0730;
      (64'h32c7407efb63fb63 & lut_mask_in) : lut = 64'h0cbc5cca046cc462;
      (64'h5ad930eae685e685 & lut_mask_in) : lut = 64'hd4a9561a849c7911;
      (64'ha176b8b54cba4cba & lut_mask_in) : lut = 64'hba3d3ecb40ad7b42;
      (64'h80c027bb47764776 & lut_mask_in) : lut = 64'ha38b00e8cfc2df34;
      (64'hadad2c22b2a2b2a2 & lut_mask_in) : lut = 64'h8061a512e0865fe1;
      (64'h0a4376e2d60ad60a & lut_mask_in) : lut = 64'h861d031dc9d9dde8;
      (64'hc1d3f3cf56d056d0 & lut_mask_in) : lut = 64'h321110a2bcff3ff0;
      (64'h68d039eaa5cca5cc & lut_mask_in) : lut = 64'h043d0bf8515e53d7;
      (64'hffbc61fc317c317c & lut_mask_in) : lut = 64'hc1c61f1104e0b3ee;
      (64'h1cdacd09e348e348 & lut_mask_in) : lut = 64'he23d38724cf43927;
      (64'hae923938a35da35d & lut_mask_in) : lut = 64'h4e42e7e0d5322dcc;
      (64'h296308e53a7e3a7e & lut_mask_in) : lut = 64'hc2bc12af4d6c3c71;
      (64'hffa6d4f426632663 & lut_mask_in) : lut = 64'h298879ac707a17f7;
      (64'ha7c2a95344fb44fb & lut_mask_in) : lut = 64'h341f03a07d92d44e;
      (64'h412610e9f2c2f2c2 & lut_mask_in) : lut = 64'h59b65d259ef22cba;
      (64'hc974e377a348a348 & lut_mask_in) : lut = 64'h34074862bc4c058a;
      (64'hed95cb0d0a6f0a6f & lut_mask_in) : lut = 64'h3fb439f9c9cbf9b0;
      (64'ha4a758ac10621062 & lut_mask_in) : lut = 64'hdd51110ec573e067;
      (64'h2c8e151dc53bc53b & lut_mask_in) : lut = 64'h1b3df7dee7b42772;
      (64'h305266dcca80ca80 & lut_mask_in) : lut = 64'h6e6fc0e6525a5cf6;
      (64'h98e43e23cf19cf19 & lut_mask_in) : lut = 64'ha347fcdbeeecbe0b;
      (64'he302cb5381958195 & lut_mask_in) : lut = 64'hbacfb4df3aabb6c8;
      (64'h0de5a27e72317231 & lut_mask_in) : lut = 64'hb028d6b3cbf354e6;
      (64'haa3525a5ef64ef64 & lut_mask_in) : lut = 64'ha86eb0ae0ed0aacf;
      (64'hb1b6f5cac0e6c0e6 & lut_mask_in) : lut = 64'h34c73414ebaf2b0f;
      (64'h250b1c4d631a631a & lut_mask_in) : lut = 64'hfc6bf103288310cd;
      (64'h9121142543d743d7 & lut_mask_in) : lut = 64'hede6a17c1aa60fc4;
      (64'h2f60b0efe4bee4be & lut_mask_in) : lut = 64'hbfe13363d4fd552c;
      (64'h677d5a6f9e029e02 & lut_mask_in) : lut = 64'h50db8d4bfd1d58d8;
      (64'h9e9e70e09a0f9a0f & lut_mask_in) : lut = 64'hb1e42498bb33ccb5;
      (64'h93da11538df78df7 & lut_mask_in) : lut = 64'h5aec10afeb64fb42;
      (64'hd58458c08db08db0 & lut_mask_in) : lut = 64'h66090f54c77df8e6;
      (64'hc03fdb8b22aa22aa & lut_mask_in) : lut = 64'hc6ddb476a48b9266;
      (64'h1c00e85cc949c949 & lut_mask_in) : lut = 64'h9db90e2404b97d01;
      (64'hf1d61a6d174a174a & lut_mask_in) : lut = 64'h57506c4d97e130cb;
      (64'h4ec6739924342434 & lut_mask_in) : lut = 64'h6216ba55671ddc41;
      (64'he58ecd6de335e335 & lut_mask_in) : lut = 64'hadb0ea2b0e97fe11;
      (64'h5bb42382ca2cca2c & lut_mask_in) : lut = 64'h6f1b63e58f1bb43e;
      (64'hd17c59a6184a184a & lut_mask_in) : lut = 64'h17537a8edf783149;
      (64'h64ca8980acdeacde & lut_mask_in) : lut = 64'h116aec5aa6f41ccc;
      (64'hdc5a6a4158eb58eb & lut_mask_in) : lut = 64'hbfaea6b130e3cb77;
      (64'hdf2f48c2c698c698 & lut_mask_in) : lut = 64'h104364e50eeeaa4e;
      (64'h1453dc064c384c38 & lut_mask_in) : lut = 64'hccccfeab5dc864ac;
      (64'h8251a42c16d516d5 & lut_mask_in) : lut = 64'h5aaa289956bfc981;
      (64'hb8328532165d165d & lut_mask_in) : lut = 64'haff84701e20bff86;
      (64'h15dec4795d3c5d3c & lut_mask_in) : lut = 64'hd58731e55e97cab9;
      (64'h6b89d23847e047e0 & lut_mask_in) : lut = 64'hd0e40de742d60ed6;
      (64'hbda86845ce54ce54 & lut_mask_in) : lut = 64'h2a189c6a0bbca0a2;
      (64'hfc73a331242f242f & lut_mask_in) : lut = 64'hf39855a922feee8f;
      (64'hd64c84f8bcedbced & lut_mask_in) : lut = 64'he4b791ef34214aaf;
      (64'h503de402a6a4a6a4 & lut_mask_in) : lut = 64'ha35b6bb2aa48f9c3;
      (64'h276aac1b8a6f8a6f & lut_mask_in) : lut = 64'h44ad77f40f31aa81;
      (64'he440be889a409a40 & lut_mask_in) : lut = 64'h152e29fefd2b3bbd;
      (64'hdfa7b88b073d073d & lut_mask_in) : lut = 64'hce79b1142ef8653f;
      (64'h53136acb44f944f9 & lut_mask_in) : lut = 64'h74b65513ad57142d;
      (64'he4dc8c6f6e7a6e7a & lut_mask_in) : lut = 64'h29ce44c2bb1837f8;
      (64'ha5ce93ae1e521e52 & lut_mask_in) : lut = 64'hbe11f4c1edb88d03;
      (64'hfb628e3fb5e8b5e8 & lut_mask_in) : lut = 64'ha3bb56a536f61664;
      (64'h4a054bbc9b399b39 & lut_mask_in) : lut = 64'h3aa4bbe3dd29cc83;
      (64'h6e04ed58e10ee10e & lut_mask_in) : lut = 64'h747de7c2d1a5f6db;
      (64'haf59d26072db72db & lut_mask_in) : lut = 64'h122804b5d29ffeda;
      (64'h60a13d73c843c843 & lut_mask_in) : lut = 64'hab3150bd9682f9ea;
      (64'h059a345ad22bd22b & lut_mask_in) : lut = 64'h0c19ecd23006eab9;
      (64'hfc6f488c426b426b & lut_mask_in) : lut = 64'h1c9add22349f0878;
      (64'h585eff42b4c0b4c0 & lut_mask_in) : lut = 64'hd3997dd3b360a416;
      (64'h049220eada27da27 & lut_mask_in) : lut = 64'h5694d5435e921596;
      (64'h162834b4538e538e & lut_mask_in) : lut = 64'h9a6bf637d477d44c;
      (64'ha25513df8fe38fe3 & lut_mask_in) : lut = 64'h600cd2f3f61094db;
      (64'h71d0f051b5e6b5e6 & lut_mask_in) : lut = 64'hef2f53d599303db2;
      (64'h93e70996322d322d & lut_mask_in) : lut = 64'h98fe9ba1bd913ba8;
      (64'hd6295b1d38aa38aa & lut_mask_in) : lut = 64'hd804395497e82cf1;
      (64'hff0f03a34e574e57 & lut_mask_in) : lut = 64'h8c80ede501a043fa;
      (64'h67d04d4a4c164c16 & lut_mask_in) : lut = 64'he4db32185c7dbcec;
      (64'h056eeda14d4d4d4d & lut_mask_in) : lut = 64'h2ac53fa0f33d8879;
      (64'ha73df5d902a602a6 & lut_mask_in) : lut = 64'h0999b609f66aa9b6;
      (64'h6aa11e491c1b1c1b & lut_mask_in) : lut = 64'ha5e04c461d28a4fd;
      (64'haec429424bd34bd3 & lut_mask_in) : lut = 64'h9568f2e4870feab6;
      (64'h206bf11a22f322f3 & lut_mask_in) : lut = 64'h02082a67cabc8c4b;
      (64'h76e88a86adc8adc8 & lut_mask_in) : lut = 64'h3f1aebf5e670b337;
      (64'hfa12ec1350285028 & lut_mask_in) : lut = 64'h7e57d39fc700df89;
      (64'heb599a4bad1bad1b & lut_mask_in) : lut = 64'hed967a28099e5410;
      (64'h290c2139e096e096 & lut_mask_in) : lut = 64'hed486072dfe51338;
      (64'h73751d29a7dba7db & lut_mask_in) : lut = 64'hc74af6434a414396;
      (64'h0c23ee6c400e400e & lut_mask_in) : lut = 64'h14e7d9ad9ef4d1db;
      (64'h2f96898f97539753 & lut_mask_in) : lut = 64'h0a2a574324ce2b56;
      (64'hc3d77616fa1cfa1c & lut_mask_in) : lut = 64'h1410e0a71ce48c06;
      (64'h28a0411a7c777c77 & lut_mask_in) : lut = 64'h719c443340862aa3;
      (64'h882fec586e226e22 & lut_mask_in) : lut = 64'h5d5578a72f78ff51;
      (64'h85987ac687fb87fb & lut_mask_in) : lut = 64'hd9bcbea7d2b6cd9c;
      (64'hc10b023078c278c2 & lut_mask_in) : lut = 64'h54e1a34d54e5e972;
      (64'h8307b912220f220f & lut_mask_in) : lut = 64'h8fc8a9eba4686a7a;
      (64'hd868c5910ab50ab5 & lut_mask_in) : lut = 64'hd6ca206dc4ac9668;
      (64'h152ea14629532953 & lut_mask_in) : lut = 64'he9b9ce11e47d8982;
      (64'h854b72b3478a478a & lut_mask_in) : lut = 64'hd3a2ea984be2ff6c;
      (64'ha31d3cd0d8f5d8f5 & lut_mask_in) : lut = 64'h7d35273e4774ce5d;
      (64'h70d05d9bc7a9c7a9 & lut_mask_in) : lut = 64'h409da66d759582d5;
      (64'hd0b823f15a155a15 & lut_mask_in) : lut = 64'hd0291ea4cd4ff115;
      (64'h7d3a566a4e5f4e5f & lut_mask_in) : lut = 64'h964473d0ed8f9aa1;
      (64'h9a3579c17fed7fed & lut_mask_in) : lut = 64'h20d85ee1efeb1aa7;
      (64'h1ac16ba1aa92aa92 & lut_mask_in) : lut = 64'h72eff20ae743a56e;
      (64'hafb7c30175cb75cb & lut_mask_in) : lut = 64'h5b65bead2eec19d2;
      (64'hf4ab52a16e0f6e0f & lut_mask_in) : lut = 64'hcf016f4f194e198f;
      (64'h3d365b0fa6f3a6f3 & lut_mask_in) : lut = 64'h9696901dce7da5bb;
      (64'h83dc741ea178a178 & lut_mask_in) : lut = 64'h5e0ded6c4cbcfd18;
      (64'hb49be449f988f988 & lut_mask_in) : lut = 64'h0a0bbc093d555b32;
      (64'h910c633e6bf76bf7 & lut_mask_in) : lut = 64'hc09cfd87c3bee5a5;
      (64'h6d32739d454e454e & lut_mask_in) : lut = 64'h306af98b790b1ba3;
      (64'h41008d0426ed26ed & lut_mask_in) : lut = 64'hfc26ce9a3bb874ad;
      (64'habd45852cf72cf72 & lut_mask_in) : lut = 64'hefbebda24623077f;
      (64'hc4fddc1c67d967d9 & lut_mask_in) : lut = 64'h6cd072046a56c21e;
      (64'hdfb6f275dbdbdbdb & lut_mask_in) : lut = 64'h168d3762ad53450e;
      (64'h988184d442a642a6 & lut_mask_in) : lut = 64'hce85091eaeff5707;
      (64'hfbcbaa1ba8d6a8d6 & lut_mask_in) : lut = 64'h00621d4eca34d6cf;
      (64'h713b4cfca89ba89b & lut_mask_in) : lut = 64'h6786f35981d9e223;
      (64'h4ecab7e1640e640e & lut_mask_in) : lut = 64'hdfb6422e2200da3a;
      (64'h29c560a1e531e531 & lut_mask_in) : lut = 64'h599786f1f2d15e35;
      (64'h93dadcaff729f729 & lut_mask_in) : lut = 64'h3b022fe4eb74df11;
      (64'ha3f03f02c8c9c8c9 & lut_mask_in) : lut = 64'h666f0038cb82f5de;
      (64'h86163763107a107a & lut_mask_in) : lut = 64'hd5ef648e24dd3a3f;
      (64'hc7cf7e58db2ddb2d & lut_mask_in) : lut = 64'h59bb314f6a1b1032;
      (64'hd7a2061ea781a781 & lut_mask_in) : lut = 64'h64b84b09a6caee1c;
      (64'h2757823437e137e1 & lut_mask_in) : lut = 64'h76687d45c081d35e;
      (64'hfc13a87ea362a362 & lut_mask_in) : lut = 64'ha1f80960d94080a5;
      (64'he91cceb9853f853f & lut_mask_in) : lut = 64'h9927388855f06d4a;
      (64'h3836fc8710d210d2 & lut_mask_in) : lut = 64'h73215d3db10f9e2d;
      (64'he79793465fc35fc3 & lut_mask_in) : lut = 64'h3fafa69090168923;
      (64'h997b09e5348e348e & lut_mask_in) : lut = 64'h513464008b778438;
      (64'ha1c441a484688468 & lut_mask_in) : lut = 64'h443c74a243d97ad1;
      (64'h6e5be8c3eb04eb04 & lut_mask_in) : lut = 64'h1e4c63b520964c54;
      (64'hba2c2be06caa6caa & lut_mask_in) : lut = 64'h366d1d10053dc228;
      (64'hc6ca3ae126f826f8 & lut_mask_in) : lut = 64'hb0922041f2b00646;
      (64'h18e4656e702c702c & lut_mask_in) : lut = 64'h0bebb555cf064608;
      (64'hc47eabbc95f095f0 & lut_mask_in) : lut = 64'h620938be85fb41e2;
      (64'h3528773cf257f257 & lut_mask_in) : lut = 64'hd68276a79e4ff998;
      (64'hda8c2f1f4c3f4c3f & lut_mask_in) : lut = 64'hfa337f7d8642275a;
      (64'h61176a5ed96bd96b & lut_mask_in) : lut = 64'h0dda524c05af699a;
      (64'hf0e67df3258d258d & lut_mask_in) : lut = 64'hb40b35d6a9268f43;
      (64'h9299781877b077b0 & lut_mask_in) : lut = 64'hda16e6be08d59342;
      (64'h1f2c02fcf18bf18b & lut_mask_in) : lut = 64'h0305fac215c4b7e8;
      (64'hca0a5d75f608f608 & lut_mask_in) : lut = 64'h4b24aef03e27815d;
      (64'h89255425bfa4bfa4 & lut_mask_in) : lut = 64'h33a1a4fe831f026d;
      (64'h846aa033ca38ca38 & lut_mask_in) : lut = 64'h2e13c3593334618c;
      (64'h9275187040a940a9 & lut_mask_in) : lut = 64'he63652727c677514;
      (64'ha236ed2b3a063a06 & lut_mask_in) : lut = 64'h4a430afc1373a892;
      (64'hc4e99fce6d3b6d3b & lut_mask_in) : lut = 64'h629ba61ff05ac3d1;
      (64'hf8c3dc1d58305830 & lut_mask_in) : lut = 64'h322de1d0c4a3f532;
      (64'h99d14a57e51fe51f & lut_mask_in) : lut = 64'h8c7c8cd70e057de4;
      (64'h66f646d98d568d56 & lut_mask_in) : lut = 64'ha62c8c4b3d39c09f;
      (64'h35f899db2dbd2dbd & lut_mask_in) : lut = 64'h55feb1e576602d1b;
      (64'h164ba400e959e959 & lut_mask_in) : lut = 64'ha8e7863f105dc6dd;
      (64'hd195e2b8006a006a & lut_mask_in) : lut = 64'hb3b2d623716d92fe;
      (64'hcf1d9b3959445944 & lut_mask_in) : lut = 64'h542f9bea562c871c;
      (64'h914fed32b97cb97c & lut_mask_in) : lut = 64'hef558921767717c4;
      (64'h02e7d905a961a961 & lut_mask_in) : lut = 64'hf7918b8d8d92b437;
      (64'ha63d5be33d383d38 & lut_mask_in) : lut = 64'h9769a066b9e91b4a;
      (64'hd36298cd59a659a6 & lut_mask_in) : lut = 64'h27eda4526e70f1a4;
      (64'h8c765e91c4b8c4b8 & lut_mask_in) : lut = 64'haa8a1de1c678a64b;
      (64'h8066828f2a4f2a4f & lut_mask_in) : lut = 64'h4438b2c77befb22c;
      (64'h0947edb1e953e953 & lut_mask_in) : lut = 64'haf93ba894da520df;
      (64'h2729de916b326b32 & lut_mask_in) : lut = 64'h96b95154d97f1682;
      (64'h710f7837d4c0d4c0 & lut_mask_in) : lut = 64'h01c6621ba0af962d;
      (64'he55b6e468c538c53 & lut_mask_in) : lut = 64'h4213473e4281da88;
      (64'hbddcf593ac26ac26 & lut_mask_in) : lut = 64'h16041820f9f8dc6b;
      (64'he27b6e7910bc10bc & lut_mask_in) : lut = 64'hd285d593b2a233f7;
      (64'hc95658e3dad1dad1 & lut_mask_in) : lut = 64'ha741506bd6f0492b;
      (64'h197aac36feabfeab & lut_mask_in) : lut = 64'hbfed47b18941aa54;
      (64'heb25634fc6bbc6bb & lut_mask_in) : lut = 64'h4d6bfb92a8fbccad;
      (64'h0e4be592369e369e & lut_mask_in) : lut = 64'h5ab54e7608429f56;
      (64'hd82137fd892f892f & lut_mask_in) : lut = 64'h4fbce5841c2d9fa1;
      (64'hc728ff99963e963e & lut_mask_in) : lut = 64'h49dd933f866252ea;
      (64'h54a36087ee63ee63 & lut_mask_in) : lut = 64'h07059fa1699cc63b;
      (64'hdff8fd32db24db24 & lut_mask_in) : lut = 64'hc7e4557649e81c98;
      (64'h990871513d343d34 & lut_mask_in) : lut = 64'h3fdc41c2eea3f46c;
      (64'h86a9939e21762176 & lut_mask_in) : lut = 64'hcd87d3983562e27b;
      (64'h8be28bf1d038d038 & lut_mask_in) : lut = 64'h418879cf97e9cf40;
      (64'h31326a7941544154 & lut_mask_in) : lut = 64'h21810362fd22d8a7;
      (64'h8fcbc706f715f715 & lut_mask_in) : lut = 64'h9011fc0041ff5e6c;
      (64'he469899ab17fb17f & lut_mask_in) : lut = 64'h6aea190cb565ce0c;
      (64'hbf0a54360c6e0c6e & lut_mask_in) : lut = 64'hb698bf0c21754986;
      (64'h24f8ea96266f266f & lut_mask_in) : lut = 64'h3acb10453b632af5;
      (64'h47d5f2c4547b547b & lut_mask_in) : lut = 64'he611c9d96afcf9e9;
      (64'h2fb97d3175407540 & lut_mask_in) : lut = 64'h031b449a30ba3f5d;
      (64'hc97503d1e089e089 & lut_mask_in) : lut = 64'hb60fd1bc507b3b59;
      (64'h4bc4ca4477d577d5 & lut_mask_in) : lut = 64'h5c7b6926610c67d3;
      (64'h16daad9c5b255b25 & lut_mask_in) : lut = 64'h7e2fd5113d69482b;
      (64'heaa17867dae4dae4 & lut_mask_in) : lut = 64'h1309f8b8052d2a31;
      (64'hfdc2f562d2cbd2cb & lut_mask_in) : lut = 64'h143b9008855c056a;
      (64'hc597524b40364036 & lut_mask_in) : lut = 64'h58446ce1861b518f;
      (64'hf1f40263c31dc31d & lut_mask_in) : lut = 64'h43db01ad63a1dafa;
      (64'h6cbd1c6dc6c7c6c7 & lut_mask_in) : lut = 64'hbd7c0582ebc5196f;
      (64'h5c09543c570d570d & lut_mask_in) : lut = 64'h9f49ac86529490eb;
      (64'h97a0a15b2de02de0 & lut_mask_in) : lut = 64'ha9d41d41a35496a6;
      (64'ha908cda7e82de82d & lut_mask_in) : lut = 64'hef477a7aa0086dd8;
      (64'hce0456d9fbdafbda & lut_mask_in) : lut = 64'h88d2c999d3a4a373;
      (64'hb4e3ae4eb466b466 & lut_mask_in) : lut = 64'he81718c3502ea43b;
      (64'h75b04f97cd79cd79 & lut_mask_in) : lut = 64'h20dd69d19a1f92f7;
      (64'hc672957bf08af08a & lut_mask_in) : lut = 64'h5c093042bfd071d2;
      (64'h12ab822b04190419 & lut_mask_in) : lut = 64'hd56eee407fa4a9c3;
      (64'h83cc4b0629702970 & lut_mask_in) : lut = 64'h3c82d8336395d03d;
      (64'h23cbb1738b6e8b6e & lut_mask_in) : lut = 64'h236f0235cfc2f284;
      (64'hcd0f50dc1cf71cf7 & lut_mask_in) : lut = 64'hc378394c3355ac59;
      (64'h972901ceb077b077 & lut_mask_in) : lut = 64'hfee923bf68bc24a7;
      (64'h0ff0b3d35a205a20 & lut_mask_in) : lut = 64'ha49e4900bdf97f32;
      (64'hcfcb9795fc20fc20 & lut_mask_in) : lut = 64'h85300e241a00298d;
      (64'h0bda28f1ae4fae4f & lut_mask_in) : lut = 64'h2f87d474cafd1a39;
      (64'hf6f26536ec40ec40 & lut_mask_in) : lut = 64'h8cf26f81a721ad2e;
      (64'h26ed65d76cdc6cdc & lut_mask_in) : lut = 64'hfcaca2917d90c111;
      (64'h68518596f47ff47f & lut_mask_in) : lut = 64'h6d97559f5cb0cc76;
      (64'h86370daff9d0f9d0 & lut_mask_in) : lut = 64'h6454ff5d20faa5a1;
      (64'h21c4e5d1dd19dd19 & lut_mask_in) : lut = 64'h24bb09e7db79d089;
      (64'ha03aa7e4cf63cf63 & lut_mask_in) : lut = 64'h53aa5b97b4ab7dfa;
      (64'hb94def70718f718f & lut_mask_in) : lut = 64'h2f4062cb6d8d7b33;
      (64'hd15e2105a48ea48e & lut_mask_in) : lut = 64'he1bd35f257c49cc1;
      (64'h21736d78c83ac83a & lut_mask_in) : lut = 64'h11576d61446930ca;
      (64'hb11ca0df70f770f7 & lut_mask_in) : lut = 64'h37318b7e7a1fcd3d;
      (64'hd1108fcc9dd49dd4 & lut_mask_in) : lut = 64'h69cd9b2435af9643;
      (64'h9a8e4c88d730d730 & lut_mask_in) : lut = 64'h8d02acfe1460fd6d;
      (64'h765eb654c697c697 & lut_mask_in) : lut = 64'hbde71953b6d04718;
      (64'h71cb9e860dfd0dfd & lut_mask_in) : lut = 64'h038cfd9fc6aacfa6;
      (64'hf40ffef664da64da & lut_mask_in) : lut = 64'h23e6d579d5e93a8c;
      (64'hfc1ce8ec3aff3aff & lut_mask_in) : lut = 64'h25f0d6304daaa346;
      (64'h8b9fb1613b823b82 & lut_mask_in) : lut = 64'hdc6ea8c4ff149c0c;
      (64'h96a0dbb6ff62ff62 & lut_mask_in) : lut = 64'h8db04d570024e4ac;
      (64'h33674301b6f6b6f6 & lut_mask_in) : lut = 64'h72a8595b2168d3e4;
      (64'h96a1893fe376e376 & lut_mask_in) : lut = 64'h07162bf985ef3aae;
      (64'h76375c6785628562 & lut_mask_in) : lut = 64'h02838180c1964fdb;
      (64'h9333213a06790679 & lut_mask_in) : lut = 64'h77c71e8f99a41421;
      (64'hebfdca620b720b72 & lut_mask_in) : lut = 64'h1a1fed2117ca3211;
      (64'h6c232151a4ffa4ff & lut_mask_in) : lut = 64'h3f47e57012627c18;
      (64'hee33651b6fb46fb4 & lut_mask_in) : lut = 64'h9c793ef6f7da89b1;
      (64'h8875eacea7a2a7a2 & lut_mask_in) : lut = 64'h23ea28798136c2b3;
      (64'hddda087f96549654 & lut_mask_in) : lut = 64'hcc51fbda462c2e4f;
      (64'h5b1f19ca8bed8bed & lut_mask_in) : lut = 64'hbb557abb564f619c;
      (64'hcae4f9efb15fb15f & lut_mask_in) : lut = 64'h7d52b72bedbf5941;
      (64'h3369ad4b090b090b & lut_mask_in) : lut = 64'hdbdd5834fdcf6cb1;
      (64'hbacd8fefc409c409 & lut_mask_in) : lut = 64'h50eb6436d1d62248;
      (64'h455487c72cd62cd6 & lut_mask_in) : lut = 64'h1ff0cf986ecab70b;
      (64'haf53023b98759875 & lut_mask_in) : lut = 64'he0251ace63e8a81a;
      (64'h976eaee64a044a04 & lut_mask_in) : lut = 64'he2b8b87cd7d4f5ab;
      (64'h6c9ebcb269886988 & lut_mask_in) : lut = 64'h2d0022e2de140361;
      (64'h0abe6a7c80a780a7 & lut_mask_in) : lut = 64'h87c1b4045ecc59d3;
      (64'hb69295b9906f906f & lut_mask_in) : lut = 64'h9a12dfacf0db2dbd;
      (64'hf0c3495e895e895e & lut_mask_in) : lut = 64'h7d29797ba05aade1;
      (64'h66a934a9a097a097 & lut_mask_in) : lut = 64'h62d936d32ce0158e;
      (64'hcaa3a43130673067 & lut_mask_in) : lut = 64'hdb173d08df2d9f14;
      (64'hd3a2ec9bd1b1d1b1 & lut_mask_in) : lut = 64'h67e38868d38f339a;
      (64'hb6fa7d52dd86dd86 & lut_mask_in) : lut = 64'hbdca1b2f054d0df3;
      (64'hf9d64ebb9ffd9ffd & lut_mask_in) : lut = 64'h3d912009da4d5c9b;
      (64'h6ab82cc1d268d268 & lut_mask_in) : lut = 64'h25a400e626086474;
      (64'h70a2567aab2cab2c & lut_mask_in) : lut = 64'h37c13fe2c8aaccdd;
      (64'h0dcf9b07f53af53a & lut_mask_in) : lut = 64'ha95ae3298497c3e7;
      (64'h3a5d70e2d085d085 & lut_mask_in) : lut = 64'h5b284f9bb602e3bd;
      (64'h973edc2bdb55db55 & lut_mask_in) : lut = 64'he3a06add068e87be;
      (64'hecdc2da9da6dda6d & lut_mask_in) : lut = 64'h32294ded9e956f6d;
      (64'h910b46af4ad34ad3 & lut_mask_in) : lut = 64'he04bfb52ea3b8d9f;
      (64'he482637a726f726f & lut_mask_in) : lut = 64'h537c721fe8c34bfd;
      (64'hbc03277210601060 & lut_mask_in) : lut = 64'haa9713b86072a7bc;
      (64'h777fbd3717c417c4 & lut_mask_in) : lut = 64'hf3705456b1a76df4;
      (64'he728595561806180 & lut_mask_in) : lut = 64'hcda426deda781bb8;
      (64'h77add8ec417b417b & lut_mask_in) : lut = 64'hd461de7507d3250b;
      (64'h480e3bc209520952 & lut_mask_in) : lut = 64'h6206ca484d3ca137;
      (64'h9a12814ffdcdfdcd & lut_mask_in) : lut = 64'hb14ef2ed9ba33320;
      (64'h9aa1b152aaf1aaf1 & lut_mask_in) : lut = 64'h36fa8916a51aea98;
      (64'hd35892f7bbe7bbe7 & lut_mask_in) : lut = 64'h23e7171ff8d3439d;
      (64'h63fc235053405340 & lut_mask_in) : lut = 64'h469845b4be813e62;
      (64'hb329b6d295669566 & lut_mask_in) : lut = 64'h365f0f6ec060583f;
      (64'h1f96ae6b7d1f7d1f & lut_mask_in) : lut = 64'he6d69bcd0da4ecf9;
      (64'h2f2224e0aacbaacb & lut_mask_in) : lut = 64'h289de535bf669f17;
      (64'hdfaf60b811301130 & lut_mask_in) : lut = 64'hd33fa41aaefa5cae;
      (64'h3302d74573fe73fe & lut_mask_in) : lut = 64'hbd6823e503b7fac2;
      (64'ha5521d9755f755f7 & lut_mask_in) : lut = 64'hee4e92d9aa41e193;
      (64'hf88e4859e608e608 & lut_mask_in) : lut = 64'h1f34a82960ab66c2;
      (64'hc28fb77a38ed38ed & lut_mask_in) : lut = 64'hdb735b489bcf712a;
      (64'h7327744958005800 & lut_mask_in) : lut = 64'ha32e4c325d871d2c;
      (64'hd80038e796f796f7 & lut_mask_in) : lut = 64'h1a53de8114ed0ea7;
      (64'h186a485665d565d5 & lut_mask_in) : lut = 64'hda4d17368b1cdfda;
      (64'hbcd7187dc0e2c0e2 & lut_mask_in) : lut = 64'h544d754eae8ccf40;
      (64'hdd18c95445844584 & lut_mask_in) : lut = 64'h247325de73ac6da1;
      (64'hfc1200ca000e000e & lut_mask_in) : lut = 64'h84d48ba7ac5e3731;
      (64'hdde88f82aaa0aaa0 & lut_mask_in) : lut = 64'hc1b636ef27bac573;
      (64'h6a56ccdf16081608 & lut_mask_in) : lut = 64'ha40075ef472f6da4;
      (64'hb06c3d267e177e17 & lut_mask_in) : lut = 64'h293f9d64205c8498;
      (64'hcc3227a954c354c3 & lut_mask_in) : lut = 64'ha5e6f52e55f709cc;
      (64'hfc16b851dc65dc65 & lut_mask_in) : lut = 64'h37acedc915bc1e3c;
      (64'h5d4625b870017001 & lut_mask_in) : lut = 64'hcd7cf57c1e6ec4ac;
      (64'h6f0ab9d18e4f8e4f & lut_mask_in) : lut = 64'h8c52714dfedd0734;
      (64'h69c68051e679e679 & lut_mask_in) : lut = 64'h0b116d6c1b1a7a25;
      (64'h033195e123882388 & lut_mask_in) : lut = 64'hf794fb27a79c9e92;
      (64'h7ab31a11cc1acc1a & lut_mask_in) : lut = 64'ha2a5f551b6cbaccc;
      (64'h05ba2a7bd1fcd1fc & lut_mask_in) : lut = 64'h32636d1359b81e0a;
      (64'h33da431138873887 & lut_mask_in) : lut = 64'h64b6f563fa1e55bd;
      (64'h4ce817244ea94ea9 & lut_mask_in) : lut = 64'h28d18a0c52d24cb6;
      (64'h2b6fc83569576957 & lut_mask_in) : lut = 64'h19753838995b9ea9;
      (64'h83ea57e1d04fd04f & lut_mask_in) : lut = 64'h3cecaeae46b3a6a7;
      (64'h7012c9a801870187 & lut_mask_in) : lut = 64'ha52bceee4e13d65c;
      (64'hf041cd2367df67df & lut_mask_in) : lut = 64'h6d9c4f1abfc94cbf;
      (64'hc8fb227f76307630 & lut_mask_in) : lut = 64'hcb081e793b25140c;
      (64'h14c894f754b554b5 & lut_mask_in) : lut = 64'hb59eaf8a071f67f1;
      (64'h1bd3d3fb62976297 & lut_mask_in) : lut = 64'he8815b50159ec068;
      (64'ha5baa440aa0eaa0e & lut_mask_in) : lut = 64'h4a6a661ef22557ee;
      (64'h4c3a8beca761a761 & lut_mask_in) : lut = 64'h5fd4ae8fc9637b4c;
      (64'h696d5a83f4a2f4a2 & lut_mask_in) : lut = 64'he88e801cf6e6b239;
      (64'h5d55f913bffabffa & lut_mask_in) : lut = 64'h5cf66ff5aaf386e3;
      (64'h7575529bf50bf50b & lut_mask_in) : lut = 64'h8cd842387dc564ac;
      (64'h341be870a5c7a5c7 & lut_mask_in) : lut = 64'hae0c976d800fe890;
      (64'h18e1c303e55de55d & lut_mask_in) : lut = 64'h4f2e4a4ee81b84f4;
      (64'h53e07d8f43674367 & lut_mask_in) : lut = 64'hd52977045e00b576;
      (64'h9c31856435f035f0 & lut_mask_in) : lut = 64'h382a86ae02005665;
      (64'h00a988082c0c2c0c & lut_mask_in) : lut = 64'hc05aa089237889a6;
      (64'h016d80dcec5eec5e & lut_mask_in) : lut = 64'hd870f0db7a09d907;
      (64'h4e97e1c80fe10fe1 & lut_mask_in) : lut = 64'hb0c56715ec19ac12;
      (64'h9ffe775580dd80dd & lut_mask_in) : lut = 64'h429e9a0306731828;
      (64'hb2c69d8945334533 & lut_mask_in) : lut = 64'h7dc716cb717a1a82;
      (64'h37a59f481d0b1d0b & lut_mask_in) : lut = 64'hb76ee19095b94393;
      (64'h9697b848d3a4d3a4 & lut_mask_in) : lut = 64'hc2206c81b67bb8a2;
      (64'h1d5cf7f9c814c814 & lut_mask_in) : lut = 64'heebb4163d79bad2e;
      (64'h855a5ae5b280b280 & lut_mask_in) : lut = 64'hec101fe4d43de8dc;
      (64'h01dc492c2d2b2d2b & lut_mask_in) : lut = 64'h0a0ee0363b051ddb;
      (64'h5370358397549754 & lut_mask_in) : lut = 64'h4ccf610fa327eb85;
      (64'h9987bcaf456d456d & lut_mask_in) : lut = 64'h6afe22628ebd9621;
      (64'h8ff588701f891f89 & lut_mask_in) : lut = 64'he6e34385bd26336f;
      (64'hb27b6f2463ce63ce & lut_mask_in) : lut = 64'h50f1401d6224c3cb;
      (64'h6af23a92a5f6a5f6 & lut_mask_in) : lut = 64'had3f29708e7a61b0;
      (64'hcbc3353bb995b995 & lut_mask_in) : lut = 64'hf11f462807c172f0;
      (64'h1eac4dce071e071e & lut_mask_in) : lut = 64'h7a0a85069c9bb8f7;
      (64'hecd226a07efa7efa & lut_mask_in) : lut = 64'h21438be719bf0fdf;
      (64'h6207f0645d715d71 & lut_mask_in) : lut = 64'h9a3523befa6dbe69;
      (64'h126b37f6b5edb5ed & lut_mask_in) : lut = 64'h0a1cbd54432e5d82;
      (64'h5621d09ae35de35d & lut_mask_in) : lut = 64'hb586a15022fbb17b;
      (64'he775764201ab01ab & lut_mask_in) : lut = 64'h9097e55ecfbac818;
      (64'hddfab438bb94bb94 & lut_mask_in) : lut = 64'haa05e7f1eb7b6b6d;
      (64'hb883606d0ad00ad0 & lut_mask_in) : lut = 64'h87f6b1321d64d34b;
      (64'hbb9029692d102d10 & lut_mask_in) : lut = 64'h1da24c2cada516fe;
      (64'h031d97dca052a052 & lut_mask_in) : lut = 64'h4feb128e369ba11f;
      (64'hda91f930a2faa2fa & lut_mask_in) : lut = 64'hec24011800616770;
      (64'h4c834f31cffbcffb & lut_mask_in) : lut = 64'h9756b71c730a42a9;
      (64'he68ec8ada13fa13f & lut_mask_in) : lut = 64'h9b2f3dbae6b09554;
      (64'h6f544b734c1b4c1b & lut_mask_in) : lut = 64'ha91275ebc0180f42;
      (64'ha7fbeb8db0a4b0a4 & lut_mask_in) : lut = 64'h1aef4a5c39fd5740;
      (64'hffa36c1de510e510 & lut_mask_in) : lut = 64'h39672c7300695c78;
      (64'h3c56c5457de07de0 & lut_mask_in) : lut = 64'hb52cc6f7a6c458db;
      (64'hc03f8ee230ba30ba & lut_mask_in) : lut = 64'h7a055ede54069b4e;
      (64'h620a0edb11e611e6 & lut_mask_in) : lut = 64'h5377871c92769a04;
      (64'hc01dc51c2f722f72 & lut_mask_in) : lut = 64'hdbc20f5d442dd4e2;
      (64'h86b2b5e7e939e939 & lut_mask_in) : lut = 64'h167e73f9843b2498;
      (64'hafdacdbaba62ba62 & lut_mask_in) : lut = 64'h5927b2db4162344b;
      (64'h2681417f7dc97dc9 & lut_mask_in) : lut = 64'h69ecfe6887801486;
      (64'hd1c63bf31d3f1d3f & lut_mask_in) : lut = 64'h0582a3d11e17455d;
      (64'hd4699ffd42dc42dc & lut_mask_in) : lut = 64'h2822ec5e51a05685;
      (64'h624a0808ae89ae89 & lut_mask_in) : lut = 64'h4435b86e0a27fd98;
      (64'hd52d310bd601d601 & lut_mask_in) : lut = 64'h254ef6c12ece991c;
      (64'h49af4a1b05d905d9 & lut_mask_in) : lut = 64'he6c3e99ff8799384;
      (64'h3c4443f71e551e55 & lut_mask_in) : lut = 64'h2b37f87ea585cca9;
      (64'h3b3b29d0824b824b & lut_mask_in) : lut = 64'h26290128cd2fa072;
      (64'hb56f6c622bb42bb4 & lut_mask_in) : lut = 64'h154cd7c2edbfb908;
      (64'h9a975a6471e271e2 & lut_mask_in) : lut = 64'h45b7928094e26a9d;
      (64'h71c0ff61b97db97d & lut_mask_in) : lut = 64'haa81dfb0a5792dc0;
      (64'h5fc92329f76af76a & lut_mask_in) : lut = 64'h616f732ca6c7a183;
      (64'hbad4d5e981248124 & lut_mask_in) : lut = 64'he629daf8decaf362;
      (64'h3cc495886c016c01 & lut_mask_in) : lut = 64'hcc87ffd068c79aed;
      (64'h7b68cc28bb80bb80 & lut_mask_in) : lut = 64'hf2e1a29dece81f02;
      (64'ha40aa14cea9aea9a & lut_mask_in) : lut = 64'h9dc57f4d8883af76;
      (64'h05902f9d271c271c & lut_mask_in) : lut = 64'h450fc62796455957;
      (64'hb9b11735c26ec26e & lut_mask_in) : lut = 64'he521475842d35172;
      (64'had9de5c0eed3eed3 & lut_mask_in) : lut = 64'hf49d4d25508c435f;
      (64'h2e6ea57e76bf76bf & lut_mask_in) : lut = 64'hb793584fe584578c;
      (64'h6ddc41ed06ac06ac & lut_mask_in) : lut = 64'h8f718b9f4858b403;
      (64'h63fb5c5316791679 & lut_mask_in) : lut = 64'he376e5adafd108d0;
      (64'h2b4b95709a609a60 & lut_mask_in) : lut = 64'h64cc08714444773c;
      (64'hf7eb9a4f439a439a & lut_mask_in) : lut = 64'hc72726c2aa089303;
      (64'h599bf3aa534f534f & lut_mask_in) : lut = 64'h3ad827c68518da91;
      (64'hdcde52017d967d96 & lut_mask_in) : lut = 64'h5708af0ca96e8d3d;
      (64'hc3e0d9a012c812c8 & lut_mask_in) : lut = 64'ha23aac0d5d03d238;
      (64'h51adc216221c221c & lut_mask_in) : lut = 64'h8168374cc2f06421;
      (64'h8a97f4f76c6d6c6d & lut_mask_in) : lut = 64'ha5915a6c2638e858;
      (64'h75f7114f965f965f & lut_mask_in) : lut = 64'h43ead1b6d729b914;
      (64'hfda0d7684b594b59 & lut_mask_in) : lut = 64'h1a87cbbd4bba1642;
      (64'h798ad0e93db73db7 & lut_mask_in) : lut = 64'hccd041302609715f;
      (64'h2592721edd58dd58 & lut_mask_in) : lut = 64'hf331c52886fab3dd;
      (64'h8b7e3079d383d383 & lut_mask_in) : lut = 64'hfa12128907f33247;
      (64'hb7d5dd4c51c351c3 & lut_mask_in) : lut = 64'h1f7af80db9010f55;
      (64'h111bbb840ad40ad4 & lut_mask_in) : lut = 64'h73ee5fdcf1000617;
      (64'h39150e4afd35fd35 & lut_mask_in) : lut = 64'hd82dc4d6b8d99b4c;
      (64'h8f789af6a3c9a3c9 & lut_mask_in) : lut = 64'hd1c47498f7723670;
      (64'h83b9ce1f16c616c6 & lut_mask_in) : lut = 64'h413a733700110897;
      (64'h01a06e3b21672167 & lut_mask_in) : lut = 64'hcc948590f971eb1d;
      (64'h722941cef68ff68f & lut_mask_in) : lut = 64'haadf1098a136e5d3;
      (64'h000f3b7351cd51cd & lut_mask_in) : lut = 64'h6dedc16f2e54de5e;
      (64'h47081b8ba33fa33f & lut_mask_in) : lut = 64'h2d0ea5d442ad87b8;
      (64'hab0425198ce68ce6 & lut_mask_in) : lut = 64'h0b0d838e4553d17c;
      (64'h4668827e7a0b7a0b & lut_mask_in) : lut = 64'h3ef3a835a71a6c6a;
      (64'h33edddcaa54da54d & lut_mask_in) : lut = 64'h5fd9fb311c351035;
      (64'h1ecfcf6166d966d9 & lut_mask_in) : lut = 64'h16be9d4896aede7b;
      (64'hcdc92a0935603560 & lut_mask_in) : lut = 64'hd3e0b53dc1264e22;
      (64'h77854c2641534153 & lut_mask_in) : lut = 64'h36a3d7f9d0ead140;
      (64'hcfb2181fc14dc14d & lut_mask_in) : lut = 64'ha21f802ba62bb7df;
      (64'ha681ce04d312d312 & lut_mask_in) : lut = 64'haf066f3fd75a8dab;
      (64'h6e7ed69b55bb55bb & lut_mask_in) : lut = 64'h88fb3f7ab3fb42c1;
      (64'ha09016cf9ac99ac9 & lut_mask_in) : lut = 64'hc203736cfeec5bec;
      (64'h897285c942514251 & lut_mask_in) : lut = 64'h496e5feb45a9c023;
      (64'he9f0eb44efc3efc3 & lut_mask_in) : lut = 64'h1babb6cc44e39787;
      (64'hf688881c0ef70ef7 & lut_mask_in) : lut = 64'hf441aace590a80d1;
      (64'h5a910676b3d7b3d7 & lut_mask_in) : lut = 64'h4c15a52d54e9180e;
      (64'h73f82c3900ab00ab & lut_mask_in) : lut = 64'he1b2aea570f0d24f;
      (64'h4c70a74fe4c5e4c5 & lut_mask_in) : lut = 64'h8bd603b1cf885f78;
      (64'hbc3791f27a267a26 & lut_mask_in) : lut = 64'h0b2f776eb5efd502;
      (64'ha9b63b9c8ea18ea1 & lut_mask_in) : lut = 64'hc69a5d52eab200e5;
      (64'h3d2cdace28cd28cd & lut_mask_in) : lut = 64'h7971ba0c1e3e4057;
      (64'h80d82a61c1dfc1df & lut_mask_in) : lut = 64'h554e4b7ed4802365;
      (64'hd32f948944f544f5 & lut_mask_in) : lut = 64'hbc664b68e25dd297;
      (64'hbe69fd836fd96fd9 & lut_mask_in) : lut = 64'h39e76824d0250b9a;
      (64'h809c7c483e783e78 & lut_mask_in) : lut = 64'hefe2a5c8a5949370;
      (64'ha65c198957655765 & lut_mask_in) : lut = 64'h94ea0921044f00a7;
      (64'hc736aaf5adaaadaa & lut_mask_in) : lut = 64'h680cac0cef39d574;
      (64'h0d3c29f28e738e73 & lut_mask_in) : lut = 64'h6c87144344351bcd;
      (64'h21e1154f5d145d14 & lut_mask_in) : lut = 64'h13358a6504174b98;
      (64'h0ab629a4f9e1f9e1 & lut_mask_in) : lut = 64'ha441477e013149eb;
      (64'h0872e06543084308 & lut_mask_in) : lut = 64'h1c06c7eb979194b7;
      (64'hff8edbb3d67cd67c & lut_mask_in) : lut = 64'he75d15085bf8f1ac;
      (64'h0967bd35748e748e & lut_mask_in) : lut = 64'h642881332e766d94;
      (64'hcd228aaa57135713 & lut_mask_in) : lut = 64'h5d37c6f684127df9;
      (64'hebf6eaeebd0dbd0d & lut_mask_in) : lut = 64'h2bc3d7e550506840;
      (64'h976937d5d691d691 & lut_mask_in) : lut = 64'h1dcba12f7289a618;
      (64'hbb30050d029a029a & lut_mask_in) : lut = 64'h87271a19232076a0;
      (64'h797144fddd1ddd1d & lut_mask_in) : lut = 64'h83e45c48da5a2254;
      (64'h56151a76aee5aee5 & lut_mask_in) : lut = 64'h5a7dbaf977b78206;
      (64'h3398ffed45e945e9 & lut_mask_in) : lut = 64'hf2b02edacc69572e;
      (64'h49840eb3f33bf33b & lut_mask_in) : lut = 64'h81dbb325dd0989b9;
      (64'h83458ceac613c613 & lut_mask_in) : lut = 64'heaa1654aec4f5ae2;
      (64'h7f27225e2a002a00 & lut_mask_in) : lut = 64'h2cb20905811616a0;
      (64'h3bab5be5a6fba6fb & lut_mask_in) : lut = 64'hf867211d09b896e6;
      (64'h8de83ad9b9c9b9c9 & lut_mask_in) : lut = 64'he433d796652eb60a;
      (64'h6fe5002c45df45df & lut_mask_in) : lut = 64'h002dbf091aba242d;
      (64'hca81a9ef5d985d98 & lut_mask_in) : lut = 64'he954447ed72efd97;
      (64'hb391ac6fa7c4a7c4 & lut_mask_in) : lut = 64'h2a76f775521d0eb4;
      (64'h9c89c47b5a095a09 & lut_mask_in) : lut = 64'hc8b25d1061981ab5;
      (64'h862129b23e463e46 & lut_mask_in) : lut = 64'he87b6ff32b43f32d;
      (64'h139bfa9067116711 & lut_mask_in) : lut = 64'h786468d5783a6452;
      (64'h44e31230b955b955 & lut_mask_in) : lut = 64'h043fc33174dabb9d;
      (64'hf1d4cef3ae4cae4c & lut_mask_in) : lut = 64'h4a4abbac9fafcf3c;
      (64'h872e6a9d1f901f90 & lut_mask_in) : lut = 64'h61c9bf7b71711dec;
      (64'hf48eef9043004300 & lut_mask_in) : lut = 64'hfca9b513a320cbfe;
      (64'h82acdc9bcddccddc & lut_mask_in) : lut = 64'h690abee3cf580bb9;
      (64'h12f54f7e5c6e5c6e & lut_mask_in) : lut = 64'hd0a96eab2145c9c3;
      (64'h51f147ca4c134c13 & lut_mask_in) : lut = 64'he0e34cb4f169dc3c;
      (64'h26ce613d80708070 & lut_mask_in) : lut = 64'h501711564b90b99a;
      (64'h8cfc384245824582 & lut_mask_in) : lut = 64'hc514000ae7142990;
      (64'h0901ab8e77317731 & lut_mask_in) : lut = 64'h9b6f10892f8d53ab;
      (64'h7864b0d951f851f8 & lut_mask_in) : lut = 64'hc6cf2aeb9a8f18f5;
      (64'ha92473401a1f1a1f & lut_mask_in) : lut = 64'h043179082650b9a1;
      (64'he0f233ff00490049 & lut_mask_in) : lut = 64'hc538b5d550096adb;
      (64'h62eee3fec247c247 & lut_mask_in) : lut = 64'h8e311081bf951d26;
      (64'h005e453ad1ded1de & lut_mask_in) : lut = 64'hbf8ab40579d136a8;
      (64'h083bfdd24e9d4e9d & lut_mask_in) : lut = 64'h77105ab6c76f5fd1;
      (64'h971eeaba29ad29ad & lut_mask_in) : lut = 64'h0e9a95a779875561;
      (64'heeeecc07445f445f & lut_mask_in) : lut = 64'hd3fd8e04fcd386d4;
      (64'hda81bad4c536c536 & lut_mask_in) : lut = 64'hae3961b8bf9b6f1c;
      (64'h67b733c37ce67ce6 & lut_mask_in) : lut = 64'h77fcc8557f1b4469;
      (64'h31875e9bfa5ffa5f & lut_mask_in) : lut = 64'h4c0921babfa59be4;
      (64'h6e0a0b72afb8afb8 & lut_mask_in) : lut = 64'h462745d3280c7c81;
      (64'ha607dc81727b727b & lut_mask_in) : lut = 64'h35ece773c1072f79;
      (64'hf43e572ffe56fe56 & lut_mask_in) : lut = 64'h3b8d7b0f232d4929;
      (64'h284eaa62caa2caa2 & lut_mask_in) : lut = 64'heae62e0f995f3590;
      (64'h585adf3656ac56ac & lut_mask_in) : lut = 64'h9e1b1a92c98cb94a;
      (64'h30d822d256705670 & lut_mask_in) : lut = 64'had7f16573697ecfe;
      (64'hae9298ef38653865 & lut_mask_in) : lut = 64'h099ccaf253060018;
      (64'h7bd214d0a8cba8cb & lut_mask_in) : lut = 64'h7b25a486b82919f3;
      (64'h977ec416d6b1d6b1 & lut_mask_in) : lut = 64'h2bcef641d0a0f16f;
      (64'h0d4e12a416f216f2 & lut_mask_in) : lut = 64'h3b34bddac092bc23;
      (64'h114eeb7b73d073d0 & lut_mask_in) : lut = 64'hce148d7fd93a4304;
      (64'heda486f786a086a0 & lut_mask_in) : lut = 64'h7d7e77ae3c6eb174;
      (64'h93be0780b10fb10f & lut_mask_in) : lut = 64'h8228ac334f04db63;
      (64'hb047247158e458e4 & lut_mask_in) : lut = 64'hd3ac46c3f8a9452a;
      (64'h1ea6dce8e195e195 & lut_mask_in) : lut = 64'h912e74b2ecad5df6;
      (64'h49ef877927f827f8 & lut_mask_in) : lut = 64'hfe6bce35203e2b71;
      (64'h10794bf62cdb2cdb & lut_mask_in) : lut = 64'h2d69da0b42f4b35f;
      (64'hc8db8043e5e5e5e5 & lut_mask_in) : lut = 64'h708841988567b10f;
      (64'h6343015433d333d3 & lut_mask_in) : lut = 64'h36e3c558b4fed195;
      (64'h32fa740d844b844b & lut_mask_in) : lut = 64'hf2c75988ec05c3f0;
      (64'h571e00826ef76ef7 & lut_mask_in) : lut = 64'hd5442fa067de9537;
      (64'hec877a1449414941 & lut_mask_in) : lut = 64'hb319eec0a6a6a842;
      (64'he1ac2fcf619a619a & lut_mask_in) : lut = 64'h5cdb3c0867a7164e;
      (64'h859f400aeef8eef8 & lut_mask_in) : lut = 64'hbb4cb1c0ffacbb36;
      (64'h6a41ad1de450e450 & lut_mask_in) : lut = 64'h031ed15028a20300;
      (64'h01c5d4295d675d67 & lut_mask_in) : lut = 64'h9ebeaf9df7345cca;
      (64'h66bad19042da42da & lut_mask_in) : lut = 64'he95aa42a4a0d66a2;
      (64'h23aa458830f330f3 & lut_mask_in) : lut = 64'h0113a4af2c8498d2;
      (64'ha3e9b6afa71da71d & lut_mask_in) : lut = 64'h5fc8e2be744a4762;
      (64'hbbea50a26a186a18 & lut_mask_in) : lut = 64'hc90e167697922c9b;
      (64'h759ada898d618d61 & lut_mask_in) : lut = 64'h6ff05f4b375b049e;
      (64'hcd6532330f6a0f6a & lut_mask_in) : lut = 64'hb8c0d6d3dc8ddc28;
      (64'ha35265ec26ec26ec & lut_mask_in) : lut = 64'hc7c6d22a4ed28fb7;
      (64'h78ec9ed08c138c13 & lut_mask_in) : lut = 64'h5c1d1fbb37330efd;
      (64'h2d31848872917291 & lut_mask_in) : lut = 64'h90edefe838e71253;
      (64'h7b87f6e6a13ea13e & lut_mask_in) : lut = 64'h16966e85e75014dd;
      (64'hd8a7e87a26502650 & lut_mask_in) : lut = 64'h52f2d0f0c595ccae;
      (64'hd74796075c755c75 & lut_mask_in) : lut = 64'hfd64c779a4267bd8;
      (64'hb84de4fd27ee27ee & lut_mask_in) : lut = 64'h879f72b0f8aacfca;
      (64'h1b48ff9783ff83ff & lut_mask_in) : lut = 64'h517cd0a22ab13923;
      (64'h8fa9be8a11b511b5 & lut_mask_in) : lut = 64'heb0f0f0c4a83af8c;
      (64'hae83560d9fb39fb3 & lut_mask_in) : lut = 64'h8f4d791907654f01;
      (64'he71b0bc9bc56bc56 & lut_mask_in) : lut = 64'h4c96c5e17afad39b;
      (64'h40ce26c8ce98ce98 & lut_mask_in) : lut = 64'he1ccbc04e88dc5c8;
      (64'hc37f35d77b0c7b0c & lut_mask_in) : lut = 64'hbc45af5fcd07e377;
      (64'ha8f483bb71ce71ce & lut_mask_in) : lut = 64'ha72d11ecdb0c6a96;
      (64'h6aa3b7f5bb27bb27 & lut_mask_in) : lut = 64'h25978da015d9fc35;
      (64'h31ed0d4159fb59fb & lut_mask_in) : lut = 64'hb33866903004d0e8;
      (64'hd73a2bb6aaecaaec & lut_mask_in) : lut = 64'h63166771c01f4cee;
      (64'h9301584e85c785c7 & lut_mask_in) : lut = 64'h264180f09c0e2ab0;
      (64'hced2aa17daa2daa2 & lut_mask_in) : lut = 64'h3d68267a83925d35;
      (64'h72757881f26df26d & lut_mask_in) : lut = 64'h1b16518547ca8123;
      (64'h864282a2f3bff3bf & lut_mask_in) : lut = 64'h7c0b39a42df176ee;
      (64'hd8f7f6b0b128b128 & lut_mask_in) : lut = 64'hde1e37909f7664d7;
      (64'h3bc19f4cd007d007 & lut_mask_in) : lut = 64'h391e226d0bbb2846;
      (64'h27d218a182d482d4 & lut_mask_in) : lut = 64'hea5fedd75e635545;
      (64'h30d532fb39583958 & lut_mask_in) : lut = 64'he6be95417fbe0030;
      (64'h7530c5a7f76cf76c & lut_mask_in) : lut = 64'hd0966458f219b3fe;
      (64'h9fb33429fa77fa77 & lut_mask_in) : lut = 64'h27e1e7b5928ea52a;
      (64'hba4d4728d2fed2fe & lut_mask_in) : lut = 64'h217575aa98e347cf;
      (64'he6dcbed62b162b16 & lut_mask_in) : lut = 64'h3dc43a2cfc7493ea;
      (64'hf2e91fb6ef0def0d & lut_mask_in) : lut = 64'he112b56023499f47;
      (64'h44c4898067d567d5 & lut_mask_in) : lut = 64'h61cdc6df9162e024;
      (64'hfe6302640d4f0d4f & lut_mask_in) : lut = 64'h9e5963a7ad022dcc;
      (64'h6237f8c5c445c445 & lut_mask_in) : lut = 64'hc10bb9c3a26d2240;
      (64'h5499d3b9cbafcbaf & lut_mask_in) : lut = 64'hc679fe4a1b011ee0;
      (64'h11df67be7fcc7fcc & lut_mask_in) : lut = 64'hda3a39c98e546952;
      (64'hf8d5179b59ce59ce & lut_mask_in) : lut = 64'ha06fb3125bf68c90;
      (64'h417eed96f470f470 & lut_mask_in) : lut = 64'ha89c5a2e9c29d6e9;
      (64'hdc8db3d60aba0aba & lut_mask_in) : lut = 64'h07a96376b0f4eccd;
      (64'h4a48049a434f434f & lut_mask_in) : lut = 64'h0dad807eed22e680;
      (64'h3696138b0a0f0a0f & lut_mask_in) : lut = 64'hfcd7fde99da9d055;
      (64'habe094907f037f03 & lut_mask_in) : lut = 64'h6113c91cd35201bf;
      (64'hcabb27c0a87ca87c & lut_mask_in) : lut = 64'h565ac3527f36e1ec;
      (64'hd5274ffe8baf8baf & lut_mask_in) : lut = 64'h86d2b205a2f10922;
      (64'h5ee44d52c23dc23d & lut_mask_in) : lut = 64'h7c329319d016d304;
      (64'h8c48d40869986998 & lut_mask_in) : lut = 64'h7880283bd7e10858;
      (64'h676a418c994c994c & lut_mask_in) : lut = 64'h47543128c05d717c;
      (64'h04e4123f85918591 & lut_mask_in) : lut = 64'hf89e6e8d80903213;
      (64'h6b68524d12b012b0 & lut_mask_in) : lut = 64'hb1b2c4d52d098479;
      (64'h67944a61e553e553 & lut_mask_in) : lut = 64'h47cf2015a39760d2;
      (64'hf2a18788d4eed4ee & lut_mask_in) : lut = 64'hbbff8a0a75985261;
      (64'h38e2704a86478647 & lut_mask_in) : lut = 64'heb0cab9de11a7f1b;
      (64'h35d77c2cb02ab02a & lut_mask_in) : lut = 64'h2fa919fcbe8cbdb5;
      (64'hb8f809c2aa6caa6c & lut_mask_in) : lut = 64'hcebab0657f51b377;
      (64'h9af35500ce3ece3e & lut_mask_in) : lut = 64'hb83c94cb1260ed3c;
      (64'hcdd4866e63356335 & lut_mask_in) : lut = 64'ha0a4a731a4581fb1;
      (64'h35938ebd42c142c1 & lut_mask_in) : lut = 64'h940af8d179f16b1d;
      (64'he775261fb52fb52f & lut_mask_in) : lut = 64'h54cb1ed56a17bf3d;
      (64'h1147df6f4d5b4d5b & lut_mask_in) : lut = 64'h52516a79567a7b81;
      (64'he6804c28a764a764 & lut_mask_in) : lut = 64'h4199644a4e5bf563;
      (64'hb4e9ae75bce2bce2 & lut_mask_in) : lut = 64'h949302723c516484;
      (64'h7b9d5102d1ffd1ff & lut_mask_in) : lut = 64'hfd8996713028925d;
      (64'h97624198f41bf41b & lut_mask_in) : lut = 64'h2118f648160ec936;
      (64'h80ebd3d245054505 & lut_mask_in) : lut = 64'hcb53547c1d72ff77;
      (64'h0741df3c72d572d5 & lut_mask_in) : lut = 64'h55a7876e117e6ca2;
      (64'h0785782203d703d7 & lut_mask_in) : lut = 64'h16068dbfcfdcae7a;
      (64'h9164f50645e645e6 & lut_mask_in) : lut = 64'h76e5e23643c363bd;
      (64'h4de4b8f6058b058b & lut_mask_in) : lut = 64'h194029c402abcb67;
      (64'hdbd6cffceb76eb76 & lut_mask_in) : lut = 64'hbc9fa8c39caffd06;
      (64'hd7b96ecbaeaaaeaa & lut_mask_in) : lut = 64'ha048e319414fe7b5;
      (64'h0302ed38270b270b & lut_mask_in) : lut = 64'h36099347449cb566;
      (64'hc72ca27d6ad36ad3 & lut_mask_in) : lut = 64'h8993f29aaf352de3;
      (64'h09771b5344d244d2 & lut_mask_in) : lut = 64'h6b08f73392f46bec;
      (64'h72cc14e3464c464c & lut_mask_in) : lut = 64'h4dd750fac744cea9;
      (64'hf4a55f4d37f137f1 & lut_mask_in) : lut = 64'hb3128d2d522399fb;
      (64'hb8ca99d2b3afb3af & lut_mask_in) : lut = 64'h9168f202d5de00ae;
      (64'hc5235d46e2e0e2e0 & lut_mask_in) : lut = 64'hcb8ac03880f6810d;
      (64'he53c036904640464 & lut_mask_in) : lut = 64'h171876525c2cd035;
      (64'h6e1c65fb48364836 & lut_mask_in) : lut = 64'h9ef8676ac6ee178f;
      (64'h303dca6ef01ff01f & lut_mask_in) : lut = 64'h27ca9c916b9b1864;
      (64'h23b968feb20eb20e & lut_mask_in) : lut = 64'h4305b0cc33c06f41;
      (64'h66c6ff55e4e4e4e4 & lut_mask_in) : lut = 64'h4c0129400d7f6b10;
      (64'h7974065059f659f6 & lut_mask_in) : lut = 64'h2808c961e360b535;
      (64'h3bf54500399b399b & lut_mask_in) : lut = 64'hb08ff32b0a405946;
      (64'h9da3897907d107d1 & lut_mask_in) : lut = 64'h44e8749a47a868fb;
      (64'ha42604ce5e915e91 & lut_mask_in) : lut = 64'hd09798b9115fbd45;
      (64'hcfed6d9a826f826f & lut_mask_in) : lut = 64'hb7355780125fd98a;
      (64'hc7780c0f6f3b6f3b & lut_mask_in) : lut = 64'hcc4f76d53e17b55e;
      (64'h158e859db9ebb9eb & lut_mask_in) : lut = 64'hf2c214807d9e52a7;
      (64'h50d9a68c080d080d & lut_mask_in) : lut = 64'h7e55ab3ae958f1f0;
      (64'h51122451b2ecb2ec & lut_mask_in) : lut = 64'h84317a786caf824c;
      (64'h3624e855d696d696 & lut_mask_in) : lut = 64'h1804db5e7bc1b4cb;
      (64'hac1bb831171d171d & lut_mask_in) : lut = 64'h7885549ae4e82cf6;
      (64'h0ad18030a82da82d & lut_mask_in) : lut = 64'h5423f5ef027f287c;
      (64'hfc1cffff48ef48ef & lut_mask_in) : lut = 64'h6e7a37ff202cd112;
      (64'hbbc3381c7ebf7ebf & lut_mask_in) : lut = 64'h0187b21e2a3b00a0;
      (64'hed5e550d38db38db & lut_mask_in) : lut = 64'hf85e61b248d0ee1b;
      (64'h2c7310c5c4dac4da & lut_mask_in) : lut = 64'h62a3a93313c45378;
      (64'h6facf404e2b9e2b9 & lut_mask_in) : lut = 64'hf61465af968ec217;
      (64'hfa43b0b4212b212b & lut_mask_in) : lut = 64'h004aeb39d75855f7;
      (64'hae6139c1c802c802 & lut_mask_in) : lut = 64'hbe9b3e336331904b;
      (64'h09f0da391be01be0 & lut_mask_in) : lut = 64'ha0effd480dd07d5b;
      (64'hf152ab0d411b411b & lut_mask_in) : lut = 64'hb7b4334b00085ca3;
      (64'h06a4ae4459015901 & lut_mask_in) : lut = 64'h22e38bfb2801f9dd;
      (64'hf91681558a828a82 & lut_mask_in) : lut = 64'hea0f137a64c239bf;
      (64'hadfdaf6b9bff9bff & lut_mask_in) : lut = 64'ha0d4ed42565cfa6a;
      (64'h7618c3a4bff2bff2 & lut_mask_in) : lut = 64'h7fb7f9a04a4131b4;
      (64'ha98ed64ab501b501 & lut_mask_in) : lut = 64'h3776ca8a08d0cd9d;
      (64'h99be658f59825982 & lut_mask_in) : lut = 64'h0d3db362b975af8e;
      (64'h9a182b7e90bc90bc & lut_mask_in) : lut = 64'h3d593fbf07c9bc53;
      (64'h9034cbb738f638f6 & lut_mask_in) : lut = 64'ha15a226b86457827;
      (64'hced93d84d5c4d5c4 & lut_mask_in) : lut = 64'h5538fd5ac8820b54;
      (64'h2ad4e02e6f746f74 & lut_mask_in) : lut = 64'h1b7a4ff099a1f2d5;
      (64'hcad9f8232c392c39 & lut_mask_in) : lut = 64'h767143160d0e7172;
      (64'h7a8ff89a589d589d & lut_mask_in) : lut = 64'hdc2845642e474c8a;
      (64'h7aaff332ac4bac4b & lut_mask_in) : lut = 64'h3cf5f92a0fdb92b2;
      (64'h59980192a686a686 & lut_mask_in) : lut = 64'h809dd01684fc3037;
      (64'hdba2c935d08dd08d & lut_mask_in) : lut = 64'h139481c23075954d;
      (64'h635b9602f1ecf1ec & lut_mask_in) : lut = 64'hdff118b8dea0fe1b;
      (64'hc7e04822c40fc40f & lut_mask_in) : lut = 64'ha7d77895800f79b5;
      (64'h2dac37c4e783e783 & lut_mask_in) : lut = 64'h2fde09d307ad9157;
      (64'hbb02b8e879a879a8 & lut_mask_in) : lut = 64'h9853c0dff3bfb1c0;
      (64'he02a7aac04ac04ac & lut_mask_in) : lut = 64'h2ee3d7977e87fe22;
      (64'h22fd55b6c86ec86e & lut_mask_in) : lut = 64'haecfe34811973e06;
      (64'hec54b430d34bd34b & lut_mask_in) : lut = 64'hce808d39a5c289a4;
      (64'h973f6b0af085f085 & lut_mask_in) : lut = 64'hc046ee92c19fb108;
      (64'h3c747212e746e746 & lut_mask_in) : lut = 64'h58de3ea7a9deee43;
      (64'hb2fd7ca6bff9bff9 & lut_mask_in) : lut = 64'hf00fb8176084164a;
      (64'h896e6f61b12ab12a & lut_mask_in) : lut = 64'h5692ff2a64e1ba00;
      (64'h2b72c8e4690f690f & lut_mask_in) : lut = 64'ha0db4a1c53337666;
      (64'h9a41a7647fb47fb4 & lut_mask_in) : lut = 64'h1981f5f212375238;
      (64'h276586411d371d37 & lut_mask_in) : lut = 64'hb3de7344f5f0861d;
      (64'hdd21d3201f4a1f4a & lut_mask_in) : lut = 64'hbd835d1f3007baf1;
      (64'h5372f63245d345d3 & lut_mask_in) : lut = 64'h7aa7b6ecde32a302;
      (64'he1cb8f8625532553 & lut_mask_in) : lut = 64'h97e61962fd04eeb2;
      (64'hb6b4a7397baf7baf & lut_mask_in) : lut = 64'hd87a47c1da4e01df;
      (64'hb2744b744cbb4cbb & lut_mask_in) : lut = 64'hf6109db1cba4f859;
      (64'hcabdb5b2be8fbe8f & lut_mask_in) : lut = 64'h93484e7bb1aa586e;
      (64'hd4a16dd5d47fd47f & lut_mask_in) : lut = 64'hbdf7b81e2074a171;
      (64'hcf6caed309f309f3 & lut_mask_in) : lut = 64'h3132b930af1dc338;
      (64'he15bf8d6566a566a & lut_mask_in) : lut = 64'hb3fe9e196d8e4d2f;
      (64'hdc9c0be8769c769c & lut_mask_in) : lut = 64'h4705bb3b88e685c5;
      (64'h0a5799ea00d000d0 & lut_mask_in) : lut = 64'h66f70063fde9da22;
      (64'hd14b17c268716871 & lut_mask_in) : lut = 64'hbeeea5ee57e5d2d0;
      (64'h49f8258512861286 & lut_mask_in) : lut = 64'h814f255f21444bac;
      (64'h9ae275b052f352f3 & lut_mask_in) : lut = 64'h9ce02c1e52399227;
      (64'h6978522208d208d2 & lut_mask_in) : lut = 64'h7e003356727c4d2f;
      (64'h781a536a2abe2abe & lut_mask_in) : lut = 64'h58b9bd1343b72982;
      (64'h749bf21d22952295 & lut_mask_in) : lut = 64'heaf70c842aa69dc9;
      (64'hd85527c08ab78ab7 & lut_mask_in) : lut = 64'hc2e6147f8bbcc2d2;
      (64'h2be69b8025322532 & lut_mask_in) : lut = 64'hbd1e6409b3542b5c;
      (64'hf6a319b209950995 & lut_mask_in) : lut = 64'h3f462df5b5de7ff1;
      (64'h2c65156344cb44cb & lut_mask_in) : lut = 64'h71b4f867bcf3c1f8;
      (64'h2f500f1898529852 & lut_mask_in) : lut = 64'h150ffe7202543c60;
      (64'h46e3c0c66b826b82 & lut_mask_in) : lut = 64'h7eb79ef7087afef3;
      (64'hc529601b44204420 & lut_mask_in) : lut = 64'h9816b01256730827;
      (64'hd2cbd786d0e7d0e7 & lut_mask_in) : lut = 64'hd125846025a92859;
      (64'h1a60ebe1f8adf8ad & lut_mask_in) : lut = 64'hbf4961e76d08aeb3;
      (64'he9b2819b53b253b2 & lut_mask_in) : lut = 64'h9f6cf6145bfbbf54;
      (64'hfed99880e18ee18e & lut_mask_in) : lut = 64'h8348b276558d7144;
      (64'h4fbb26e0410d410d & lut_mask_in) : lut = 64'h9b784c3aebca988f;
      (64'h6fc1e391cf44cf44 & lut_mask_in) : lut = 64'h17723d4fff41eb64;
      (64'hf67b7ec5a5d5a5d5 & lut_mask_in) : lut = 64'h5664a21ddda545b2;
      (64'hdeedcacb60d060d0 & lut_mask_in) : lut = 64'he5fb118ff7e5c257;
      (64'hd4bac6f0291d291d & lut_mask_in) : lut = 64'hcf6a38eb1b1d0f43;
      (64'h4592654738673867 & lut_mask_in) : lut = 64'h8a7a1d5476a4a81a;
      (64'h7f7b8545208d208d & lut_mask_in) : lut = 64'hfc7fc8dcc1dd726e;
      (64'h8d5d0ce43f313f31 & lut_mask_in) : lut = 64'h18746b8939751360;
      (64'hf5b9a478e2f5e2f5 & lut_mask_in) : lut = 64'h710fbeb5b0a7562d;
      (64'h3bd798b358c358c3 & lut_mask_in) : lut = 64'h90c72f49728bb0b9;
      (64'hf35115339f399f39 & lut_mask_in) : lut = 64'hafd6c9d409558331;
      (64'h80b20bdf8a018a01 & lut_mask_in) : lut = 64'h93a3689afa816706;
      (64'hda27ec5d58565856 & lut_mask_in) : lut = 64'h34bdde6a781d72f9;
      (64'h3e319c24a973a973 & lut_mask_in) : lut = 64'he6026a77eff31912;
      (64'h24bcc25fbd7dbd7d & lut_mask_in) : lut = 64'h2a591d7281edb557;
      (64'hfb1b4a9e92dd92dd & lut_mask_in) : lut = 64'h162feb314389b2e2;
      (64'h81db73adf7bbf7bb & lut_mask_in) : lut = 64'hb0c77262dda89181;
      (64'h8d51f72446fa46fa & lut_mask_in) : lut = 64'he2bb5b40c698e9d9;
      (64'h2851a374cef3cef3 & lut_mask_in) : lut = 64'h94c311ef701319bf;
      (64'h9b5bbb8ae987e987 & lut_mask_in) : lut = 64'hcaa12be5b09da298;
      (64'h857c3008d935d935 & lut_mask_in) : lut = 64'h3b95d537a18391ab;
      (64'h6da8ccfe26a226a2 & lut_mask_in) : lut = 64'h94ee4538fc9b3576;
      (64'he564a1938bac8bac & lut_mask_in) : lut = 64'h4fc8862aa34a0c6c;
      (64'h3046eec609180918 & lut_mask_in) : lut = 64'he793bbbe8cb861eb;
      (64'ha5e3704c44c044c0 & lut_mask_in) : lut = 64'ha708fd4c57acf100;
      (64'hb83e2db49f499f49 & lut_mask_in) : lut = 64'h000d00d28b6a0e09;
      (64'h392067bf94929492 & lut_mask_in) : lut = 64'h5c658ec9218ca19c;
      (64'hb79828d850b850b8 & lut_mask_in) : lut = 64'h9539232dd04f8ba4;
      (64'h5c1fda62886a886a & lut_mask_in) : lut = 64'h7d0fc4a6157535fb;
      (64'h1fd78876fe67fe67 & lut_mask_in) : lut = 64'hd96b53877e7190a2;
      (64'h3cf10f6b44104410 & lut_mask_in) : lut = 64'hba94bc75cb5e0414;
      (64'h211780f090899089 & lut_mask_in) : lut = 64'h0a3ef6ccdb7d8f5b;
      (64'hf577ac6c254a254a & lut_mask_in) : lut = 64'h9cb1ddbc38915b84;
      (64'he08d435628cf28cf & lut_mask_in) : lut = 64'hf4d3e5c1b34a6226;
      (64'h09fc61166a416a41 & lut_mask_in) : lut = 64'h3dbae4d49195a4f4;
      (64'h730c8d40f7d9f7d9 & lut_mask_in) : lut = 64'h99775aaf25df332a;
      (64'h6a80771204f704f7 & lut_mask_in) : lut = 64'hbfe6f8368d3e2650;
      (64'hf929bdc11e501e50 & lut_mask_in) : lut = 64'ha1fb285b4bdf2c44;
      (64'he20091812a612a61 & lut_mask_in) : lut = 64'h976551a2d7c79ee9;
      (64'hc4bc9df372417241 & lut_mask_in) : lut = 64'h970a0d7d99ac2299;
      (64'hf87d31fd47b447b4 & lut_mask_in) : lut = 64'ha8a21f637c6605bc;
      (64'hef5e5326831b831b & lut_mask_in) : lut = 64'h6c3b1c62e6af15df;
      (64'h1ee8c15e67966796 & lut_mask_in) : lut = 64'h50a07f409cd536e7;
      (64'h8ff363dab8e2b8e2 & lut_mask_in) : lut = 64'hb8b988c29471b73b;
      (64'h32c2a90b1e921e92 & lut_mask_in) : lut = 64'hc4d5fca9e1756c09;
      (64'h47068d2f3efd3efd & lut_mask_in) : lut = 64'h0835058b65980242;
      (64'h93e3fc89546b546b & lut_mask_in) : lut = 64'h36f4e6a869c4211e;
      (64'h6e5a0d883f703f70 & lut_mask_in) : lut = 64'h62e6862ac517fda6;
      (64'h6b40ef4cdc63dc63 & lut_mask_in) : lut = 64'hc1dcd2aeae915d07;
      (64'hd0a47ca712e512e5 & lut_mask_in) : lut = 64'he491bdb555f6d8a9;
      (64'hcc1207f299aa99aa & lut_mask_in) : lut = 64'h2b3e739cfb1aeca3;
      (64'h74f325a5a776a776 & lut_mask_in) : lut = 64'ha3a4da348ea42136;
      (64'h277996474a8d4a8d & lut_mask_in) : lut = 64'hf4353266dd139617;
      (64'h6c83fc0b81658165 & lut_mask_in) : lut = 64'h7e3b736f0a8411de;
      (64'h9cb1720c21472147 & lut_mask_in) : lut = 64'hc08ed6ac7def42df;
      (64'h6074d408ea97ea97 & lut_mask_in) : lut = 64'ha795ba1438a4830e;
      (64'h41854e0d6d626d62 & lut_mask_in) : lut = 64'hc985d9a876979948;
      (64'hd23a5198d4acd4ac & lut_mask_in) : lut = 64'he840b5ddf9b8e567;
      (64'hd19bea7d83908390 & lut_mask_in) : lut = 64'h3db8edd540b446d4;
      (64'ha8600fd291959195 & lut_mask_in) : lut = 64'he0eafe7dd0a848c6;
      (64'hc4f048b202570257 & lut_mask_in) : lut = 64'h3501349d09a57a3c;
      (64'h9ef2fc98dcd0dcd0 & lut_mask_in) : lut = 64'hb20c8588f20a42be;
      (64'h4a983709e83ee83e & lut_mask_in) : lut = 64'h8b8a066f1fbe542c;
      (64'heb572f5a54185418 & lut_mask_in) : lut = 64'h4108d436a856c3e0;
      (64'h5318785232a232a2 & lut_mask_in) : lut = 64'he21c73ca047c6a49;
      (64'h9ceb9eb1463e463e & lut_mask_in) : lut = 64'hd83c7d0c3d2d2e52;
      (64'h083352d8990f990f & lut_mask_in) : lut = 64'h1c20a31e2f848bad;
      (64'h7671a7c1d267d267 & lut_mask_in) : lut = 64'h7429e750a91213a0;
      (64'h2e763c4e81f781f7 & lut_mask_in) : lut = 64'h3320ec4701ac7cde;
      (64'h204aa639c074c074 & lut_mask_in) : lut = 64'h1d9d4764a89a1115;
      (64'h55e5469609150915 & lut_mask_in) : lut = 64'h6130a2506d114bd8;
      (64'hcdce9fb342174217 & lut_mask_in) : lut = 64'hedb96a419a7caf5b;
      (64'h8894188bf654f654 & lut_mask_in) : lut = 64'hb39b70ff4ed4b06b;
      (64'he0fdbe552d7b2d7b & lut_mask_in) : lut = 64'hb7cdae14a49e3f30;
      (64'hd3431950ed6ced6c & lut_mask_in) : lut = 64'h56de607bfe77f73d;
      (64'h86573e13883e883e & lut_mask_in) : lut = 64'h23ea796a3153ca8e;
      (64'h206af197aed6aed6 & lut_mask_in) : lut = 64'ha81d6384fc5d19d1;
      (64'h931249657c9c7c9c & lut_mask_in) : lut = 64'hc389489fed8faa2e;
      (64'h906e6166b824b824 & lut_mask_in) : lut = 64'h7bdf22c065662cdd;
      (64'h0f74781e5bac5bac & lut_mask_in) : lut = 64'h1bdc29dfce49b994;
      (64'he1422eaea860a860 & lut_mask_in) : lut = 64'h4e22afd337d5ca92;
      (64'hd2a5be1e3df43df4 & lut_mask_in) : lut = 64'hc047ec3dd1865a37;
      (64'h6673af4382d282d2 & lut_mask_in) : lut = 64'h5c56f4c7d6ac1e04;
      (64'h3a463ac0b9b1b9b1 & lut_mask_in) : lut = 64'he9eadf5fe5e7cc9f;
      (64'h5e7d1de32af92af9 & lut_mask_in) : lut = 64'h70d7e620701e71e4;
      (64'h881a4c7857445744 & lut_mask_in) : lut = 64'h28ada2dc5d177bf2;
      (64'h01e7973863c263c2 & lut_mask_in) : lut = 64'h75db94c2c19aedcf;
      (64'hae99b8fc6fc26fc2 & lut_mask_in) : lut = 64'hf9d3641a86e5d69b;
      (64'ha3d99b482b0f2b0f & lut_mask_in) : lut = 64'hd376ee6ba1700312;
      (64'hd02c02a501430143 & lut_mask_in) : lut = 64'h6f50d6beb1df0397;
      (64'he2e71f7fdd8cdd8c & lut_mask_in) : lut = 64'h3f8ebaf9ea9caed4;
      (64'hd7f59b0e13531353 & lut_mask_in) : lut = 64'h7aed7ee746973f89;
      (64'hd3886672c5c1c5c1 & lut_mask_in) : lut = 64'h0257aa850fbe86d5;
      (64'hc649c3540c400c40 & lut_mask_in) : lut = 64'h46cae6b8fda310cc;
      (64'hd0b581d9418e418e & lut_mask_in) : lut = 64'h4e923f3b4d611db4;
      (64'hdb6a5417d42ad42a & lut_mask_in) : lut = 64'h9df852af57b54d8c;
      (64'h22e33d4b507f507f & lut_mask_in) : lut = 64'hb2d10fab82a89921;
      (64'hee33d16f02200220 & lut_mask_in) : lut = 64'h8de45716e9e38739;
      (64'hc67b8c47b89fb89f & lut_mask_in) : lut = 64'h994143d224b6cd34;
      (64'hf2158f02e260e260 & lut_mask_in) : lut = 64'h351d1e7bae676e7c;
      (64'hdf2d3ea52d082d08 & lut_mask_in) : lut = 64'ha0b722fffccd0361;
      (64'h7eaa5b6999d399d3 & lut_mask_in) : lut = 64'hdc836a2dc0a0defd;
      (64'h55822a6cf8f1f8f1 & lut_mask_in) : lut = 64'h61ef00a1f6a5e8c9;
      (64'h585ab599b60bb60b & lut_mask_in) : lut = 64'h38066ef3ec05b924;
      (64'hc4d42db18fee8fee & lut_mask_in) : lut = 64'h936523d94c6365bc;
      (64'hb9c6d5b276c476c4 & lut_mask_in) : lut = 64'h4f5ec87cbb3dad8f;
      (64'he803bebe3dff3dff & lut_mask_in) : lut = 64'hf91b54cbb4ca585e;
      (64'hcf1d97bc37f237f2 & lut_mask_in) : lut = 64'h209010874b987b08;
      (64'h7672df7417751775 & lut_mask_in) : lut = 64'habe20ec1965e75fa;
      (64'h7335b6b612cf12cf & lut_mask_in) : lut = 64'h679339951e25d05b;
      (64'h3cacffd2e537e537 & lut_mask_in) : lut = 64'h09ed9a86bbff7e5f;
      (64'h395ea81daec5aec5 & lut_mask_in) : lut = 64'hadb52f8093eb675b;
      (64'h12114f2c25ea25ea & lut_mask_in) : lut = 64'h80acc9a17bb95347;
      (64'h93d1ac1c34c534c5 & lut_mask_in) : lut = 64'ha3bfbbe415d6849f;
      (64'h3d9587f2932a932a & lut_mask_in) : lut = 64'h7670b922522b3577;
      (64'h40f2be62c718c718 & lut_mask_in) : lut = 64'h580d1ee5b9a9eb67;
      (64'h073eed7225ed25ed & lut_mask_in) : lut = 64'h09842b80c17993fc;
      (64'hc0ebd0abeec4eec4 & lut_mask_in) : lut = 64'hcef98dd57dc3b33d;
      (64'h8e637e769f529f52 & lut_mask_in) : lut = 64'h73ec0609f2a44699;
      (64'he445ab20e2f7e2f7 & lut_mask_in) : lut = 64'hadb0fcbc4addad43;
      (64'hd4832dd8040e040e & lut_mask_in) : lut = 64'hd353675446c11dc8;
      (64'h670a019e504a504a & lut_mask_in) : lut = 64'h3da3951b04d600de;
      (64'hb776a80842af42af & lut_mask_in) : lut = 64'hc678b636d883de1b;
      (64'ha20d12af2df02df0 & lut_mask_in) : lut = 64'hf0b097b8908b2ffd;
      (64'hc53cd02310691069 & lut_mask_in) : lut = 64'hcdfb1e6af8eb0529;
      (64'h7f334b586fd76fd7 & lut_mask_in) : lut = 64'hd507b48630342033;
      (64'h1308ca819b299b29 & lut_mask_in) : lut = 64'h593a6299c1768ed6;
      (64'h876700add3ebd3eb & lut_mask_in) : lut = 64'h01ba3fcecbf887ec;
      (64'h186f67ce0b4f0b4f & lut_mask_in) : lut = 64'hcdb7a2ac828b5f38;
      (64'h43a3e8f1715e715e & lut_mask_in) : lut = 64'h34f0bfec5f4983be;
      (64'h11e89ba309f109f1 & lut_mask_in) : lut = 64'h189eb6059e25a953;
      (64'hfc85692cd4efd4ef & lut_mask_in) : lut = 64'h5b53fb5888cf7ff8;
      (64'h4eb6b514b3c4b3c4 & lut_mask_in) : lut = 64'h3a032508d0b1ba92;
      (64'h074bc7fe40ed40ed & lut_mask_in) : lut = 64'hb0c7442c4cbddb76;
      (64'h56c3174baf3faf3f & lut_mask_in) : lut = 64'h8614ac1cbc041cb1;
      (64'he64c903e74f674f6 & lut_mask_in) : lut = 64'ha7d720be7467c51e;
      (64'h62b13bc6de1ede1e & lut_mask_in) : lut = 64'h53061b0ac9f588b3;
      (64'h2389dbcbbaa5baa5 & lut_mask_in) : lut = 64'hf27a241d45cbf769;
      (64'h0def3da8db13db13 & lut_mask_in) : lut = 64'h9654cfe46ca1f82d;
      (64'he3548cadecf2ecf2 & lut_mask_in) : lut = 64'h7c7c6e1a4d08a1b8;
      (64'h4ec1e241142a142a & lut_mask_in) : lut = 64'he397f76423ac8f36;
      (64'hbfc3f859f0a6f0a6 & lut_mask_in) : lut = 64'h8c3ad4eebb9bdc27;
      (64'hd0435af93c273c27 & lut_mask_in) : lut = 64'h6e2691ceb4cbff1c;
      (64'h2a0987c74d614d61 & lut_mask_in) : lut = 64'h3c989ec3d24cc696;
      (64'hcbca20b3567a567a & lut_mask_in) : lut = 64'h6d40c88c55d77b8c;
      (64'h59c2ac8968886888 & lut_mask_in) : lut = 64'hd14c9d6a8904fbd9;
      (64'h2723dd5ddc86dc86 & lut_mask_in) : lut = 64'h8c063b4a74c16be0;
      (64'hb5dd14601dad1dad & lut_mask_in) : lut = 64'h5efd5d7b88580009;
      (64'h699943f077ea77ea & lut_mask_in) : lut = 64'hf55543c08b31c139;
      (64'h8159c072b504b504 & lut_mask_in) : lut = 64'h14037740b95c1963;
      (64'h992fec5422772277 & lut_mask_in) : lut = 64'ha05903ae89aa1e1f;
      (64'ha9e646b36fb36fb3 & lut_mask_in) : lut = 64'ha79b193be9d66389;
      (64'h8f54de4c71797179 & lut_mask_in) : lut = 64'h438bc2e10006dfbd;
      (64'ha02d6bf4fd41fd41 & lut_mask_in) : lut = 64'hb744eba19346f069;
      (64'h4a0fdcf8c775c775 & lut_mask_in) : lut = 64'h1b95710575da4eb9;
      (64'hbb4401a0ebd0ebd0 & lut_mask_in) : lut = 64'h2d58dba8665a7517;
      (64'h54c80b2fcddbcddb & lut_mask_in) : lut = 64'h0d5665a46dc44dbf;
      (64'hec5bc76d147a147a & lut_mask_in) : lut = 64'h0bfe9985ee6e7ec9;
      (64'h6a066bf4831a831a & lut_mask_in) : lut = 64'h9da2fbbad48bde07;
      (64'hd0800da134103410 & lut_mask_in) : lut = 64'h32757f201dcda17d;
      (64'h3b29bd743a5d3a5d & lut_mask_in) : lut = 64'h05d1a6a27e0113b3;
      (64'hc1a3fc1cba83ba83 & lut_mask_in) : lut = 64'hc7c7fdae090cc230;
      (64'h921bdf330ed20ed2 & lut_mask_in) : lut = 64'hd50d21c4657230f2;
      (64'h2c4e57ef38623862 & lut_mask_in) : lut = 64'h87d928ef8360f0de;
      (64'h7decdde7b65bb65b & lut_mask_in) : lut = 64'h7a267d0359571fe6;
      (64'he3715a7d1bcc1bcc & lut_mask_in) : lut = 64'hd4c92b68e65220f9;
      (64'h39600158114f114f & lut_mask_in) : lut = 64'h736555a3fb21de14;
      (64'hb754f6f67e417e41 & lut_mask_in) : lut = 64'haa342ce94a7c0047;
      (64'h1d2b78ae06bd06bd & lut_mask_in) : lut = 64'h8de6a817b0b6335b;
      (64'h677f28b089098909 & lut_mask_in) : lut = 64'hddd245a71fe6e2fc;
      (64'h32d924c5b6a4b6a4 & lut_mask_in) : lut = 64'hf74b979d6ab86282;
      (64'hc73562aadb2bdb2b & lut_mask_in) : lut = 64'h982a15a390148c98;
      (64'h99d41551e501e501 & lut_mask_in) : lut = 64'h5118772159db54c5;
      (64'h8e5407bba94da94d & lut_mask_in) : lut = 64'h870a6883cd1a3d90;
      (64'h18e8d0b83aa93aa9 & lut_mask_in) : lut = 64'h26e566dc496460ec;
      (64'hb5b9bdad396e396e & lut_mask_in) : lut = 64'h58ae7a49d3bab8d1;
      (64'h33ca0aa68e188e18 & lut_mask_in) : lut = 64'hdb52faa2070d2085;
      (64'hcc921f1109050905 & lut_mask_in) : lut = 64'hd9b86e1f506e86ca;
      (64'h5c32f8fb29372937 & lut_mask_in) : lut = 64'h24594de1bb20f255;
      (64'h8c07856c02660266 & lut_mask_in) : lut = 64'h748f42c036844f2d;
      (64'h9aad8d0280938093 & lut_mask_in) : lut = 64'hd8746ccc69befa53;
      (64'h4f37aac85f715f71 & lut_mask_in) : lut = 64'he521250a2982c0f1;
      (64'h03220772276f276f & lut_mask_in) : lut = 64'ha14de9dc59e9ca02;
      (64'h01cde3ce04250425 & lut_mask_in) : lut = 64'hc7f377657f126da1;
      (64'he5c043814d054d05 & lut_mask_in) : lut = 64'h093f9b5d4f65dfd9;
      (64'h9c32074ab881b881 & lut_mask_in) : lut = 64'he662e534845cbb25;
      (64'h959043c24bb74bb7 & lut_mask_in) : lut = 64'hb7e5b9e6879a3928;
      (64'h609449f015901590 & lut_mask_in) : lut = 64'h59725008f848c56b;
      (64'h6b014cc6a2b9a2b9 & lut_mask_in) : lut = 64'hbe3d1a3526a81c8f;
      (64'h8df7bee022a422a4 & lut_mask_in) : lut = 64'h3aaa25ea2a6c714f;
      (64'hc4c18f1d55e855e8 & lut_mask_in) : lut = 64'h4ab7ccdf557a7f30;
      (64'hcdbc3c60fbc6fbc6 & lut_mask_in) : lut = 64'h230d2fe4714b2082;
      (64'h1ca85137a0b0a0b0 & lut_mask_in) : lut = 64'hd733afd9f6df6c11;
      (64'h7f535a2294ef94ef & lut_mask_in) : lut = 64'h26ee363a39e62b7d;
      (64'h7c7c148afd34fd34 & lut_mask_in) : lut = 64'h77562340cf65e88a;
      (64'h8b87b97461d661d6 & lut_mask_in) : lut = 64'hee04222dab388085;
      (64'h70007e8964206420 & lut_mask_in) : lut = 64'hd895a6f73b4e4340;
      (64'h92604b44a02da02d & lut_mask_in) : lut = 64'h8a6b0302c80debff;
      (64'h15e6a6a2090f090f & lut_mask_in) : lut = 64'h0672e26f3ea5b504;
      (64'h5c475b7cc0cfc0cf & lut_mask_in) : lut = 64'h624a094f9a8a70a9;
      (64'h28fcf7bb608a608a & lut_mask_in) : lut = 64'h287c508c4193d1ba;
      (64'hd31ef20f07a107a1 & lut_mask_in) : lut = 64'h79bc29933bfc57b5;
      (64'hd0072bf0f739f739 & lut_mask_in) : lut = 64'hb5e57b7effa87bdd;
      (64'h10f1ecdeecdaecda & lut_mask_in) : lut = 64'hc631d153abfe681e;
      (64'h0206be0f0ce60ce6 & lut_mask_in) : lut = 64'h066a3592c83dea4e;
      (64'hbcbc1fc1daa7daa7 & lut_mask_in) : lut = 64'h30c693d733b8e7c4;
      (64'h531250e625572557 & lut_mask_in) : lut = 64'h8090296c4a97cc00;
      (64'h53c4aca4b323b323 & lut_mask_in) : lut = 64'hb89af962fcb587ca;
      (64'hb632ae79d952d952 & lut_mask_in) : lut = 64'h5a361b8b8997afa9;
      (64'hab93bdcc977a977a & lut_mask_in) : lut = 64'h06b23dbf5b554e34;
      (64'h2ce0971afe3afe3a & lut_mask_in) : lut = 64'h1b35e1f64efd5438;
      (64'h70e361deb4b7b4b7 & lut_mask_in) : lut = 64'ha40f8fa528b17a1d;
      (64'hb413f1ad8b078b07 & lut_mask_in) : lut = 64'h79dbe0efa5d774d6;
      (64'hf7ef28848c858c85 & lut_mask_in) : lut = 64'h4e1ea969736094a3;
      (64'h378dd3b985fe85fe & lut_mask_in) : lut = 64'hb7447bd456eb15f4;
      (64'h0458ef5a08c608c6 & lut_mask_in) : lut = 64'hd6de0c511dde3b12;
      (64'ha2ec97fa15421542 & lut_mask_in) : lut = 64'h4d8c1b2945bf5297;
      (64'h7ee851dcb8d3b8d3 & lut_mask_in) : lut = 64'hacde8580e5fac2c0;
      (64'h224b3bf44f3b4f3b & lut_mask_in) : lut = 64'hdf0adf15625d82f7;
      (64'h75712820bae2bae2 & lut_mask_in) : lut = 64'h56985c85e1ff8d9f;
      (64'h382256275ea35ea3 & lut_mask_in) : lut = 64'h6afb4fd28e4c5fe4;
      (64'h8a7890f8272d272d & lut_mask_in) : lut = 64'hf065fc541bf3da9b;
      (64'h0af6abdc0a540a54 & lut_mask_in) : lut = 64'h15659b9bdb0aca3a;
      (64'h357eb68e358d358d & lut_mask_in) : lut = 64'hd3dc797c1b8403a8;
      (64'hb5cb3d8cf3a7f3a7 & lut_mask_in) : lut = 64'h25d63c2a9ca94059;
      (64'hfc23277e8ed48ed4 & lut_mask_in) : lut = 64'h3820f16d283d964b;
      (64'h45a3f6930bb80bb8 & lut_mask_in) : lut = 64'hf386a80d7945eb04;
      (64'h95d8f42475fa75fa & lut_mask_in) : lut = 64'hebd5e276ce96c524;
      (64'h929818b6a258a258 & lut_mask_in) : lut = 64'h8dc6bee8649665a1;
      (64'h8b96c54663f963f9 & lut_mask_in) : lut = 64'h50d7aee59eb55305;
      (64'h99cb7d1fae17ae17 & lut_mask_in) : lut = 64'he6bd25e9e5c519bd;
      (64'h379c929786328632 & lut_mask_in) : lut = 64'ha3d2d1a43f4119f9;
      (64'hc1ab458f55245524 & lut_mask_in) : lut = 64'hd45c5acbec8dc6ba;
      (64'ha8522049c07dc07d & lut_mask_in) : lut = 64'hf14337b33013cf8c;
      (64'h6d6865c859b859b8 & lut_mask_in) : lut = 64'h113428519565f29e;
      (64'h2b418f887a6b7a6b & lut_mask_in) : lut = 64'h0971f7030359e59e;
      (64'ha6ce02c03d0e3d0e & lut_mask_in) : lut = 64'h5531bae2ef4d42d2;
      (64'hdf5a372697eb97eb & lut_mask_in) : lut = 64'h53129a7005109753;
      (64'h1c36f8b090919091 & lut_mask_in) : lut = 64'hfe2f83cc3c182ed3;
      (64'h62c3d0453ec63ec6 & lut_mask_in) : lut = 64'hc6434fd71c88004e;
      (64'ha241898946944694 & lut_mask_in) : lut = 64'h5edd0ea8c9178412;
      (64'h34be0217a1e6a1e6 & lut_mask_in) : lut = 64'ha1812012ce02d92f;
      (64'hed923c3d34573457 & lut_mask_in) : lut = 64'hcbc6d4fb1d65114e;
      (64'h395a45d75ae85ae8 & lut_mask_in) : lut = 64'ha3bd83b04a14500c;
      (64'ha096d3b76c696c69 & lut_mask_in) : lut = 64'hc5241d12fd5df9fb;
      (64'h4c9acc56a2f6a2f6 & lut_mask_in) : lut = 64'hb98ccecc7db821ce;
      (64'h0f3c9bdec4b9c4b9 & lut_mask_in) : lut = 64'h8a0441850b90621b;
      (64'he4ad46df68e268e2 & lut_mask_in) : lut = 64'h769392372a4654f3;
      (64'h26aeb487d628d628 & lut_mask_in) : lut = 64'h26d662ac037e7b68;
      (64'h9ad6d90bf913f913 & lut_mask_in) : lut = 64'h0a590157931b748f;
      (64'h2b208b4879847984 & lut_mask_in) : lut = 64'h882dc60ddef55b76;
      (64'h86675e08de74de74 & lut_mask_in) : lut = 64'h86bc3fef7cd3ff9c;
      (64'he46ac234c491c491 & lut_mask_in) : lut = 64'h416b798d01d11038;
      (64'h4fb1085244cc44cc & lut_mask_in) : lut = 64'hd0c7de61fee6079d;
      (64'he8afd6e7ccc4ccc4 & lut_mask_in) : lut = 64'ha350bdb00b8a75d5;
      (64'h8751ffbf6beb6beb & lut_mask_in) : lut = 64'hf0ea190604380b80;
      (64'hb6689ee03c453c45 & lut_mask_in) : lut = 64'hfe6397a9112c99f6;
      (64'h023a39c6fbb4fbb4 & lut_mask_in) : lut = 64'h5259dab36dd565dc;
      (64'he3445dd327622762 & lut_mask_in) : lut = 64'h66cb670859248f3e;
      (64'hc70ea1a695699569 & lut_mask_in) : lut = 64'h16ee894852b39644;
      (64'h238c785d461e461e & lut_mask_in) : lut = 64'h1f12fe9d6135f4f6;
      (64'h56e7ef4b89bf89bf & lut_mask_in) : lut = 64'hf924c5b1c1167733;
      (64'h07a6bcc83bfd3bfd & lut_mask_in) : lut = 64'h0bb5000066c84bd8;
      (64'h835bd69f8b898b89 & lut_mask_in) : lut = 64'hf9ccd1020645cf5d;
      (64'h7cccf6dae256e256 & lut_mask_in) : lut = 64'hfe11fd1b91d447ac;
      (64'h7bb612f0bcffbcff & lut_mask_in) : lut = 64'h1081fef3de3f18fe;
      (64'h349db1600d5a0d5a & lut_mask_in) : lut = 64'hd87166bc91872fbe;
      (64'h88e7e6119aeb9aeb & lut_mask_in) : lut = 64'hd343758284282805;
      (64'h09a90c2bca03ca03 & lut_mask_in) : lut = 64'hc5bd876f660b6e19;
      (64'h9d0f3823ae8eae8e & lut_mask_in) : lut = 64'hf33501a4f139678f;
      (64'h20465d671f3b1f3b & lut_mask_in) : lut = 64'hfd601cf8e7a9d957;
      (64'h2977d31d71987198 & lut_mask_in) : lut = 64'he75fd49acaa35798;
      (64'hb1b03c0df0cdf0cd & lut_mask_in) : lut = 64'hb283ff9d5244cd0e;
      (64'hb9fdefb25b775b77 & lut_mask_in) : lut = 64'h9d594b31ec53bf5e;
      (64'hae9a557104150415 & lut_mask_in) : lut = 64'h8b0a4f94a20a1037;
      (64'h5f9e4350098d098d & lut_mask_in) : lut = 64'h0d05bdaa071faf93;
      (64'h9795d87724982498 & lut_mask_in) : lut = 64'he78c056fbf28c2b8;
      (64'h3b77ae68b213b213 & lut_mask_in) : lut = 64'h0629b45fd4d0087b;
      (64'haf22737b2b4e2b4e & lut_mask_in) : lut = 64'h9cb2c3200f1315b4;
      (64'h28d2a13317de17de & lut_mask_in) : lut = 64'hc19dfa1d8aaffb45;
      (64'h7e46534f2d632d63 & lut_mask_in) : lut = 64'hdbfc32fe0fbc5286;
      (64'h15699dc5ef20ef20 & lut_mask_in) : lut = 64'h3e7d5c4e8ae7c542;
      (64'hd756b8b6359c359c & lut_mask_in) : lut = 64'hd6a958eb7ad18858;
      (64'h885cf7bccd5fcd5f & lut_mask_in) : lut = 64'h027ce54017888b4b;
      (64'h562a4755544e544e & lut_mask_in) : lut = 64'hb55b487375de04c2;
      (64'h164177f7f6c9f6c9 & lut_mask_in) : lut = 64'h1b165495fc80412d;
      (64'h2f5063c50fbb0fbb & lut_mask_in) : lut = 64'h6b15f225ac975d55;
      (64'hefc23dc7d89fd89f & lut_mask_in) : lut = 64'h42295e17adc8d531;
      (64'ha66a99e1d8eed8ee & lut_mask_in) : lut = 64'ha1f0140603ac94b1;
      (64'h736c93ff09c909c9 & lut_mask_in) : lut = 64'h8a94be6fa294f62f;
      (64'hda59ff8aab60ab60 & lut_mask_in) : lut = 64'h0f6b1ce9e09b4817;
      (64'hcc0547994de64de6 & lut_mask_in) : lut = 64'h5dd50cefc13e9d5e;
      (64'h1ecb681863746374 & lut_mask_in) : lut = 64'hf7f7456587bfb6d9;
      (64'h47f6b1ca69c569c5 & lut_mask_in) : lut = 64'h37a62076df06a309;
      (64'hfbeda5fe0d110d11 & lut_mask_in) : lut = 64'h4d284fe5873fb9ca;
      (64'he7cba5990ea10ea1 & lut_mask_in) : lut = 64'he2be5b92be24d268;
      (64'h17eb5b3184a284a2 & lut_mask_in) : lut = 64'habd48e1bdd8d65da;
      (64'h40e20d9eabe0abe0 & lut_mask_in) : lut = 64'he8a4ff199241dee1;
      (64'h06a586d1344c344c & lut_mask_in) : lut = 64'h35d6edf0d8b7600c;
      (64'h5454b329a7c8a7c8 & lut_mask_in) : lut = 64'h1f128d27da149858;
      (64'hf4160ee576a676a6 & lut_mask_in) : lut = 64'h65c293bd9589df6d;
      (64'h158eb9a194a794a7 & lut_mask_in) : lut = 64'h47e0984260bb28c0;
      (64'hc8d0d2e567cb67cb & lut_mask_in) : lut = 64'h643e2f3d74b901c6;
      (64'hb927322759e559e5 & lut_mask_in) : lut = 64'hd63b540b594fde67;
      (64'h3435d174dd7fdd7f & lut_mask_in) : lut = 64'h3e1623437a5f9161;
      (64'h97cf45e4eebeeebe & lut_mask_in) : lut = 64'hc174e2812dc59859;
      (64'ha416dfcb17311731 & lut_mask_in) : lut = 64'h9bbec19ea343cc48;
      (64'hf74ad8ee92e292e2 & lut_mask_in) : lut = 64'h5f8eabfccce42e58;
      (64'hb1b766a074117411 & lut_mask_in) : lut = 64'hc7dd2f4eba498f67;
      (64'h4713b12e3a243a24 & lut_mask_in) : lut = 64'h35d824b2bd68337e;
      (64'h7f4003631f501f50 & lut_mask_in) : lut = 64'he771265e94404c8c;
      (64'hbbbadda2ece8ece8 & lut_mask_in) : lut = 64'h6324269a7de4f051;
      (64'h7489120a95fe95fe & lut_mask_in) : lut = 64'h8a0b6df729a6ec66;
      (64'h5920efcc64686468 & lut_mask_in) : lut = 64'hdc319384e54a65d6;
      (64'h884541b712781278 & lut_mask_in) : lut = 64'h9c9f30c839d26b3c;
      (64'he669cb929a859a85 & lut_mask_in) : lut = 64'hb9c4108d197bf91d;
      (64'h89c004e9c8d9c8d9 & lut_mask_in) : lut = 64'h044d10196f67b484;
      (64'h44c75d584f314f31 & lut_mask_in) : lut = 64'hef984e2b32d58e67;
      (64'h3019f8fb29c929c9 & lut_mask_in) : lut = 64'h77c6df9b9d09ee72;
      (64'h245c72cd728c728c & lut_mask_in) : lut = 64'hf5459ad4940f2cfc;
      (64'he34db7444c454c45 & lut_mask_in) : lut = 64'h84cb40e1c6a4148b;
      (64'hb6e13cdc64246424 & lut_mask_in) : lut = 64'h1badf6cdb69c9f74;
      (64'hb9a30d62ab5eab5e & lut_mask_in) : lut = 64'he676cfa34bc29d16;
      (64'hc18162d5c884c884 & lut_mask_in) : lut = 64'h5ad8d1e62b1e362a;
      (64'h27bd281785f885f8 & lut_mask_in) : lut = 64'hf510de3b917d0939;
      (64'h93cf144880038003 & lut_mask_in) : lut = 64'h405d26d83ea61f59;
      (64'h82b5bed855f855f8 & lut_mask_in) : lut = 64'h8a7453e7bf023ea1;
      (64'h5078dd3b24d324d3 & lut_mask_in) : lut = 64'h9699cba035711d3b;
      (64'he87756f1bf89bf89 & lut_mask_in) : lut = 64'hbca481a214c81132;
      (64'hfae7d010c529c529 & lut_mask_in) : lut = 64'h2aad0134d2848099;
      (64'h79a9f97924bc24bc & lut_mask_in) : lut = 64'h4398cfe61f9e49eb;
      (64'ha2e2effcdb14db14 & lut_mask_in) : lut = 64'he799054002f8b1f3;
      (64'hdc5e1ac2273f273f & lut_mask_in) : lut = 64'hc5ac181f6625cd12;
      (64'h1c7dc427b266b266 & lut_mask_in) : lut = 64'h554f9227bb48552b;
      (64'h0027df404c9f4c9f & lut_mask_in) : lut = 64'hf165b7b5680319c7;
      (64'h49b754c07ec37ec3 & lut_mask_in) : lut = 64'hc83895317223b006;
      (64'hbb2003a24bce4bce & lut_mask_in) : lut = 64'h02977ab1b25b36b9;
      (64'h43830d83d4c7d4c7 & lut_mask_in) : lut = 64'h7d30904c754378d7;
      (64'h7aae13cb5c105c10 & lut_mask_in) : lut = 64'h8141b43e39fb4beb;
      (64'h2dc6f01d25552555 & lut_mask_in) : lut = 64'h9b414f0843ff3e41;
      (64'h6f8ecedef648f648 & lut_mask_in) : lut = 64'h5b96de21dc3f1208;
      (64'h6f2de44518d418d4 & lut_mask_in) : lut = 64'h415291cd88ae1163;
      (64'h402f81003bea3bea & lut_mask_in) : lut = 64'ha913a099aff3f00c;
      (64'h37e13563a1b3a1b3 & lut_mask_in) : lut = 64'h687a5c8adc1ea9ec;
      (64'h3333285610ed10ed & lut_mask_in) : lut = 64'h469a602d3d2978be;
      (64'h52595623733e733e & lut_mask_in) : lut = 64'h68b2a53db1529198;
      (64'h1684933b1f961f96 & lut_mask_in) : lut = 64'hda50ed43f68637a0;
      (64'h4a09d8b0bc36bc36 & lut_mask_in) : lut = 64'h4d925a217298c8a3;
      (64'h08e9d2d2ee40ee40 & lut_mask_in) : lut = 64'h463de2be79de0302;
      (64'h859456f7d0efd0ef & lut_mask_in) : lut = 64'h037993bb57b2d7fd;
      (64'h1c0901e31f4c1f4c & lut_mask_in) : lut = 64'h75c7553af2c09e49;
      (64'h384e6faeefbdefbd & lut_mask_in) : lut = 64'h8e38b1ea60c7b654;
      (64'h1bfa39f99a3f9a3f & lut_mask_in) : lut = 64'hffa9afa371d6e565;
      (64'h0310ce2ddbfcdbfc & lut_mask_in) : lut = 64'hadf7a523a3cb3ee6;
      (64'h29cf414180088008 & lut_mask_in) : lut = 64'h0e99476cea12f24e;
      (64'hbf357cb6ab12ab12 & lut_mask_in) : lut = 64'he40ae5eb67a260f8;
      (64'ha2d05fe4521c521c & lut_mask_in) : lut = 64'h8b6daf5b0f8f2090;
      (64'hcc8bc6eccc76cc76 & lut_mask_in) : lut = 64'hb879fdec4144e1a9;
      (64'h1c1c181d7f187f18 & lut_mask_in) : lut = 64'h1b85503a7a2d9778;
      (64'he67cd6053b9f3b9f & lut_mask_in) : lut = 64'h3df21b31776bdf4a;
      (64'h83c6fd9970347034 & lut_mask_in) : lut = 64'h66ffa16ac6bc7572;
      (64'heea313dc73c173c1 & lut_mask_in) : lut = 64'h03b2f3cc79b716bb;
      (64'h0f5cb551bc6dbc6d & lut_mask_in) : lut = 64'h0438a8052edc8b1d;
      (64'h20771a3bd546d546 & lut_mask_in) : lut = 64'he16953c9d1e67eb9;
      (64'hab96e9cd06a806a8 & lut_mask_in) : lut = 64'h1e214422b19f2980;
      (64'h2253186f242c242c & lut_mask_in) : lut = 64'hfb86976bc46c8ce7;
      (64'ha3fb37fcf2f7f2f7 & lut_mask_in) : lut = 64'h722126a236f9f53f;
      (64'h4cfaedc160fb60fb & lut_mask_in) : lut = 64'h7f186374cc4fd541;
      (64'hf6ef01fa03580358 & lut_mask_in) : lut = 64'h59ec9640e9c1ee73;
      (64'h55139ee3c07fc07f & lut_mask_in) : lut = 64'he5920380f6b95789;
      (64'h90e20aa3bedbbedb & lut_mask_in) : lut = 64'h9e410dda451f0d74;
      (64'hb208fce33d7a3d7a & lut_mask_in) : lut = 64'h10456b9114fe64e5;
      (64'h3ad34426327f327f & lut_mask_in) : lut = 64'h53ef70dfdf51f51b;
      (64'hc98998d846364636 & lut_mask_in) : lut = 64'hf1432522436a8029;
      (64'h77789eccb16bb16b & lut_mask_in) : lut = 64'hc51294feee8573e9;
      (64'hf17f43241a4b1a4b & lut_mask_in) : lut = 64'h8c96e667a256f499;
      (64'h6f81f5ec3d513d51 & lut_mask_in) : lut = 64'h6472f4f6155e90b7;
      (64'hef67b0f2d03fd03f & lut_mask_in) : lut = 64'hd34d85cbd2f7926f;
      (64'h653f7f19e212e212 & lut_mask_in) : lut = 64'h128d314a271a22c6;
      (64'h7e42e731383f383f & lut_mask_in) : lut = 64'h01f2420bc2fc5d13;
      (64'h0cf4e67cddffddff & lut_mask_in) : lut = 64'hd24ecbb8dcdb79ca;
      (64'hb31d0853a6e6a6e6 & lut_mask_in) : lut = 64'hdb5fec3e277a7600;
      (64'h7372785a55755575 & lut_mask_in) : lut = 64'h8b87f0f5732e7168;

      default  : lut = 0;
    endcase
  end

endmodule

////////////////////////////////////////////////////////////////////////////////
// End Of File
////////////////////////////////////////////////////////////////////////////////
