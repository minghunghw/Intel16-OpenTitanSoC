


# |---------------------|-----------------|
# | Item                | Value           |
# |---------------------|-----------------|
# | Process             | p1222           |
# | Dot Process         | dotp1222_4_opt1 |
# | Library             | 108pp           |
# | Library ID          | b15             |
# | Track Pattern       | tp0             |
# | Redbook DRM Version | 4.0.9           |
# | Ptech Revision      | 31cd5367        |
# | Date                | Jan 31, 2022    |
# | Tech File Version   | 22.05.1-18.44   |
# |---------------------|-----------------|


VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

USEMINSPACING OBS OFF ;

PROPERTYDEFINITIONS
 LAYER techCstId STRING ;
 LAYER sheetResistance REAL ;
 LAYER LEF58_TYPE STRING ;
 LAYER LEF58_ENCLOSURE STRING ;
 LAYER LEF58_ENCLOSURETABLE STRING ;
 LAYER LEF58_CUTCLASS STRING ;
 LAYER LEF58_SPACINGTABLE STRING ;
 LAYER LEF58_WIDTH STRING ;
 LAYER LEF58_MINWIDTH STRING ;
 LAYER LEF58_WIDTHTABLE STRING ;
 LAYER LEF58_EOLKEEPOUT STRING ;
 LAYER LEF58_OPPOSITEEOLSPACING STRING ;
 LAYER LEF58_SPACING STRING ;
 LAYER LEF58_FILLTOFILLSPACING STRING ;
 LAYER LEF58_CORNERSPACING STRING ;
 LAYER LEF58_FORBIDDENSPACING STRING ;
 LAYER LEF58_RECTONLY STRING ;
 LAYER LEF58_AREA STRING ;
 LAYER LEF58_EOLEXTENSIONSPACING STRING ;
 LAYER LEF58_MINSTEP STRING ;
 LAYER LEF58_MAXVIASTACK STRING ;
 LAYER LEF58_FORBIDDENSPACING STRING ;
 LAYER LEF58_KEEPOUTZONE STRING ;
 LAYER LEF58_CUTONCENTERLINE STRING ;
END PROPERTYDEFINITIONS

#################################################
# Overlap layer definitions
#################################################
LAYER OVERLAP
 TYPE OVERLAP ;
END OVERLAP

LAYER OverlapCheck
 TYPE OVERLAP ;
END OverlapCheck

#################################################
# Masterslice layer definitions
#################################################
LAYER diffCheck
 TYPE MASTERSLICE ;
END diffCheck

LAYER deepnwell
 TYPE MASTERSLICE ;
END deepnwell

LAYER nwell
 TYPE MASTERSLICE ;
 PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER ndiff
 TYPE MASTERSLICE ;
END ndiff

LAYER pdiff
 TYPE MASTERSLICE ;
END pdiff

LAYER poly
 TYPE MASTERSLICE ;
END poly

LAYER eoa
 TYPE MASTERSLICE ;
END eoa

LAYER esd_id
 TYPE MASTERSLICE ;
END esd_id

LAYER dummy273
 TYPE MASTERSLICE ;
END dummy273

LAYER dummy81
 TYPE MASTERSLICE ;
END dummy81

LAYER dummy82
 TYPE MASTERSLICE ;
END dummy82

LAYER gcn
 TYPE MASTERSLICE ;
END gcn

LAYER tcn
 TYPE MASTERSLICE ;
END tcn

LAYER emib2bump_zone
 TYPE MASTERSLICE ;
END emib2bump_zone

LAYER emib3bump_zone
 TYPE MASTERSLICE ;
END emib3bump_zone

LAYER TGOXID
 TYPE MASTERSLICE ;
END TGOXID

LAYER emibbump_boundary
 TYPE MASTERSLICE ;
END emibbump_boundary

LAYER GLOBALFILLKOR
 TYPE MASTERSLICE ;
END GLOBALFILLKOR

LAYER v3e7
 TYPE MASTERSLICE ;
END v3e7

LAYER v0_fillBlockage
 TYPE MASTERSLICE ;
END v0_fillBlockage

LAYER m1_fillBlockage
 TYPE MASTERSLICE ;
END m1_fillBlockage

LAYER v1_fillBlockage
 TYPE MASTERSLICE ;
END v1_fillBlockage

LAYER m2_fillBlockage
 TYPE MASTERSLICE ;
END m2_fillBlockage

LAYER v2_fillBlockage
 TYPE MASTERSLICE ;
END v2_fillBlockage

LAYER m3_fillBlockage
 TYPE MASTERSLICE ;
END m3_fillBlockage

LAYER v3_fillBlockage
 TYPE MASTERSLICE ;
END v3_fillBlockage

LAYER m4_fillBlockage
 TYPE MASTERSLICE ;
END m4_fillBlockage

LAYER v4_fillBlockage
 TYPE MASTERSLICE ;
END v4_fillBlockage

LAYER m5_fillBlockage
 TYPE MASTERSLICE ;
END m5_fillBlockage

LAYER v5_fillBlockage
 TYPE MASTERSLICE ;
END v5_fillBlockage

LAYER m6_fillBlockage
 TYPE MASTERSLICE ;
END m6_fillBlockage

LAYER v6_fillBlockage
 TYPE MASTERSLICE ;
END v6_fillBlockage

LAYER m7_fillBlockage
 TYPE MASTERSLICE ;
END m7_fillBlockage

LAYER v7_fillBlockage
 TYPE MASTERSLICE ;
END v7_fillBlockage

LAYER m8_fillBlockage
 TYPE MASTERSLICE ;
END m8_fillBlockage

LAYER v8_fillBlockage
 TYPE MASTERSLICE ;
END v8_fillBlockage

LAYER gmz_fillBlockage
 TYPE MASTERSLICE ;
END gmz_fillBlockage

LAYER vmz_fillBlockage
 TYPE MASTERSLICE ;
END vmz_fillBlockage

LAYER gm0_fillBlockage
 TYPE MASTERSLICE ;
END gm0_fillBlockage

LAYER gv0_fillBlockage
 TYPE MASTERSLICE ;
END gv0_fillBlockage

LAYER gmb_fillBlockage
 TYPE MASTERSLICE ;
END gmb_fillBlockage

LAYER gv1_fillBlockage
 TYPE MASTERSLICE ;
END gv1_fillBlockage

LAYER c4_fillBlockage
 TYPE MASTERSLICE ;
END c4_fillBlockage

LAYER IP
 TYPE MASTERSLICE ;
END IP

#################################################
# Layer definition : v0
#################################################
LAYER v0
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS Via0tcn_64x44 WIDTH 0.0440 LENGTH 0.0640 ;
  CUTCLASS Via0tcn_68x44S WIDTH 0.0440 LENGTH 0.0680 ;
  CUTCLASS Via0gcn_100x44S WIDTH 0.0440 LENGTH 0.1000 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 0.04 ; # V0_23 ;
 # +-----------------------+------------+--------------------------------------------------------------------------------------------+
 # |                                Via spacing table for vias on the same metal segment (SAMEMETAL)                                 |
 # +-----------------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name             | Rule Value | Rule Description                                                                           |
 # +-----------------------+------------+--------------------------------------------------------------------------------------------+
 # | V0_22 - 0.022 - 0.022 | 0.0900     |                                                                                            |
 # | V0_22 - 0.044         | 0.0900     |                                                                                            |
 # | V0_23                 | 0.0400     | Minimum via0 metal aligned edges space in OGD = minimum metal space, when the other edges  |
 # |                       |            | (non-metal limited edges) are perfectly aligned                                            |
 # | V0_24                 | 0.0540     | via0 corner-to-corner space                                                                |
 # | V0_25                 | 0.0840     | via0 edge-to-edge space (V0_23 and V0_26 are exceptions to this rule)                      |
 # | V0_26                 | 0.1520     | Via0_64x44 to Via0_64x44 space in OGD                                                      |
 # +-----------------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0540 
   CUTCLASS                   Via0tcn_64x44 SIDE       Via0tcn_64x44 END       Via0tcn_68x44S SIDE      Via0tcn_68x44S END      Via0gcn_100x44S SIDE     Via0gcn_100x44S END      
   Via0tcn_64x44 SIDE         -       0.0900           -       0.1520          -       0.0900           -       0.1520          -       0.0900           -       0.1520           
   Via0tcn_64x44 END          -       0.1520           -       0.1520          -       0.1520           -       0.0840          -       0.1520           -       0.0840           
   Via0tcn_68x44S SIDE        -       0.0900           -       0.1520          -       0.0900           -       0.1520          -       0.0900           -       0.1520           
   Via0tcn_68x44S END         -       0.1520           -       0.0840          -       0.1520           -       0.0400          -       0.1520           -       0.0400           
   Via0gcn_100x44S SIDE       -       0.0900           -       0.1520          -       0.0900           -       0.1520          -       0.0900           -       0.1520           
   Via0gcn_100x44S END        -       0.1520           -       0.0840          -       0.1520           -       0.0400          -       0.1520           -       0.0400           
  ; " ;
 # +---------------------------------------------------------------------------------------------------------------------+
 # | Forbidden spacing between full facing aligned spacing and standard spacing                                          |
 # +---------------------------------------------------------------------------------------------------------------------+
 # | For each same mask Via spacing at Vx_23 value, a forbidden region must be created to limit spacing from the spacing |
 # | just beyond the Via (Vx_23 + the Via width or height + 0.001) up to the Vx_128 value.                               |
 # +---------------------------------------------------------------------------------------------------------------------+
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                     Forbidden spacing between full facing aligned spacing and standard spacing                      |
 # |                      For each same mask Via spacing at Vx_23 value, a forbidden region must be                      |
 # |                   created to limit spacing from the spacing just beyond the Via (Vx_23 + the Via                    |
 # |                                  width or height + 0.001) up to the Vx_128 value.                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | V0_23     | 0.0400     | Minimum Via0 metal aligned edges space in OGD = minimum metal space, when the other edges  |
 # |           |            | (non-metal limited edges) are perfectly aligned                                            |
 # | V0_25     | 0.0840     | Via0 edge-to-edge space (V0_23 and V0_26 are exceptions to this rule)                      |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_FORBIDDENSPACING "
   FORBIDDENSPACING CUTCLASS Via0gcn_100x44S 0.0410 0.1510  SHORTEDGEONLY    PRL  -0.002 TO Via0tcn_68x44S -0.002 TO Via0gcn_100x44S ;
 " ;
 # -----------------------------------------------------------
 # No clr table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No clr_samenet table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No stack table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 9 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 9 ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 9 ;

END v0








#################################################
# Layer definition : m1
#################################################
LAYER m1
 TYPE ROUTING ;
 DIRECTION VERTICAL ;
 # ------------------------------------------------------------------
 # Width 
 # ------------------------------------------------------------------
 WIDTH    0.0680 ;
 MINWIDTH 0.044 ; # M1_01 ;
 MAXWIDTH 0.1 ; # M1_03 ;
 PROPERTY LEF58_WIDTHTABLE "
  WIDTHTABLE 0.068 0.1 ;
  WIDTHTABLE 0.044 0.1 WRONGDIRECTION ;
 " ;
 # ------------------------------------------------------------------
 # Spacing
 # ------------------------------------------------------------------
 SPACING  0.04 ; # M1_31 ;
 PITCH    0.1080 ; # WIDTH + SPACING 
 # -----------------------------
 # | Width Based Spacing Table |
 # -----------------------------
 # | M1 Width | 68     | 100   |
 # -----------------------------
 # | 68       | 40+    | 50+   |
 # | 100      | 50+    | 50+   |
 # -----------------------------
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE TWOWIDTHS
   WIDTH  0.0000 0.0400 0.0500
   WIDTH  0.0680 0.0500 0.0500
  ; " ; 
 
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                     Metal end-to-end spacing for aligned lines                                      |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | M1_44     | 0.0460     | width_02/03 to width_02/03 end-to-end space PGD (min)                                      |
 # | M1_03     | 0.1000     | width_03 value (PGD/OGD)                                                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.0460 ENDOFLINE  0.1010 WRONGDIRSPACING 0.001  WITHIN 0.0010  ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | M1_80     | 0.0560     | Corner-to-corner space, when corners have no overlap                                       |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.0560 ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                        Metal concave and convex corner rules                                        |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | M1_70     | 0.0170     | Minimum segment length                                                                     |
 # | M1_71     | 0.1080     | Minimum segment lengths, when both adjacent at a concave corner (i.e., length of one of    |
 # |           |            | the edges needs to be greater than M1_71)                                                  |
 # | M1_74     | 0.0700     | Minimum segment lengths, when both adjacent at a convex corner (i.e., length of one of the |
 # |           |            | edges needs to be greater than M1_74)                                                      |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 MINSTEP 0.0170 MAXEDGES 0 ;
 PROPERTY LEF58_MINSTEP "
  MINSTEP 0.1080 MAXEDGES 1 MINADJACENTLENGTH 0.1080 CONCAVECORNER ;
  MINSTEP 0.0700 MAXEDGES 1 MINADJACENTLENGTH 0.0700 CONVEXCORNER ;
 " ;

 # ------------------------------------------------------------------
 # Area and size
 # ------------------------------------------------------------------
 AREA     0.00528000 ; # M1_01 * M1_60 ;
 PROPERTY LEF58_AREA "
  AREA 0.00528 RECTWIDTH 0.044 ;
  AREA 0.00816 RECTWIDTH 0.068 ;
  AREA 0.012 RECTWIDTH 0.1 ;
 " ;
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 5000 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 3000  ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 10000 ;

END m1



#################################################
# Layer definition : v1
#################################################
LAYER v1
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS Via1_60Sx44  WIDTH 0.0440 LENGTH 0.0600 ;
  CUTCLASS Via1_60Sx56  WIDTH 0.0560 LENGTH 0.0600 ;
  CUTCLASS Via1_60Sx76  WIDTH 0.0600 LENGTH 0.0760 ;
  CUTCLASS Via1_60Sx90  WIDTH 0.0600 LENGTH 0.0900 ;
  CUTCLASS Via1_60Sx108 WIDTH 0.0600 LENGTH 0.1080 ;
  CUTCLASS Via1_70x70   WIDTH 0.0700 ;
  CUTCLASS Via1_76x52S  WIDTH 0.0520 LENGTH 0.0760 ;
  CUTCLASS Via1_90x52S  WIDTH 0.0520 LENGTH 0.0900 ;
  CUTCLASS Via1_108x52S WIDTH 0.0520 LENGTH 0.1080 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 0.046 ; # v1_Vm1xa_23 ;
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # |                            Via spacing table for vias on the same metal segment (SAMEMETAL)                            |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name    | Rule Value | Rule Description                                                                           |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | v1_Vm1xa_124 | 0.0880     | v1 min corner-to-corner spacing between via with SA edge in PGD and via with SA edge in    |
 # |              |            | OGD                                                                                        |
 # | v1_Vm1xa_128 | 0.1360     | Unrestricted min v1 edge-to-edge space (SA edges, SA to non-SA edges)                      |
 # | v1_Vm1xa_23  | 0.0460     | Parallel full-facing metal-aligned v1 edges can be as closely spaced as the minimum        |
 # |              |            | allowed m2 space. Min value in PGD.                                                        |
 # | v1_Vm1xa_24  | 0.0660     | Min v1 corner-to-corner space                                                              |
 # | v1_Vm1xa_28  | 0.1560     | Unrestricted min v1 edge-to-edge space (non-SA edges)                                      |
 # | v1_Vm1xa_31  | 0.1100     | Min Via1_70x70-to-Via1_70x70 space                                                         |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0660 
  EXACTALIGNEDSPACING VERTICAL  Via1_70x70 0.11
   CUTCLASS                Via1_60Sx44 SIDE      Via1_60Sx44 END       Via1_60Sx56 SIDE      Via1_60Sx56 END       Via1_60Sx76 SIDE      Via1_60Sx76 END       Via1_60Sx90 SIDE      Via1_60Sx90 END       Via1_60Sx108 SIDE     Via1_60Sx108 END      Via1_70x70            Via1_76x52S SIDE      Via1_76x52S END       Via1_90x52S SIDE      Via1_90x52S END       Via1_108x52S SIDE     Via1_108x52S END      
   Via1_60Sx44 SIDE        -       0.0460        -       0.1560        -       0.0460        -       0.1560        -       0.1560        -       0.0460        -       0.1560        -       0.0460        -       0.1560        -       0.0460        -       0.1360        0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         
   Via1_60Sx44 END         -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         
   Via1_60Sx56 SIDE        -       0.0460        -       0.1560        -       0.0460        -       0.1560        -       0.1560        -       0.0460        -       0.1560        -       0.0460        -       0.1560        -       0.0460        -       0.1360        0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         
   Via1_60Sx56 END         -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         
   Via1_60Sx76 SIDE        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         
   Via1_60Sx76 END         -       0.0460        -       0.1560        -       0.0460        -       0.1560        -       0.1560        -       0.0460        -       0.1560        -       0.0460        -       0.1560        -       0.0460        -       0.1360        0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         
   Via1_60Sx90 SIDE        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         
   Via1_60Sx90 END         -       0.0460        -       0.1560        -       0.0460        -       0.1560        -       0.1560        -       0.0460        -       0.1560        -       0.0460        -       0.1560        -       0.0460        -       0.1360        0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         
   Via1_60Sx108 SIDE       -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         
   Via1_60Sx108 END        -       0.0460        -       0.1560        -       0.0460        -       0.1560        -       0.1560        -       0.0460        -       0.1560        -       0.0460        -       0.1560        -       0.0460        -       0.1360        0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         
   Via1_70x70              -       0.1360        -       0.1560        -       0.1360        -       0.1560        -       0.1560        -       0.1360        -       0.1560        -       0.1360        -       0.1560        -       0.1360        0.1100 0.1100         -       0.1560        -       0.1360        -       0.1560        -       0.1360        -       0.1560        -       0.1360        
   Via1_76x52S SIDE        0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        
   Via1_76x52S END         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         -       0.1360        -       0.1560        -       0.1360        -       0.1560        -       0.1360        -       0.1560        -       0.1360        
   Via1_90x52S SIDE        0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        
   Via1_90x52S END         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         -       0.1360        -       0.1560        -       0.1360        -       0.1560        -       0.1360        -       0.1560        -       0.1360        
   Via1_108x52S SIDE       0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        -       0.1560        
   Via1_108x52S END        0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         0.0880 0.1360         0.0880 0.1560         -       0.1360        -       0.1560        -       0.1360        -       0.1560        -       0.1360        -       0.1560        -       0.1360        
  ; " ;
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # |            Center aligned forbidden spacing limits via spacing from the Mx_25 value up to the Vx_128 value             |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name    | Rule Value | Rule Description                                                                           |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | v1_Vm1xa_23  | 0.0460     | Parallel full-facing metal-aligned v1 edges can be as closely spaced as the minimum        |
 # |              |            | allowed m2 space. Min value in PGD.                                                        |
 # | v1_Vm1xa_128 | 0.1360     | Unrestricted min v1 edge-to-edge space (SA edges, SA to non-SA edges)                      |
 # | m2_Mxa_25    | 0.0600     | width_04/05 OGD to width_04/05 OGD unrestricted space (min)                                |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_FORBIDDENSPACING "
  FORBIDDENSPACING CUTCLASS Via1_60Sx44 0.001 0.0195   PRL  -0.100 TO Via1_60Sx44 -0.100 TO Via1_60Sx56 -0.100 TO Via1_60Sx76 -0.100 TO Via1_60Sx90 -0.100 TO Via1_60Sx108 -0.100 TO Via1_70x70 -0.100 TO Via1_76x52S -0.100 TO Via1_90x52S -0.100 TO Via1_108x52S ;
  FORBIDDENSPACING CUTCLASS Via1_60Sx56 0.001 0.0195   PRL  -0.100 TO Via1_60Sx44 -0.100 TO Via1_60Sx56 -0.100 TO Via1_60Sx76 -0.100 TO Via1_60Sx90 -0.100 TO Via1_60Sx108 -0.100 TO Via1_70x70 -0.100 TO Via1_76x52S -0.100 TO Via1_90x52S -0.100 TO Via1_108x52S ;
  FORBIDDENSPACING CUTCLASS Via1_60Sx76 0.001 0.0195   PRL  -0.100 TO Via1_60Sx44 -0.100 TO Via1_60Sx56 -0.100 TO Via1_60Sx76 -0.100 TO Via1_60Sx90 -0.100 TO Via1_60Sx108 -0.100 TO Via1_70x70 -0.100 TO Via1_76x52S -0.100 TO Via1_90x52S -0.100 TO Via1_108x52S ;
  FORBIDDENSPACING CUTCLASS Via1_60Sx90 0.001 0.0195   PRL  -0.100 TO Via1_60Sx44 -0.100 TO Via1_60Sx56 -0.100 TO Via1_60Sx76 -0.100 TO Via1_60Sx90 -0.100 TO Via1_60Sx108 -0.100 TO Via1_70x70 -0.100 TO Via1_76x52S -0.100 TO Via1_90x52S -0.100 TO Via1_108x52S ;
  FORBIDDENSPACING CUTCLASS Via1_60Sx108 0.001 0.0195   PRL  -0.100 TO Via1_60Sx44 -0.100 TO Via1_60Sx56 -0.100 TO Via1_60Sx76 -0.100 TO Via1_60Sx90 -0.100 TO Via1_60Sx108 -0.100 TO Via1_70x70 -0.100 TO Via1_76x52S -0.100 TO Via1_90x52S -0.100 TO Via1_108x52S ;
  FORBIDDENSPACING CUTCLASS Via1_70x70 0.001 0.0195   PRL  -0.100 TO Via1_60Sx44 -0.100 TO Via1_60Sx44 -0.100 TO Via1_60Sx56 -0.100 TO Via1_60Sx56 -0.100 TO Via1_60Sx76 -0.100 TO Via1_60Sx76 -0.100 TO Via1_60Sx90 -0.100 TO Via1_60Sx90 -0.100 TO Via1_60Sx108 -0.100 TO Via1_60Sx108 -0.100 TO Via1_70x70 -0.100 TO Via1_76x52S -0.100 TO Via1_76x52S -0.100 TO Via1_90x52S -0.100 TO Via1_90x52S -0.100 TO Via1_108x52S -0.100 TO Via1_108x52S ;
  FORBIDDENSPACING CUTCLASS Via1_76x52S 0.001 0.0195   PRL  -0.100 TO Via1_60Sx44 -0.100 TO Via1_60Sx56 -0.100 TO Via1_60Sx76 -0.100 TO Via1_60Sx90 -0.100 TO Via1_60Sx108 -0.100 TO Via1_70x70 -0.100 TO Via1_76x52S -0.100 TO Via1_90x52S -0.100 TO Via1_108x52S ;
  FORBIDDENSPACING CUTCLASS Via1_90x52S 0.001 0.0195   PRL  -0.100 TO Via1_60Sx44 -0.100 TO Via1_60Sx56 -0.100 TO Via1_60Sx76 -0.100 TO Via1_60Sx90 -0.100 TO Via1_60Sx108 -0.100 TO Via1_70x70 -0.100 TO Via1_76x52S -0.100 TO Via1_90x52S -0.100 TO Via1_108x52S ;
  FORBIDDENSPACING CUTCLASS Via1_108x52S 0.001 0.0195   PRL  -0.100 TO Via1_60Sx44 -0.100 TO Via1_60Sx56 -0.100 TO Via1_60Sx76 -0.100 TO Via1_60Sx90 -0.100 TO Via1_60Sx108 -0.100 TO Via1_70x70 -0.100 TO Via1_76x52S -0.100 TO Via1_90x52S -0.100 TO Via1_108x52S ;
 " ;
 # +--------------------------------------------------------------------------+
 # | Via clearance spacing table (Vn to Vn-1)                                 |
 # +--------------------------------------------------------------------------+
 # | This table defines the inter-cut-layer spacing between a className1      |
 # | via in the first row of the table on the layer that this spacing table   |
 # | is being defined to another className2 via in the first column           |
 # | on secondLayerName cut layer.                                            |
 # |                                                                          |
 # | This second layer must be a previously defined                           |
 # | cut layer immediately below the layer that this spacing table is         |
 # | being defined, that is,  one layer look ahead  is not supported.         |
 # |                                                                          |
 # | **NOTE** This cut spacing is ignored for same-net.                       |
 # +--------------------------------------------------------------------------+
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name   | Rule Value | Rule Description                                                                           |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | v1_Vm1xa_32 | 0.0360     | Min v1 to v0 space (on different m1, all-directional check)                                |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0360 LAYER v0
   CUTCLASS                   Via1_60Sx44 SIDE         Via1_60Sx44 END          Via1_60Sx56 SIDE         Via1_60Sx56 END          Via1_60Sx76 SIDE         Via1_60Sx76 END          Via1_60Sx90 SIDE         Via1_60Sx90 END          Via1_60Sx108 SIDE        Via1_60Sx108 END         Via1_70x70               Via1_76x52S SIDE         Via1_76x52S END          Via1_90x52S SIDE         Via1_90x52S END          Via1_108x52S SIDE        Via1_108x52S END         
   Via0tcn_64x44 SIDE         - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0tcn_64x44 END          - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0tcn_68x44S SIDE        - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0tcn_68x44S END         - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0gcn_100x44S SIDE       - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0gcn_100x44S END        - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
  ; " ;
 # +--------------------------------------------------------------------------+
 # | Via clearance spacing table (Vn to Vn-1) for SAMENET                     |
 # +--------------------------------------------------------------------------+
 # | If an inter-cut-layer spacing table is defined for same-net cuts         |
 # | using the SAMENET keyword, the cuts on two different layers can          |
 # | always be stacked if they are exactly aligned (that is, the centers      |
 # | of the cuts are aligned) for same sized cuts. For different sized        |
 # | cuts, it is legal if the smaller cut is completely covered by the        |
 # | bigger cut. Otherwise, the cuts must have cutSpacing                     |
 # | between them.                                                            |
 # +--------------------------------------------------------------------------+
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name   | Rule Value | Rule Description                                                                           |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | v1_Vm1xa_32 | 0.0360     | Min v1 to v0 space (on different m1, all-directional check)                                |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0360 SAMENET LAYER v0
   CUTCLASS                   Via1_60Sx44 SIDE         Via1_60Sx44 END          Via1_60Sx56 SIDE         Via1_60Sx56 END          Via1_60Sx76 SIDE         Via1_60Sx76 END          Via1_60Sx90 SIDE         Via1_60Sx90 END          Via1_60Sx108 SIDE        Via1_60Sx108 END         Via1_70x70               Via1_76x52S SIDE         Via1_76x52S END          Via1_90x52S SIDE         Via1_90x52S END          Via1_108x52S SIDE        Via1_108x52S END         
   Via0tcn_64x44 SIDE         - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0tcn_64x44 END          - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0tcn_68x44S SIDE        - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0tcn_68x44S END         - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0gcn_100x44S SIDE       - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0gcn_100x44S END        - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
  ; " ;
# +-------------------------------------------------------+
# | Via stacking table (Vn to Vn-1 on same metal segment) |
# +-------------------------------------------------------+
# | v1 may stack on v0                               |
# +-------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0000 SAMEMETAL LAYER v0
   CUTCLASS                   Via1_60Sx44 SIDE         Via1_60Sx44 END          Via1_60Sx56 SIDE         Via1_60Sx56 END          Via1_60Sx76 SIDE         Via1_60Sx76 END          Via1_60Sx90 SIDE         Via1_60Sx90 END          Via1_60Sx108 SIDE        Via1_60Sx108 END         Via1_70x70               Via1_76x52S SIDE         Via1_76x52S END          Via1_90x52S SIDE         Via1_90x52S END          Via1_108x52S SIDE        Via1_108x52S END         
   Via0tcn_64x44 SIDE         - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0tcn_64x44 END          - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0tcn_68x44S SIDE        - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0tcn_68x44S END         - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0gcn_100x44S SIDE       - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
   Via0gcn_100x44S END        - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      - -                      
  ; " ;



 # ------------------------------------------------------------------
 # v1_Vm1xa_54 and v1_Vm1xa_154
 # ------------------------------------------------------------------
 PROPERTY LEF58_SPACING "
  SPACING 0.026  LAYER m2 CUTCLASS Via1_60Sx44  CONCAVECORNER ;
  SPACING 0.026  LAYER m2 CUTCLASS Via1_60Sx56  CONCAVECORNER ;
  SPACING 0.026  LAYER m2 CUTCLASS Via1_60Sx76  CONCAVECORNER ;
  SPACING 0.026  LAYER m2 CUTCLASS Via1_60Sx90  CONCAVECORNER ;
  SPACING 0.026  LAYER m2 CUTCLASS Via1_60Sx108 CONCAVECORNER ;
  SPACING 0.019  LAYER m2 CUTCLASS Via1_70x70   CONCAVECORNER ;
  SPACING 0.026  LAYER m2 CUTCLASS Via1_76x52S  CONCAVECORNER ;
  SPACING 0.026  LAYER m2 CUTCLASS Via1_90x52S  CONCAVECORNER ;
  SPACING 0.026  LAYER m2 CUTCLASS Via1_108x52S CONCAVECORNER ;
" ; 




 # ------------------------------------------------------------------
 # v1_Vm1xa_128
 # ------------------------------------------------------------------
 PROPERTY LEF58_KEEPOUTZONE "
  KEEPOUTZONE CUTCLASS Via1_60Sx44  TO Via1_60Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx44  TO Via1_60Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx44  TO Via1_60Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx44  TO Via1_60Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx44  TO Via1_60Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx44  TO Via1_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx44  TO Via1_76x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx44  TO Via1_90x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx44  TO Via1_108x52S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx56  TO Via1_60Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx56  TO Via1_60Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx56  TO Via1_60Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx56  TO Via1_60Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx56  TO Via1_60Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx56  TO Via1_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx56  TO Via1_76x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx56  TO Via1_90x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx56  TO Via1_108x52S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.136 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx76  TO Via1_60Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx76  TO Via1_60Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx76  TO Via1_60Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx76  TO Via1_60Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx76  TO Via1_60Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx76  TO Via1_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx76  TO Via1_76x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx76  TO Via1_90x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx76  TO Via1_108x52S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx90  TO Via1_60Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx90  TO Via1_60Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx90  TO Via1_60Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx90  TO Via1_60Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx90  TO Via1_60Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx90  TO Via1_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx90  TO Via1_76x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx90  TO Via1_90x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx90  TO Via1_108x52S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx108 TO Via1_60Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx108 TO Via1_60Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx108 TO Via1_60Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx108 TO Via1_60Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx108 TO Via1_60Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx108 TO Via1_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx108 TO Via1_76x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx108 TO Via1_90x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_60Sx108 TO Via1_108x52S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_76x52S  TO Via1_60Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_76x52S  TO Via1_60Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_76x52S  TO Via1_60Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_76x52S  TO Via1_60Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_76x52S  TO Via1_60Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_76x52S  TO Via1_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_76x52S  TO Via1_76x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_76x52S  TO Via1_90x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_76x52S  TO Via1_108x52S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_90x52S  TO Via1_60Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_90x52S  TO Via1_60Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_90x52S  TO Via1_60Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_90x52S  TO Via1_60Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_90x52S  TO Via1_60Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_90x52S  TO Via1_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_90x52S  TO Via1_76x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_90x52S  TO Via1_90x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_90x52S  TO Via1_108x52S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_108x52S TO Via1_60Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_108x52S TO Via1_60Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_108x52S TO Via1_60Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_108x52S TO Via1_60Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_108x52S TO Via1_60Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_108x52S TO Via1_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_108x52S TO Via1_76x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_108x52S TO Via1_90x52S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via1_108x52S TO Via1_108x52S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.136 SPIRALEXTENSION 0.0 ;
" ;


 
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 360 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 360 ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 360 ;

END v1








#################################################
# Layer definition : m2
#################################################
LAYER m2
 TYPE ROUTING ;
 DIRECTION HORIZONTAL ;
 # ------------------------------------------------------------------
 # Width 
 # ------------------------------------------------------------------
 WIDTH    0.0440 ;
 MINWIDTH 0.044 ; # m2_Mxa_01 ;
 MAXWIDTH 0.108 ; # m2_Mxa_05 ;
 PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
 PROPERTY LEF58_WIDTHTABLE "
  WIDTHTABLE 0.044 0.056 0.076 0.09 0.108 ;
 " ;
 # ------------------------------------------------------------------
 # Spacing
 # ------------------------------------------------------------------
 SPACING  0.046 ; # m2_Mxa_24 ;
 PITCH    0.0900 ; # WIDTH + SPACING 
 # ----------------------------------
 # |   Width Based Spacing Table    |
 # ----------------------------------
 # | M2 Width | 44/56/76 | 90/108   |
 # ----------------------------------
 # | 44/56/76 | 46+, 46+ | 46+, 46+ |
 # | 90/108   | 46+, 46+ | 60+, 46+ |
 # ----------------------------------
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE TWOWIDTHS
   WIDTH  0.0000 0.0460 0.0460 0.0460 0.0460 0.0460
   WIDTH  0.0440 0.0460 0.0460 0.0460 0.0460 0.0460
   WIDTH  0.0560 0.0460 0.0460 0.0460 0.0460 0.0460
   WIDTH  0.0760 0.0460 0.0460 0.0460 0.0600 0.0600
   WIDTH  0.0900 0.0460 0.0460 0.0460 0.0600 0.0600
  ; " ; 
 
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m2_Mxa_38 | 0.0600     | width_01 OGD to width_04/05 OGD space on one side, when width_01 OGD is sandwiched between |
 # |           |            | width_04/05 OGD on both sides (min)                                                        |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_FORBIDDENSPACING "
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.0890 WITHIN 0.1640 ;
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.1070 WITHIN 0.1640 ;
 " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                     Metal end-to-end spacing for aligned lines                                      |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m2_Mxa_41 | 0.0800     | m2 end-to-end space (min)                                                                  |
 # | m2_Mxa_05 | 0.1080     | width_05 value (OGD/PGD)                                                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.0800 ENDOFLINE  0.1090 WRONGDIRSPACING 0.001  WITHIN 0.0010  ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m2_Mxa_44 | 0.1600     | Width_01 to any width end-to-end space (min) if overlap between facing ends is < m2_Mxa_45 |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.0800 ENDOFLINE 0.0450 WITHIN 0.0010 ENDPRLSPACING 0.1600 PRL 0.0290 ; " ;
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # |                                  Metal end-to-end spacing for misaligned lines                                   |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                        |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # | m2_Mxa_47 | 0.1000     | Min ETE space between a <=m2_Mxa_01 line and a <=m2_Mxa_02 line, when the line ends are |
 # |           |            | not facing each other (The line ends of the <=m2_Mxa_01 wide lines are extended by      |
 # |           |            | m2_Mxa_48 prior to this check)                                                          |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.0570 EXTENSION 0.000 0.0125 0.1000 EXCEPTWITHIN -0.010 -0.001 CLASS M2_C2C ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m2_Mxa_80 | 0.0560     | Min Corner-to-corner space, when corners have no overlap                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.0560 ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                        Metal concave and convex corner rules                                        |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m2_Mxa_70 | 0.0180     | Minimum segment length                                                                     |
 # | m2_Mxa_71 | 0.1000     | Minimum length of at least one segment, when two segments are adjacent at a corner         |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 MINSTEP 0.0180 MAXEDGES 0 ;
 PROPERTY LEF58_MINSTEP "
  MINSTEP 0.1000 MAXEDGES 1 MINADJACENTLENGTH 0.1000 CONCAVECORNER ;
 " ;

 # ------------------------------------------------------------------
 # Area and size
 # ------------------------------------------------------------------
 AREA     0.00704000 ; # m2_Mxa_01 * m2_Mxa_60 ;
 PROPERTY LEF58_AREA "
  AREA 0.00704 RECTWIDTH 0.044 ;
  AREA 0.00896 RECTWIDTH 0.056 ;
  AREA 0.01216 RECTWIDTH 0.076 ;
  AREA 0.0144 RECTWIDTH 0.09 ;
  AREA 0.01728 RECTWIDTH 0.108 ;
 " ;
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 5000 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 3000  ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 10000 ;

END m2



#################################################
# Layer definition : v2
#################################################
LAYER v2
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS Via2_44x58S  WIDTH 0.0440 LENGTH 0.0580 ;
  CUTCLASS Via2_56x58S  WIDTH 0.0560 LENGTH 0.0580 ;
  CUTCLASS Via2_76x58S  WIDTH 0.0580 LENGTH 0.0760 ;
  CUTCLASS Via2_90x58S  WIDTH 0.0580 LENGTH 0.0900 ;
  CUTCLASS Via2_108x58S WIDTH 0.0580 LENGTH 0.1080 ;
  CUTCLASS Via2_70x70   WIDTH 0.0700 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 0.046 ; # v2_Vxa_23 ;
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # |                           Via spacing table for vias on the same metal segment (SAMEMETAL)                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name  | Rule Value | Rule Description                                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | v2_Vxa_128 | 0.1200     | Unrestricted min v2 edge-to-edge space (SA edges, SA to non-SA edges)                      |
 # | v2_Vxa_23  | 0.0460     | Parallel full-facing metal-aligned v2 edges can be as closely spaced as the minimum        |
 # |            |            | allowed m3 space. Min value in OGD.                                                        |
 # | v2_Vxa_24  | 0.0560     | Min v2 corner-to-corner space                                                              |
 # | v2_Vxa_28  | 0.1000     | Unrestricted min v2 edge-to-edge space (non-SA edges)                                      |
 # | v2_Vxa_31  | 0.1100     | Min Via2_70x70-to-Via2_70x70 space                                                         |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0560 
  EXACTALIGNEDSPACING HORIZONTAL  Via2_70x70 0.11
   CUTCLASS                Via2_44x58S SIDE      Via2_44x58S END       Via2_56x58S SIDE      Via2_56x58S END       Via2_76x58S SIDE      Via2_76x58S END       Via2_90x58S SIDE      Via2_90x58S END       Via2_108x58S SIDE     Via2_108x58S END      Via2_70x70            
   Via2_44x58S SIDE        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        
   Via2_44x58S END         -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        
   Via2_56x58S SIDE        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        
   Via2_56x58S END         -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        
   Via2_76x58S SIDE        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        
   Via2_76x58S END         -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        
   Via2_90x58S SIDE        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        
   Via2_90x58S END         -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        
   Via2_108x58S SIDE       -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        
   Via2_108x58S END        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        
   Via2_70x70              -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        0.1100 0.1100         
  ; " ;
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # |           Center aligned forbidden spacing limits via spacing from the Mx_25 value up to the Vx_128 value            |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name  | Rule Value | Rule Description                                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | v2_Vxa_23  | 0.0460     | Parallel full-facing metal-aligned v2 edges can be as closely spaced as the minimum        |
 # |            |            | allowed m3 space. Min value in OGD.                                                        |
 # | v2_Vxa_128 | 0.1200     | Unrestricted min v2 edge-to-edge space (SA edges, SA to non-SA edges)                      |
 # | m3_Mxa_25  | 0.0600     | width_04/05 PGD to width_04/05 PGD unrestricted space (min)                                |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_FORBIDDENSPACING "
  FORBIDDENSPACING CUTCLASS Via2_44x58S 0.001 0.0195   PRL  -0.100 TO Via2_44x58S -0.100 TO Via2_56x58S -0.100 TO Via2_76x58S -0.100 TO Via2_90x58S -0.100 TO Via2_108x58S -0.100 TO Via2_70x70 ;
  FORBIDDENSPACING CUTCLASS Via2_56x58S 0.001 0.0195   PRL  -0.100 TO Via2_44x58S -0.100 TO Via2_56x58S -0.100 TO Via2_76x58S -0.100 TO Via2_90x58S -0.100 TO Via2_108x58S -0.100 TO Via2_70x70 ;
  FORBIDDENSPACING CUTCLASS Via2_76x58S 0.001 0.0195   PRL  -0.100 TO Via2_44x58S -0.100 TO Via2_56x58S -0.100 TO Via2_76x58S -0.100 TO Via2_90x58S -0.100 TO Via2_108x58S -0.100 TO Via2_70x70 ;
  FORBIDDENSPACING CUTCLASS Via2_90x58S 0.001 0.0195   PRL  -0.100 TO Via2_44x58S -0.100 TO Via2_56x58S -0.100 TO Via2_76x58S -0.100 TO Via2_90x58S -0.100 TO Via2_108x58S -0.100 TO Via2_70x70 ;
  FORBIDDENSPACING CUTCLASS Via2_108x58S 0.001 0.0195   PRL  -0.100 TO Via2_44x58S -0.100 TO Via2_56x58S -0.100 TO Via2_76x58S -0.100 TO Via2_90x58S -0.100 TO Via2_108x58S -0.100 TO Via2_70x70 ;
  FORBIDDENSPACING CUTCLASS Via2_70x70 0.001 0.0195   PRL  -0.100 TO Via2_44x58S -0.100 TO Via2_44x58S -0.100 TO Via2_56x58S -0.100 TO Via2_56x58S -0.100 TO Via2_76x58S -0.100 TO Via2_76x58S -0.100 TO Via2_90x58S -0.100 TO Via2_90x58S -0.100 TO Via2_108x58S -0.100 TO Via2_108x58S -0.100 TO Via2_70x70 ;
 " ;
 # +--------------------------------------------------------------------------+
 # | Via clearance spacing table (Vn to Vn-1)                                 |
 # +--------------------------------------------------------------------------+
 # | This table defines the inter-cut-layer spacing between a className1      |
 # | via in the first row of the table on the layer that this spacing table   |
 # | is being defined to another className2 via in the first column           |
 # | on secondLayerName cut layer.                                            |
 # |                                                                          |
 # | This second layer must be a previously defined                           |
 # | cut layer immediately below the layer that this spacing table is         |
 # | being defined, that is,  one layer look ahead  is not supported.         |
 # |                                                                          |
 # | **NOTE** This cut spacing is ignored for same-net.                       |
 # +--------------------------------------------------------------------------+
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | v2_Vxa_32 | 0.0360     | Min v2 to v1 space (on different m2, all-directional check)                                |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0360 LAYER v1
   CUTCLASS                Via2_44x58S SIDE      Via2_44x58S END       Via2_56x58S SIDE      Via2_56x58S END       Via2_76x58S SIDE      Via2_76x58S END       Via2_90x58S SIDE      Via2_90x58S END       Via2_108x58S SIDE     Via2_108x58S END      Via2_70x70            
   Via1_60Sx44 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx44 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx56 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx56 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx76 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx76 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx90 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx90 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx108 SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx108 END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_76x52S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_76x52S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_90x52S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_90x52S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_108x52S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_108x52S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;
 # +--------------------------------------------------------------------------+
 # | Via clearance spacing table (Vn to Vn-1) for SAMENET                     |
 # +--------------------------------------------------------------------------+
 # | If an inter-cut-layer spacing table is defined for same-net cuts         |
 # | using the SAMENET keyword, the cuts on two different layers can          |
 # | always be stacked if they are exactly aligned (that is, the centers      |
 # | of the cuts are aligned) for same sized cuts. For different sized        |
 # | cuts, it is legal if the smaller cut is completely covered by the        |
 # | bigger cut. Otherwise, the cuts must have cutSpacing                     |
 # | between them.                                                            |
 # +--------------------------------------------------------------------------+
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | v2_Vxa_32 | 0.0360     | Min v2 to v1 space (on different m2, all-directional check)                                |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0360 SAMENET LAYER v1
   CUTCLASS                Via2_44x58S SIDE      Via2_44x58S END       Via2_56x58S SIDE      Via2_56x58S END       Via2_76x58S SIDE      Via2_76x58S END       Via2_90x58S SIDE      Via2_90x58S END       Via2_108x58S SIDE     Via2_108x58S END      Via2_70x70            
   Via1_60Sx44 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx44 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx56 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx56 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx76 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx76 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx90 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx90 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx108 SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx108 END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_76x52S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_76x52S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_90x52S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_90x52S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_108x52S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_108x52S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;
# +-------------------------------------------------------+
# | Via stacking table (Vn to Vn-1 on same metal segment) |
# +-------------------------------------------------------+
# | v2 may stack on v1                               |
# +-------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0000 SAMEMETAL LAYER v1
   CUTCLASS                Via2_44x58S SIDE      Via2_44x58S END       Via2_56x58S SIDE      Via2_56x58S END       Via2_76x58S SIDE      Via2_76x58S END       Via2_90x58S SIDE      Via2_90x58S END       Via2_108x58S SIDE     Via2_108x58S END      Via2_70x70            
   Via1_60Sx44 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx44 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx56 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx56 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx76 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx76 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx90 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx90 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx108 SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_60Sx108 END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_76x52S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_76x52S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_90x52S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_90x52S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_108x52S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via1_108x52S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;



 # ------------------------------------------------------------------
 # v2_Vxa_54 and v2_Vxa_154
 # ------------------------------------------------------------------
 PROPERTY LEF58_SPACING "
  SPACING 0.026  LAYER m3 CUTCLASS Via2_44x58S  CONCAVECORNER ;
  SPACING 0.026  LAYER m3 CUTCLASS Via2_56x58S  CONCAVECORNER ;
  SPACING 0.026  LAYER m3 CUTCLASS Via2_76x58S  CONCAVECORNER ;
  SPACING 0.026  LAYER m3 CUTCLASS Via2_90x58S  CONCAVECORNER ;
  SPACING 0.026  LAYER m3 CUTCLASS Via2_108x58S CONCAVECORNER ;
  SPACING 0.019  LAYER m3 CUTCLASS Via2_70x70   CONCAVECORNER ;
" ; 




 # ------------------------------------------------------------------
 # v2_Vxa_128
 # ------------------------------------------------------------------
 PROPERTY LEF58_KEEPOUTZONE "
  KEEPOUTZONE CUTCLASS Via2_44x58S  TO Via2_44x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_44x58S  TO Via2_56x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_44x58S  TO Via2_76x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_44x58S  TO Via2_90x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_44x58S  TO Via2_108x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_44x58S  TO Via2_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_56x58S  TO Via2_44x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_56x58S  TO Via2_56x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_56x58S  TO Via2_76x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_56x58S  TO Via2_90x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_56x58S  TO Via2_108x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_56x58S  TO Via2_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_76x58S  TO Via2_44x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_76x58S  TO Via2_56x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_76x58S  TO Via2_76x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_76x58S  TO Via2_90x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_76x58S  TO Via2_108x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_76x58S  TO Via2_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_90x58S  TO Via2_44x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_90x58S  TO Via2_56x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_90x58S  TO Via2_76x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_90x58S  TO Via2_90x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_90x58S  TO Via2_108x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_90x58S  TO Via2_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_108x58S TO Via2_44x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_108x58S TO Via2_56x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_108x58S TO Via2_76x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_108x58S TO Via2_90x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_108x58S TO Via2_108x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via2_108x58S TO Via2_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
" ;


 
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 360 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 360 ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 360 ;

END v2








#################################################
# Layer definition : m3
#################################################
LAYER m3
 TYPE ROUTING ;
 DIRECTION VERTICAL ;
 # ------------------------------------------------------------------
 # Width 
 # ------------------------------------------------------------------
 WIDTH    0.0440 ;
 MINWIDTH 0.044 ; # m3_Mxa_01 ;
 MAXWIDTH 0.108 ; # m3_Mxa_05 ;
 PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
 PROPERTY LEF58_WIDTHTABLE "
  WIDTHTABLE 0.044 0.056 0.076 0.09 0.108 ;
 " ;
 # ------------------------------------------------------------------
 # Spacing
 # ------------------------------------------------------------------
 SPACING  0.046 ; # m3_Mxa_24 ;
 PITCH    0.0900 ; # WIDTH + SPACING 
 # ----------------------------------
 # |   Width Based Spacing Table    |
 # ----------------------------------
 # | M3 Width | 44/56/76 | 90/108   |
 # ----------------------------------
 # | 44/56/76 | 46+, 46+ | 46+, 46+ |
 # | 90/108   | 46+, 46+ | 60+, 46+ |
 # ----------------------------------
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE TWOWIDTHS
   WIDTH  0.0000 0.0460 0.0460 0.0460 0.0460 0.0460
   WIDTH  0.0440 0.0460 0.0460 0.0460 0.0460 0.0460
   WIDTH  0.0560 0.0460 0.0460 0.0460 0.0460 0.0460
   WIDTH  0.0760 0.0460 0.0460 0.0460 0.0600 0.0600
   WIDTH  0.0900 0.0460 0.0460 0.0460 0.0600 0.0600
  ; " ; 
 
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m3_Mxa_38 | 0.0600     | width_01 PGD to width_04/05 PGD space on one side, when width_01 PGD is sandwiched between |
 # |           |            | width_04/05 PGD on both sides (min)                                                        |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_FORBIDDENSPACING "
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.0890 WITHIN 0.1640 ;
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.1070 WITHIN 0.1640 ;
 " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                     Metal end-to-end spacing for aligned lines                                      |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m3_Mxa_41 | 0.0800     | m3 end-to-end space (min)                                                                  |
 # | m3_Mxa_05 | 0.1080     | width_05 value (PGD/OGD)                                                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.0800 ENDOFLINE  0.1090 WRONGDIRSPACING 0.001  WITHIN 0.0010  ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m3_Mxa_44 | 0.1600     | Width_01 to any width end-to-end space (min) if overlap between facing ends is < m3_Mxa_45 |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.0800 ENDOFLINE 0.0450 WITHIN 0.0010 ENDPRLSPACING 0.1600 PRL 0.0290 ; " ;
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # |                                  Metal end-to-end spacing for misaligned lines                                   |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                        |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # | m3_Mxa_47 | 0.1000     | Min ETE space between a <=m3_Mxa_01 line and a <=m3_Mxa_02 line, when the line ends are |
 # |           |            | not facing each other (The line ends of the <=m3_Mxa_01 wide lines are extended by      |
 # |           |            | m3_Mxa_48 prior to this check)                                                          |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.0570 EXTENSION 0.000 0.0125 0.1000 EXCEPTWITHIN -0.010 -0.001 CLASS M3_C2C ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m3_Mxa_80 | 0.0560     | Min Corner-to-corner space, when corners have no overlap                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.0560 ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                        Metal concave and convex corner rules                                        |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m3_Mxa_70 | 0.0180     | Minimum segment length                                                                     |
 # | m3_Mxa_71 | 0.1000     | Minimum length of at least one segment, when two segments are adjacent at a corner         |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 MINSTEP 0.0180 MAXEDGES 0 ;
 PROPERTY LEF58_MINSTEP "
  MINSTEP 0.1000 MAXEDGES 1 MINADJACENTLENGTH 0.1000 CONCAVECORNER ;
 " ;

 # ------------------------------------------------------------------
 # Area and size
 # ------------------------------------------------------------------
 AREA     0.00704000 ; # m3_Mxa_01 * m3_Mxa_60 ;
 PROPERTY LEF58_AREA "
  AREA 0.00704 RECTWIDTH 0.044 ;
  AREA 0.00896 RECTWIDTH 0.056 ;
  AREA 0.01216 RECTWIDTH 0.076 ;
  AREA 0.0144 RECTWIDTH 0.09 ;
  AREA 0.01728 RECTWIDTH 0.108 ;
 " ;
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 5000 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 3000  ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 10000 ;

END m3



#################################################
# Layer definition : v3
#################################################
LAYER v3
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS Via3_58Sx44  WIDTH 0.0440 LENGTH 0.0580 ;
  CUTCLASS Via3_58Sx56  WIDTH 0.0560 LENGTH 0.0580 ;
  CUTCLASS Via3_58Sx76  WIDTH 0.0580 LENGTH 0.0760 ;
  CUTCLASS Via3_58Sx90  WIDTH 0.0580 LENGTH 0.0900 ;
  CUTCLASS Via3_58Sx108 WIDTH 0.0580 LENGTH 0.1080 ;
  CUTCLASS Via3_70x70   WIDTH 0.0700 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 0.046 ; # v3_Vxa_23 ;
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # |                           Via spacing table for vias on the same metal segment (SAMEMETAL)                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name  | Rule Value | Rule Description                                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | v3_Vxa_128 | 0.1200     | Unrestricted min v3 edge-to-edge space (SA edges, SA to non-SA edges)                      |
 # | v3_Vxa_23  | 0.0460     | Parallel full-facing metal-aligned v3 edges can be as closely spaced as the minimum        |
 # |            |            | allowed m4 space. Min value in PGD.                                                        |
 # | v3_Vxa_24  | 0.0560     | Min v3 corner-to-corner space                                                              |
 # | v3_Vxa_28  | 0.1000     | Unrestricted min v3 edge-to-edge space (non-SA edges)                                      |
 # | v3_Vxa_31  | 0.1100     | Min Via3_70x70-to-Via3_70x70 space                                                         |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0560 
  EXACTALIGNEDSPACING VERTICAL  Via3_70x70 0.11
   CUTCLASS                Via3_58Sx44 SIDE      Via3_58Sx44 END       Via3_58Sx56 SIDE      Via3_58Sx56 END       Via3_58Sx76 SIDE      Via3_58Sx76 END       Via3_58Sx90 SIDE      Via3_58Sx90 END       Via3_58Sx108 SIDE     Via3_58Sx108 END      Via3_70x70            
   Via3_58Sx44 SIDE        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        
   Via3_58Sx44 END         -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        
   Via3_58Sx56 SIDE        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        
   Via3_58Sx56 END         -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        
   Via3_58Sx76 SIDE        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        
   Via3_58Sx76 END         -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        
   Via3_58Sx90 SIDE        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        
   Via3_58Sx90 END         -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        
   Via3_58Sx108 SIDE       -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        
   Via3_58Sx108 END        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        
   Via3_70x70              -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        0.1100 0.1100         
  ; " ;
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # |           Center aligned forbidden spacing limits via spacing from the Mx_25 value up to the Vx_128 value            |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name  | Rule Value | Rule Description                                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | v3_Vxa_23  | 0.0460     | Parallel full-facing metal-aligned v3 edges can be as closely spaced as the minimum        |
 # |            |            | allowed m4 space. Min value in PGD.                                                        |
 # | v3_Vxa_128 | 0.1200     | Unrestricted min v3 edge-to-edge space (SA edges, SA to non-SA edges)                      |
 # | m4_Mxa_25  | 0.0600     | width_04/05 OGD to width_04/05 OGD unrestricted space (min)                                |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_FORBIDDENSPACING "
  FORBIDDENSPACING CUTCLASS Via3_58Sx44 0.001 0.0195   PRL  -0.100 TO Via3_58Sx44 -0.100 TO Via3_58Sx56 -0.100 TO Via3_58Sx76 -0.100 TO Via3_58Sx90 -0.100 TO Via3_58Sx108 -0.100 TO Via3_70x70 ;
  FORBIDDENSPACING CUTCLASS Via3_58Sx56 0.001 0.0195   PRL  -0.100 TO Via3_58Sx44 -0.100 TO Via3_58Sx56 -0.100 TO Via3_58Sx76 -0.100 TO Via3_58Sx90 -0.100 TO Via3_58Sx108 -0.100 TO Via3_70x70 ;
  FORBIDDENSPACING CUTCLASS Via3_58Sx76 0.001 0.0195   PRL  -0.100 TO Via3_58Sx44 -0.100 TO Via3_58Sx56 -0.100 TO Via3_58Sx76 -0.100 TO Via3_58Sx90 -0.100 TO Via3_58Sx108 -0.100 TO Via3_70x70 ;
  FORBIDDENSPACING CUTCLASS Via3_58Sx90 0.001 0.0195   PRL  -0.100 TO Via3_58Sx44 -0.100 TO Via3_58Sx56 -0.100 TO Via3_58Sx76 -0.100 TO Via3_58Sx90 -0.100 TO Via3_58Sx108 -0.100 TO Via3_70x70 ;
  FORBIDDENSPACING CUTCLASS Via3_58Sx108 0.001 0.0195   PRL  -0.100 TO Via3_58Sx44 -0.100 TO Via3_58Sx56 -0.100 TO Via3_58Sx76 -0.100 TO Via3_58Sx90 -0.100 TO Via3_58Sx108 -0.100 TO Via3_70x70 ;
  FORBIDDENSPACING CUTCLASS Via3_70x70 0.001 0.0195   PRL  -0.100 TO Via3_58Sx44 -0.100 TO Via3_58Sx44 -0.100 TO Via3_58Sx56 -0.100 TO Via3_58Sx56 -0.100 TO Via3_58Sx76 -0.100 TO Via3_58Sx76 -0.100 TO Via3_58Sx90 -0.100 TO Via3_58Sx90 -0.100 TO Via3_58Sx108 -0.100 TO Via3_58Sx108 -0.100 TO Via3_70x70 ;
 " ;
 # +--------------------------------------------------------------------------+
 # | Via clearance spacing table (Vn to Vn-1)                                 |
 # +--------------------------------------------------------------------------+
 # | This table defines the inter-cut-layer spacing between a className1      |
 # | via in the first row of the table on the layer that this spacing table   |
 # | is being defined to another className2 via in the first column           |
 # | on secondLayerName cut layer.                                            |
 # |                                                                          |
 # | This second layer must be a previously defined                           |
 # | cut layer immediately below the layer that this spacing table is         |
 # | being defined, that is,  one layer look ahead  is not supported.         |
 # |                                                                          |
 # | **NOTE** This cut spacing is ignored for same-net.                       |
 # +--------------------------------------------------------------------------+
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | v3_Vxa_32 | 0.0360     | Min v3 to v2 space (on different m3, all-directional check)                                |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0360 LAYER v2
   CUTCLASS                Via3_58Sx44 SIDE      Via3_58Sx44 END       Via3_58Sx56 SIDE      Via3_58Sx56 END       Via3_58Sx76 SIDE      Via3_58Sx76 END       Via3_58Sx90 SIDE      Via3_58Sx90 END       Via3_58Sx108 SIDE     Via3_58Sx108 END      Via3_70x70            
   Via2_44x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_44x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_56x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_56x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_76x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_76x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_90x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_90x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_108x58S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_108x58S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;
 # +--------------------------------------------------------------------------+
 # | Via clearance spacing table (Vn to Vn-1) for SAMENET                     |
 # +--------------------------------------------------------------------------+
 # | If an inter-cut-layer spacing table is defined for same-net cuts         |
 # | using the SAMENET keyword, the cuts on two different layers can          |
 # | always be stacked if they are exactly aligned (that is, the centers      |
 # | of the cuts are aligned) for same sized cuts. For different sized        |
 # | cuts, it is legal if the smaller cut is completely covered by the        |
 # | bigger cut. Otherwise, the cuts must have cutSpacing                     |
 # | between them.                                                            |
 # +--------------------------------------------------------------------------+
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | v3_Vxa_32 | 0.0360     | Min v3 to v2 space (on different m3, all-directional check)                                |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0360 SAMENET LAYER v2
   CUTCLASS                Via3_58Sx44 SIDE      Via3_58Sx44 END       Via3_58Sx56 SIDE      Via3_58Sx56 END       Via3_58Sx76 SIDE      Via3_58Sx76 END       Via3_58Sx90 SIDE      Via3_58Sx90 END       Via3_58Sx108 SIDE     Via3_58Sx108 END      Via3_70x70            
   Via2_44x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_44x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_56x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_56x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_76x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_76x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_90x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_90x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_108x58S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_108x58S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;
# +-------------------------------------------------------+
# | Via stacking table (Vn to Vn-1 on same metal segment) |
# +-------------------------------------------------------+
# | v3 may stack on v2                               |
# +-------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0000 SAMEMETAL LAYER v2
   CUTCLASS                Via3_58Sx44 SIDE      Via3_58Sx44 END       Via3_58Sx56 SIDE      Via3_58Sx56 END       Via3_58Sx76 SIDE      Via3_58Sx76 END       Via3_58Sx90 SIDE      Via3_58Sx90 END       Via3_58Sx108 SIDE     Via3_58Sx108 END      Via3_70x70            
   Via2_44x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_44x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_56x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_56x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_76x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_76x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_90x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_90x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_108x58S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_108x58S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via2_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;



 # ------------------------------------------------------------------
 # v3_Vxa_54 and v3_Vxa_154
 # ------------------------------------------------------------------
 PROPERTY LEF58_SPACING "
  SPACING 0.026  LAYER m4 CUTCLASS Via3_58Sx44  CONCAVECORNER ;
  SPACING 0.026  LAYER m4 CUTCLASS Via3_58Sx56  CONCAVECORNER ;
  SPACING 0.026  LAYER m4 CUTCLASS Via3_58Sx76  CONCAVECORNER ;
  SPACING 0.026  LAYER m4 CUTCLASS Via3_58Sx90  CONCAVECORNER ;
  SPACING 0.026  LAYER m4 CUTCLASS Via3_58Sx108 CONCAVECORNER ;
  SPACING 0.019  LAYER m4 CUTCLASS Via3_70x70   CONCAVECORNER ;
" ; 




 # ------------------------------------------------------------------
 # v3_Vxa_128
 # ------------------------------------------------------------------
 PROPERTY LEF58_KEEPOUTZONE "
  KEEPOUTZONE CUTCLASS Via3_58Sx44  TO Via3_58Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx44  TO Via3_58Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx44  TO Via3_58Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx44  TO Via3_58Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx44  TO Via3_58Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx44  TO Via3_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx56  TO Via3_58Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx56  TO Via3_58Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx56  TO Via3_58Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx56  TO Via3_58Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx56  TO Via3_58Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx56  TO Via3_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx76  TO Via3_58Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx76  TO Via3_58Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx76  TO Via3_58Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx76  TO Via3_58Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx76  TO Via3_58Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx76  TO Via3_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx90  TO Via3_58Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx90  TO Via3_58Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx90  TO Via3_58Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx90  TO Via3_58Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx90  TO Via3_58Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx90  TO Via3_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx108 TO Via3_58Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx108 TO Via3_58Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx108 TO Via3_58Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx108 TO Via3_58Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx108 TO Via3_58Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via3_58Sx108 TO Via3_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
" ;


 
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 360 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 360 ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 360 ;

END v3








#################################################
# Layer definition : m4
#################################################
LAYER m4
 TYPE ROUTING ;
 DIRECTION HORIZONTAL ;
 # ------------------------------------------------------------------
 # Width 
 # ------------------------------------------------------------------
 WIDTH    0.0440 ;
 MINWIDTH 0.044 ; # m4_Mxa_01 ;
 MAXWIDTH 0.108 ; # m4_Mxa_05 ;
 PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
 PROPERTY LEF58_WIDTHTABLE "
  WIDTHTABLE 0.044 0.056 0.076 0.09 0.108 ;
 " ;
 # ------------------------------------------------------------------
 # Spacing
 # ------------------------------------------------------------------
 SPACING  0.046 ; # m4_Mxa_24 ;
 PITCH    0.0900 ; # WIDTH + SPACING 
 # ----------------------------------
 # |   Width Based Spacing Table    |
 # ----------------------------------
 # | M4 Width | 44/56/76 | 90/108   |
 # ----------------------------------
 # | 44/56/76 | 46+, 46+ | 46+, 46+ |
 # | 90/108   | 46+, 46+ | 60+, 46+ |
 # ----------------------------------
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE TWOWIDTHS
   WIDTH  0.0000 0.0460 0.0460 0.0460 0.0460 0.0460
   WIDTH  0.0440 0.0460 0.0460 0.0460 0.0460 0.0460
   WIDTH  0.0560 0.0460 0.0460 0.0460 0.0460 0.0460
   WIDTH  0.0760 0.0460 0.0460 0.0460 0.0600 0.0600
   WIDTH  0.0900 0.0460 0.0460 0.0460 0.0600 0.0600
  ; " ; 
 
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m4_Mxa_38 | 0.0600     | width_01 OGD to width_04/05 OGD space on one side, when width_01 OGD is sandwiched between |
 # |           |            | width_04/05 OGD on both sides (min)                                                        |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_FORBIDDENSPACING "
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.0890 WITHIN 0.1640 ;
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.1070 WITHIN 0.1640 ;
 " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                     Metal end-to-end spacing for aligned lines                                      |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m4_Mxa_41 | 0.0800     | m4 end-to-end space (min)                                                                  |
 # | m4_Mxa_05 | 0.1080     | width_05 value (OGD/PGD)                                                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.1090 EXTENSION 0.000 0.010 0.0800 CLASS M4_E2E ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m4_Mxa_44 | 0.1600     | Width_01 to any width end-to-end space (min) if overlap between facing ends is < m4_Mxa_45 |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.0800 ENDOFLINE 0.0450 WITHIN 0.0010 ENDPRLSPACING 0.1600 PRL 0.0290 ; " ;
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # |                                  Metal end-to-end spacing for misaligned lines                                   |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                        |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # | m4_Mxa_47 | 0.1000     | Min ETE space between a <=m4_Mxa_01 line and a <=m4_Mxa_02 line, when the line ends are |
 # |           |            | not facing each other (The line ends of the <=m4_Mxa_01 wide lines are extended by      |
 # |           |            | m4_Mxa_48 prior to this check)                                                          |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.0570 EXTENSION 0.000 0.0125 0.1000 EXCEPTWITHIN -0.010 -0.001 CLASS M4_C2C ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m4_Mxa_80 | 0.0560     | Min Corner-to-corner space, when corners have no overlap                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.0560 ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                        Metal concave and convex corner rules                                        |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m4_Mxa_70 | 0.0180     | Minimum segment length                                                                     |
 # | m4_Mxa_71 | 0.1000     | Minimum length of at least one segment, when two segments are adjacent at a corner         |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 MINSTEP 0.0180 MAXEDGES 0 ;
 PROPERTY LEF58_MINSTEP "
  MINSTEP 0.1000 MAXEDGES 1 MINADJACENTLENGTH 0.1000 CONCAVECORNER ;
 " ;

 # ------------------------------------------------------------------
 # Area and size
 # ------------------------------------------------------------------
 AREA     0.00704000 ; # m4_Mxa_01 * m4_Mxa_60 ;
 PROPERTY LEF58_AREA "
  AREA 0.00704 RECTWIDTH 0.044 ;
  AREA 0.00896 RECTWIDTH 0.056 ;
  AREA 0.01216 RECTWIDTH 0.076 ;
  AREA 0.0144 RECTWIDTH 0.09 ;
  AREA 0.01728 RECTWIDTH 0.108 ;
 " ;
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 5000 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 3000  ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 10000 ;

END m4



#################################################
# Layer definition : v4
#################################################
LAYER v4
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS Via4_44x58S  WIDTH 0.0440 LENGTH 0.0580 ;
  CUTCLASS Via4_56x58S  WIDTH 0.0560 LENGTH 0.0580 ;
  CUTCLASS Via4_76x58S  WIDTH 0.0580 LENGTH 0.0760 ;
  CUTCLASS Via4_90x58S  WIDTH 0.0580 LENGTH 0.0900 ;
  CUTCLASS Via4_108x58S WIDTH 0.0580 LENGTH 0.1080 ;
  CUTCLASS Via4_160x58S WIDTH 0.0580 LENGTH 0.1600 ;
  CUTCLASS Via4_70x70   WIDTH 0.0700 ;
  CUTCLASS Via4_90x90   WIDTH 0.0900 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 0.046 ; # v4_Vxaxb_23 ;
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # |                            Via spacing table for vias on the same metal segment (SAMEMETAL)                            |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name    | Rule Value | Rule Description                                                                           |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | v4_Vxaxb_128 | 0.1200     | Unrestricted min v4 edge-to-edge space (SA edges, SA to non-SA edges)                      |
 # | v4_Vxaxb_23  | 0.0460     | Parallel full-facing metal-aligned v4 edges can be as closely spaced as the minimum        |
 # |              |            | allowed m5 space. Min value in OGD.                                                        |
 # | v4_Vxaxb_24  | 0.0560     | Min v4 corner-to-corner space                                                              |
 # | v4_Vxaxb_28  | 0.1000     | Unrestricted min v4 edge-to-edge space (non-SA edges)                                      |
 # | v4_Vxaxb_31  | 0.1100     | Min Via4_70x70-to-Via4_70x70 space                                                         |
 # | v4_Vxaxb_34  | 0.1300     | Min Via4_90x90 to any other v4 space                                                       |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0560 
  EXACTALIGNEDSPACING HORIZONTAL  Via4_70x70 0.11 Via4_90x90 0.13
   CUTCLASS                Via4_44x58S SIDE      Via4_44x58S END       Via4_56x58S SIDE      Via4_56x58S END       Via4_76x58S SIDE      Via4_76x58S END       Via4_90x58S SIDE      Via4_90x58S END       Via4_108x58S SIDE     Via4_108x58S END      Via4_160x58S SIDE     Via4_160x58S END      Via4_70x70            Via4_90x90            
   Via4_44x58S SIDE        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via4_44x58S END         -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via4_56x58S SIDE        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via4_56x58S END         -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via4_76x58S SIDE        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via4_76x58S END         -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via4_90x58S SIDE        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via4_90x58S END         -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via4_108x58S SIDE       -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via4_108x58S END        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via4_160x58S SIDE       -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via4_160x58S END        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via4_70x70              -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        0.1100 0.1100         0.1300 0.1300         
   Via4_90x90              0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         
  ; " ;
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # |            Center aligned forbidden spacing limits via spacing from the Mx_25 value up to the Vx_128 value             |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name    | Rule Value | Rule Description                                                                           |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | v4_Vxaxb_23  | 0.0460     | Parallel full-facing metal-aligned v4 edges can be as closely spaced as the minimum        |
 # |              |            | allowed m5 space. Min value in OGD.                                                        |
 # | v4_Vxaxb_128 | 0.1200     | Unrestricted min v4 edge-to-edge space (SA edges, SA to non-SA edges)                      |
 # | m5_Mxb_25    | 0.0600     | width_04/05 PGD to width_04/05 PGD unrestricted space (min)                                |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_FORBIDDENSPACING "
  FORBIDDENSPACING CUTCLASS Via4_44x58S 0.001 0.0195   PRL  -0.100 TO Via4_44x58S -0.100 TO Via4_56x58S -0.100 TO Via4_76x58S -0.100 TO Via4_90x58S -0.100 TO Via4_108x58S -0.100 TO Via4_160x58S -0.100 TO Via4_70x70 -0.100 TO Via4_90x90 ;
  FORBIDDENSPACING CUTCLASS Via4_56x58S 0.001 0.0195   PRL  -0.100 TO Via4_44x58S -0.100 TO Via4_56x58S -0.100 TO Via4_76x58S -0.100 TO Via4_90x58S -0.100 TO Via4_108x58S -0.100 TO Via4_160x58S -0.100 TO Via4_70x70 -0.100 TO Via4_90x90 ;
  FORBIDDENSPACING CUTCLASS Via4_76x58S 0.001 0.0195   PRL  -0.100 TO Via4_44x58S -0.100 TO Via4_56x58S -0.100 TO Via4_76x58S -0.100 TO Via4_90x58S -0.100 TO Via4_108x58S -0.100 TO Via4_160x58S -0.100 TO Via4_70x70 -0.100 TO Via4_90x90 ;
  FORBIDDENSPACING CUTCLASS Via4_90x58S 0.001 0.0195   PRL  -0.100 TO Via4_44x58S -0.100 TO Via4_56x58S -0.100 TO Via4_76x58S -0.100 TO Via4_90x58S -0.100 TO Via4_108x58S -0.100 TO Via4_160x58S -0.100 TO Via4_70x70 -0.100 TO Via4_90x90 ;
  FORBIDDENSPACING CUTCLASS Via4_108x58S 0.001 0.0195   PRL  -0.100 TO Via4_44x58S -0.100 TO Via4_56x58S -0.100 TO Via4_76x58S -0.100 TO Via4_90x58S -0.100 TO Via4_108x58S -0.100 TO Via4_160x58S -0.100 TO Via4_70x70 -0.100 TO Via4_90x90 ;
  FORBIDDENSPACING CUTCLASS Via4_160x58S 0.001 0.0195   PRL  -0.100 TO Via4_44x58S -0.100 TO Via4_56x58S -0.100 TO Via4_76x58S -0.100 TO Via4_90x58S -0.100 TO Via4_108x58S -0.100 TO Via4_160x58S -0.100 TO Via4_70x70 -0.100 TO Via4_90x90 ;
  FORBIDDENSPACING CUTCLASS Via4_70x70 0.001 0.0195   PRL  -0.100 TO Via4_44x58S -0.100 TO Via4_44x58S -0.100 TO Via4_56x58S -0.100 TO Via4_56x58S -0.100 TO Via4_76x58S -0.100 TO Via4_76x58S -0.100 TO Via4_90x58S -0.100 TO Via4_90x58S -0.100 TO Via4_108x58S -0.100 TO Via4_108x58S -0.100 TO Via4_160x58S -0.100 TO Via4_160x58S -0.100 TO Via4_70x70 -0.100 TO Via4_90x90 ;
  FORBIDDENSPACING CUTCLASS Via4_90x90 0.001 0.0195   PRL  -0.100 TO Via4_44x58S -0.100 TO Via4_44x58S -0.100 TO Via4_56x58S -0.100 TO Via4_56x58S -0.100 TO Via4_76x58S -0.100 TO Via4_76x58S -0.100 TO Via4_90x58S -0.100 TO Via4_90x58S -0.100 TO Via4_108x58S -0.100 TO Via4_108x58S -0.100 TO Via4_160x58S -0.100 TO Via4_160x58S -0.100 TO Via4_70x70 -0.100 TO Via4_90x90 ;
 " ;
 # +--------------------------------------------------------------------------+
 # | Via clearance spacing table (Vn to Vn-1)                                 |
 # +--------------------------------------------------------------------------+
 # | This table defines the inter-cut-layer spacing between a className1      |
 # | via in the first row of the table on the layer that this spacing table   |
 # | is being defined to another className2 via in the first column           |
 # | on secondLayerName cut layer.                                            |
 # |                                                                          |
 # | This second layer must be a previously defined                           |
 # | cut layer immediately below the layer that this spacing table is         |
 # | being defined, that is,  one layer look ahead  is not supported.         |
 # |                                                                          |
 # | **NOTE** This cut spacing is ignored for same-net.                       |
 # +--------------------------------------------------------------------------+
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name   | Rule Value | Rule Description                                                                           |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | v4_Vxaxb_32 | 0.0360     | Min v4 to v3 space (on different m4, all-directional check)                                |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0360 LAYER v3
   CUTCLASS                Via4_44x58S SIDE      Via4_44x58S END       Via4_56x58S SIDE      Via4_56x58S END       Via4_76x58S SIDE      Via4_76x58S END       Via4_90x58S SIDE      Via4_90x58S END       Via4_108x58S SIDE     Via4_108x58S END      Via4_160x58S SIDE     Via4_160x58S END      Via4_70x70            Via4_90x90            
   Via3_58Sx44 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx44 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx56 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx56 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx76 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx76 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx90 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx90 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx108 SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx108 END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;
 # +--------------------------------------------------------------------------+
 # | Via clearance spacing table (Vn to Vn-1) for SAMENET                     |
 # +--------------------------------------------------------------------------+
 # | If an inter-cut-layer spacing table is defined for same-net cuts         |
 # | using the SAMENET keyword, the cuts on two different layers can          |
 # | always be stacked if they are exactly aligned (that is, the centers      |
 # | of the cuts are aligned) for same sized cuts. For different sized        |
 # | cuts, it is legal if the smaller cut is completely covered by the        |
 # | bigger cut. Otherwise, the cuts must have cutSpacing                     |
 # | between them.                                                            |
 # +--------------------------------------------------------------------------+
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name   | Rule Value | Rule Description                                                                           |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | v4_Vxaxb_32 | 0.0360     | Min v4 to v3 space (on different m4, all-directional check)                                |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0360 SAMENET LAYER v3
   CUTCLASS                Via4_44x58S SIDE      Via4_44x58S END       Via4_56x58S SIDE      Via4_56x58S END       Via4_76x58S SIDE      Via4_76x58S END       Via4_90x58S SIDE      Via4_90x58S END       Via4_108x58S SIDE     Via4_108x58S END      Via4_160x58S SIDE     Via4_160x58S END      Via4_70x70            Via4_90x90            
   Via3_58Sx44 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx44 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx56 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx56 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx76 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx76 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx90 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx90 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx108 SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx108 END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;
# +-------------------------------------------------------+
# | Via stacking table (Vn to Vn-1 on same metal segment) |
# +-------------------------------------------------------+
# | v4 may stack on v3                               |
# +-------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0000 SAMEMETAL LAYER v3
   CUTCLASS                Via4_44x58S SIDE      Via4_44x58S END       Via4_56x58S SIDE      Via4_56x58S END       Via4_76x58S SIDE      Via4_76x58S END       Via4_90x58S SIDE      Via4_90x58S END       Via4_108x58S SIDE     Via4_108x58S END      Via4_160x58S SIDE     Via4_160x58S END      Via4_70x70            Via4_90x90            
   Via3_58Sx44 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx44 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx56 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx56 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx76 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx76 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx90 SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx90 END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx108 SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_58Sx108 END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via3_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;



 # ------------------------------------------------------------------
 # v4_Vxaxb_54 and v4_Vxaxb_154
 # ------------------------------------------------------------------
 PROPERTY LEF58_SPACING "
  SPACING 0.026  LAYER m5 CUTCLASS Via4_44x58S  CONCAVECORNER ;
  SPACING 0.026  LAYER m5 CUTCLASS Via4_56x58S  CONCAVECORNER ;
  SPACING 0.026  LAYER m5 CUTCLASS Via4_76x58S  CONCAVECORNER ;
  SPACING 0.026  LAYER m5 CUTCLASS Via4_90x58S  CONCAVECORNER ;
  SPACING 0.026  LAYER m5 CUTCLASS Via4_108x58S CONCAVECORNER ;
  SPACING 0.026  LAYER m5 CUTCLASS Via4_160x58S CONCAVECORNER ;
  SPACING 0.019  LAYER m5 CUTCLASS Via4_70x70   CONCAVECORNER ;
  SPACING 0.026  LAYER m5 CUTCLASS Via4_90x90   CONCAVECORNER ;
" ; 




 # ------------------------------------------------------------------
 # v4_Vxaxb_128
 # ------------------------------------------------------------------
 PROPERTY LEF58_KEEPOUTZONE "
  KEEPOUTZONE CUTCLASS Via4_44x58S  TO Via4_44x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_44x58S  TO Via4_56x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_44x58S  TO Via4_76x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_44x58S  TO Via4_90x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_44x58S  TO Via4_108x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_44x58S  TO Via4_160x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_44x58S  TO Via4_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_44x58S  TO Via4_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_56x58S  TO Via4_44x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_56x58S  TO Via4_56x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_56x58S  TO Via4_76x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_56x58S  TO Via4_90x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_56x58S  TO Via4_108x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_56x58S  TO Via4_160x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_56x58S  TO Via4_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_56x58S  TO Via4_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_76x58S  TO Via4_44x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_76x58S  TO Via4_56x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_76x58S  TO Via4_76x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_76x58S  TO Via4_90x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_76x58S  TO Via4_108x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_76x58S  TO Via4_160x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_76x58S  TO Via4_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_76x58S  TO Via4_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_90x58S  TO Via4_44x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_90x58S  TO Via4_56x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_90x58S  TO Via4_76x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_90x58S  TO Via4_90x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_90x58S  TO Via4_108x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_90x58S  TO Via4_160x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_90x58S  TO Via4_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_90x58S  TO Via4_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_108x58S TO Via4_44x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_108x58S TO Via4_56x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_108x58S TO Via4_76x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_108x58S TO Via4_90x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_108x58S TO Via4_108x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_108x58S TO Via4_160x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_108x58S TO Via4_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_108x58S TO Via4_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_160x58S TO Via4_44x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_160x58S TO Via4_56x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_160x58S TO Via4_76x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_160x58S TO Via4_90x58S  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_160x58S TO Via4_108x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_160x58S TO Via4_160x58S EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_160x58S TO Via4_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via4_160x58S TO Via4_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
" ;


 
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 420 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 420 ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 420 ;

END v4








#################################################
# Layer definition : m5
#################################################
LAYER m5
 TYPE ROUTING ;
 DIRECTION VERTICAL ;
 # ------------------------------------------------------------------
 # Width 
 # ------------------------------------------------------------------
 WIDTH    0.0440 ;
 MINWIDTH 0.044 ; # m5_Mxb_01 ;
 MAXWIDTH 0.2 ; # m5_Mxb_07 ;
 PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
 PROPERTY LEF58_WIDTHTABLE "
  WIDTHTABLE 0.044 0.056 0.076 0.09 0.108 0.16 0.2 ;
 " ;
 # ------------------------------------------------------------------
 # Spacing
 # ------------------------------------------------------------------
 SPACING  0.046 ; # m5_Mxb_24 ;
 PITCH    0.0900 ; # WIDTH + SPACING 
 # -----------------------------------------------------------------------------
 # |                         Width Based Spacing Table                         |
 # -----------------------------------------------------------------------------
 # | M5 Width | 44            | 56/76    | 90/108   | 160      | 200           |
 # -----------------------------------------------------------------------------
 # | 44       | 46+, 46+      | 46+, 46+ | 46+, 46+ | 60+, 46+ | 60+, 58+, 46+ |
 # | 56/76    | 46+, 46+      | 46+, 46+ | 46+, 46+ | 60+, 46+ | 60+, 46+      |
 # | 90/108   | 46+, 46+      | 46+, 46+ | 60+, 46+ | 60+, 46+ | 60+, 46+      |
 # | 160      | 60+, 46+      | 60+, 46+ | 60+, 46+ | 60+, 46+ | 60+, 46+      |
 # | 200      | 60+, 58+, 46+ | 60+, 46+ | 60+, 46+ | 60+, 46+ | 60+, 46+      |
 # -----------------------------------------------------------------------------
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE TWOWIDTHS
   WIDTH  0.0000 0.0460 0.0460 0.0460 0.0460 0.0460 0.0600 0.0580
   WIDTH  0.0440 0.0460 0.0460 0.0460 0.0460 0.0460 0.0600 0.0600
   WIDTH  0.0560 0.0460 0.0460 0.0460 0.0460 0.0460 0.0600 0.0600
   WIDTH  0.0760 0.0460 0.0460 0.0460 0.0600 0.0600 0.0600 0.0600
   WIDTH  0.0900 0.0460 0.0460 0.0460 0.0600 0.0600 0.0600 0.0600
   WIDTH  0.1080 0.0600 0.0600 0.0600 0.0600 0.0600 0.0600 0.0600
   WIDTH  0.1600 0.0580 0.0600 0.0600 0.0600 0.0600 0.0600 0.0600
  ; " ; 
 
 # +-----------+------------+------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                         |
 # +-----------+------------+------------------------------------------------------------------------------------------+
 # | m5_Mxb_38 | 0.0600     | width_01 PGD to width >= width_04 PGD space on one side, when width_01 PGD is sandwiched |
 # |           |            | between width >= width_04 PGD on both sides (min)                                        |
 # +-----------+------------+------------------------------------------------------------------------------------------+
 PROPERTY LEF58_FORBIDDENSPACING "
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.0890 WITHIN 0.1640 ;
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.1070 WITHIN 0.1640 ;
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.1590 WITHIN 0.1640 ;
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.1990 WITHIN 0.1640 ;
 " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                     Metal end-to-end spacing for aligned lines                                      |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m5_Mxb_41 | 0.0800     | m5 end-to-end space (min)                                                                  |
 # | m5_Mxb_07 | 0.2000     | width_07 value (OGD/PGD)                                                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.0800 ENDOFLINE  0.2010 WRONGDIRSPACING 0.001  WITHIN 0.0010  ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m5_Mxb_44 | 0.1600     | Width_01 to any width end-to-end space (min) if overlap between facing ends is < m5_Mxb_45 |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.0800 ENDOFLINE 0.0450 WITHIN 0.0010 ENDPRLSPACING 0.1600 PRL 0.0290 ; " ;
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # |                                  Metal end-to-end spacing for misaligned lines                                   |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                        |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # | m5_Mxb_47 | 0.1000     | Min ETE space between a <=m5_Mxb_01 line and a <=m5_Mxb_02 line, when the line ends are |
 # |           |            | not facing each other (The line ends of the <=m5_Mxb_01 wide lines are extended by      |
 # |           |            | m5_Mxb_48 prior to this check)                                                          |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.0570 EXTENSION 0.000 0.0125 0.1000 EXCEPTWITHIN -0.010 -0.001 CLASS M5_C2C ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m5_Mxb_80 | 0.0560     | Min Corner-to-corner space, when corners have no overlap                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.0560 ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                        Metal concave and convex corner rules                                        |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m5_Mxb_70 | 0.0180     | Minimum segment length                                                                     |
 # | m5_Mxb_71 | 0.1000     | Minimum length of at least one segment, when two segments are adjacent at a corner         |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 MINSTEP 0.0180 MAXEDGES 0 ;
 PROPERTY LEF58_MINSTEP "
  MINSTEP 0.1000 MAXEDGES 1 MINADJACENTLENGTH 0.1000 CONCAVECORNER ;
 " ;

 # ------------------------------------------------------------------
 # Area and size
 # ------------------------------------------------------------------
 AREA     0.00704000 ; # m5_Mxb_01 * m5_Mxb_60 ;
 PROPERTY LEF58_AREA "
  AREA 0.00704 RECTWIDTH 0.044 ;
  AREA 0.00896 RECTWIDTH 0.056 ;
  AREA 0.01216 RECTWIDTH 0.076 ;
  AREA 0.0144 RECTWIDTH 0.09 ;
  AREA 0.01728 RECTWIDTH 0.108 ;
  AREA 0.0256 RECTWIDTH 0.16 ;
  AREA 0.04 RECTWIDTH 0.2 ;
 " ;
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 5000 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 3000  ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 10000 ;

END m5



#################################################
# Layer definition : v5
#################################################
LAYER v5
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS Via5_58Sx44  WIDTH 0.0440 LENGTH 0.0580 ;
  CUTCLASS Via5_58Sx56  WIDTH 0.0560 LENGTH 0.0580 ;
  CUTCLASS Via5_58Sx76  WIDTH 0.0580 LENGTH 0.0760 ;
  CUTCLASS Via5_58Sx90  WIDTH 0.0580 LENGTH 0.0900 ;
  CUTCLASS Via5_58Sx108 WIDTH 0.0580 LENGTH 0.1080 ;
  CUTCLASS Via5_58Sx160 WIDTH 0.0580 LENGTH 0.1600 ;
  CUTCLASS Via5_70x70   WIDTH 0.0700 ;
  CUTCLASS Via5_90x90   WIDTH 0.0900 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 0.046 ; # v5_Vxbxc_23 ;
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # |                            Via spacing table for vias on the same metal segment (SAMEMETAL)                            |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name    | Rule Value | Rule Description                                                                           |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | v5_Vxbxc_128 | 0.1200     | Unrestricted min v5 edge-to-edge space (SA edges, SA to non-SA edges)                      |
 # | v5_Vxbxc_23  | 0.0460     | Parallel full-facing metal-aligned v5 edges can be as closely spaced as the minimum        |
 # |              |            | allowed m6 space. Min value in PGD.                                                        |
 # | v5_Vxbxc_24  | 0.0560     | Min v5 corner-to-corner space                                                              |
 # | v5_Vxbxc_28  | 0.1000     | Unrestricted min v5 edge-to-edge space (non-SA edges)                                      |
 # | v5_Vxbxc_31  | 0.1100     | Min Via5_70x70-to-Via5_70x70 space                                                         |
 # | v5_Vxbxc_34  | 0.1300     | Min Via5_90x90 to any other v5 space                                                       |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0560 
  EXACTALIGNEDSPACING VERTICAL  Via5_70x70 0.11 Via5_90x90 0.13
   CUTCLASS                Via5_58Sx44 SIDE      Via5_58Sx44 END       Via5_58Sx56 SIDE      Via5_58Sx56 END       Via5_58Sx76 SIDE      Via5_58Sx76 END       Via5_58Sx90 SIDE      Via5_58Sx90 END       Via5_58Sx108 SIDE     Via5_58Sx108 END      Via5_58Sx160 SIDE     Via5_58Sx160 END      Via5_70x70            Via5_90x90            
   Via5_58Sx44 SIDE        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via5_58Sx44 END         -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via5_58Sx56 SIDE        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via5_58Sx56 END         -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via5_58Sx76 SIDE        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via5_58Sx76 END         -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via5_58Sx90 SIDE        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via5_58Sx90 END         -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via5_58Sx108 SIDE       -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via5_58Sx108 END        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via5_58Sx160 SIDE       -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        0.1300 0.1300         
   Via5_58Sx160 END        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        -       0.0460        -       0.1200        0.1300 0.1300         
   Via5_70x70              -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        -       0.1000        -       0.1200        0.1100 0.1100         0.1300 0.1300         
   Via5_90x90              0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         0.1300 0.1300         
  ; " ;
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # |            Center aligned forbidden spacing limits via spacing from the Mx_25 value up to the Vx_128 value             |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name    | Rule Value | Rule Description                                                                           |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | v5_Vxbxc_23  | 0.0460     | Parallel full-facing metal-aligned v5 edges can be as closely spaced as the minimum        |
 # |              |            | allowed m6 space. Min value in PGD.                                                        |
 # | v5_Vxbxc_128 | 0.1200     | Unrestricted min v5 edge-to-edge space (SA edges, SA to non-SA edges)                      |
 # | m6_Mxc_27    | 0.1000     | width_08 OGD to any width OGD unrestricted space (min)                                     |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_FORBIDDENSPACING "
  FORBIDDENSPACING CUTCLASS Via5_58Sx44 0.001 0.0195   PRL  -0.100 TO Via5_58Sx44 -0.100 TO Via5_58Sx56 -0.100 TO Via5_58Sx76 -0.100 TO Via5_58Sx90 -0.100 TO Via5_58Sx108 -0.100 TO Via5_58Sx160 -0.100 TO Via5_70x70 -0.100 TO Via5_90x90 ;
  FORBIDDENSPACING CUTCLASS Via5_58Sx56 0.001 0.0195   PRL  -0.100 TO Via5_58Sx44 -0.100 TO Via5_58Sx56 -0.100 TO Via5_58Sx76 -0.100 TO Via5_58Sx90 -0.100 TO Via5_58Sx108 -0.100 TO Via5_58Sx160 -0.100 TO Via5_70x70 -0.100 TO Via5_90x90 ;
  FORBIDDENSPACING CUTCLASS Via5_58Sx76 0.001 0.0195   PRL  -0.100 TO Via5_58Sx44 -0.100 TO Via5_58Sx56 -0.100 TO Via5_58Sx76 -0.100 TO Via5_58Sx90 -0.100 TO Via5_58Sx108 -0.100 TO Via5_58Sx160 -0.100 TO Via5_70x70 -0.100 TO Via5_90x90 ;
  FORBIDDENSPACING CUTCLASS Via5_58Sx90 0.001 0.0195   PRL  -0.100 TO Via5_58Sx44 -0.100 TO Via5_58Sx56 -0.100 TO Via5_58Sx76 -0.100 TO Via5_58Sx90 -0.100 TO Via5_58Sx108 -0.100 TO Via5_58Sx160 -0.100 TO Via5_70x70 -0.100 TO Via5_90x90 ;
  FORBIDDENSPACING CUTCLASS Via5_58Sx108 0.001 0.0195   PRL  -0.100 TO Via5_58Sx44 -0.100 TO Via5_58Sx56 -0.100 TO Via5_58Sx76 -0.100 TO Via5_58Sx90 -0.100 TO Via5_58Sx108 -0.100 TO Via5_58Sx160 -0.100 TO Via5_70x70 -0.100 TO Via5_90x90 ;
  FORBIDDENSPACING CUTCLASS Via5_58Sx160 0.001 0.0195   PRL  -0.100 TO Via5_58Sx44 -0.100 TO Via5_58Sx56 -0.100 TO Via5_58Sx76 -0.100 TO Via5_58Sx90 -0.100 TO Via5_58Sx108 -0.100 TO Via5_58Sx160 -0.100 TO Via5_70x70 -0.100 TO Via5_90x90 ;
  FORBIDDENSPACING CUTCLASS Via5_70x70 0.001 0.0195   PRL  -0.100 TO Via5_58Sx44 -0.100 TO Via5_58Sx44 -0.100 TO Via5_58Sx56 -0.100 TO Via5_58Sx56 -0.100 TO Via5_58Sx76 -0.100 TO Via5_58Sx76 -0.100 TO Via5_58Sx90 -0.100 TO Via5_58Sx90 -0.100 TO Via5_58Sx108 -0.100 TO Via5_58Sx108 -0.100 TO Via5_58Sx160 -0.100 TO Via5_58Sx160 -0.100 TO Via5_70x70 -0.100 TO Via5_90x90 ;
  FORBIDDENSPACING CUTCLASS Via5_90x90 0.001 0.0195   PRL  -0.100 TO Via5_58Sx44 -0.100 TO Via5_58Sx44 -0.100 TO Via5_58Sx56 -0.100 TO Via5_58Sx56 -0.100 TO Via5_58Sx76 -0.100 TO Via5_58Sx76 -0.100 TO Via5_58Sx90 -0.100 TO Via5_58Sx90 -0.100 TO Via5_58Sx108 -0.100 TO Via5_58Sx108 -0.100 TO Via5_58Sx160 -0.100 TO Via5_58Sx160 -0.100 TO Via5_70x70 -0.100 TO Via5_90x90 ;
 " ;
 # +--------------------------------------------------------------------------+
 # | Via clearance spacing table (Vn to Vn-1)                                 |
 # +--------------------------------------------------------------------------+
 # | This table defines the inter-cut-layer spacing between a className1      |
 # | via in the first row of the table on the layer that this spacing table   |
 # | is being defined to another className2 via in the first column           |
 # | on secondLayerName cut layer.                                            |
 # |                                                                          |
 # | This second layer must be a previously defined                           |
 # | cut layer immediately below the layer that this spacing table is         |
 # | being defined, that is,  one layer look ahead  is not supported.         |
 # |                                                                          |
 # | **NOTE** This cut spacing is ignored for same-net.                       |
 # +--------------------------------------------------------------------------+
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name   | Rule Value | Rule Description                                                                           |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | v5_Vxbxc_32 | 0.0360     | Min v5 to v4 space (on different m5, all-directional check)                                |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0360 LAYER v4
   CUTCLASS                Via5_58Sx44 SIDE      Via5_58Sx44 END       Via5_58Sx56 SIDE      Via5_58Sx56 END       Via5_58Sx76 SIDE      Via5_58Sx76 END       Via5_58Sx90 SIDE      Via5_58Sx90 END       Via5_58Sx108 SIDE     Via5_58Sx108 END      Via5_58Sx160 SIDE     Via5_58Sx160 END      Via5_70x70            Via5_90x90            
   Via4_44x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_44x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_56x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_56x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_76x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_76x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_90x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_90x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_108x58S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_108x58S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_160x58S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_160x58S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_90x90              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;
 # +--------------------------------------------------------------------------+
 # | Via clearance spacing table (Vn to Vn-1) for SAMENET                     |
 # +--------------------------------------------------------------------------+
 # | If an inter-cut-layer spacing table is defined for same-net cuts         |
 # | using the SAMENET keyword, the cuts on two different layers can          |
 # | always be stacked if they are exactly aligned (that is, the centers      |
 # | of the cuts are aligned) for same sized cuts. For different sized        |
 # | cuts, it is legal if the smaller cut is completely covered by the        |
 # | bigger cut. Otherwise, the cuts must have cutSpacing                     |
 # | between them.                                                            |
 # +--------------------------------------------------------------------------+
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name   | Rule Value | Rule Description                                                                           |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | v5_Vxbxc_32 | 0.0360     | Min v5 to v4 space (on different m5, all-directional check)                                |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0360 SAMENET LAYER v4
   CUTCLASS                Via5_58Sx44 SIDE      Via5_58Sx44 END       Via5_58Sx56 SIDE      Via5_58Sx56 END       Via5_58Sx76 SIDE      Via5_58Sx76 END       Via5_58Sx90 SIDE      Via5_58Sx90 END       Via5_58Sx108 SIDE     Via5_58Sx108 END      Via5_58Sx160 SIDE     Via5_58Sx160 END      Via5_70x70            Via5_90x90            
   Via4_44x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_44x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_56x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_56x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_76x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_76x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_90x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_90x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_108x58S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_108x58S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_160x58S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_160x58S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_90x90              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;
# +-------------------------------------------------------+
# | Via stacking table (Vn to Vn-1 on same metal segment) |
# +-------------------------------------------------------+
# | v5 may stack on v4                               |
# +-------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.0000 SAMEMETAL LAYER v4
   CUTCLASS                Via5_58Sx44 SIDE      Via5_58Sx44 END       Via5_58Sx56 SIDE      Via5_58Sx56 END       Via5_58Sx76 SIDE      Via5_58Sx76 END       Via5_58Sx90 SIDE      Via5_58Sx90 END       Via5_58Sx108 SIDE     Via5_58Sx108 END      Via5_58Sx160 SIDE     Via5_58Sx160 END      Via5_70x70            Via5_90x90            
   Via4_44x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_44x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_56x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_56x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_76x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_76x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_90x58S SIDE        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_90x58S END         - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_108x58S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_108x58S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_160x58S SIDE       - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_160x58S END        - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_70x70              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
   Via4_90x90              - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   - -                   
  ; " ;



 # ------------------------------------------------------------------
 # v5_Vxbxc_54 and v5_Vxbxc_154
 # ------------------------------------------------------------------
 PROPERTY LEF58_SPACING "
  SPACING 0.026  LAYER m6 CUTCLASS Via5_58Sx44  CONCAVECORNER ;
  SPACING 0.026  LAYER m6 CUTCLASS Via5_58Sx56  CONCAVECORNER ;
  SPACING 0.026  LAYER m6 CUTCLASS Via5_58Sx76  CONCAVECORNER ;
  SPACING 0.026  LAYER m6 CUTCLASS Via5_58Sx90  CONCAVECORNER ;
  SPACING 0.026  LAYER m6 CUTCLASS Via5_58Sx108 CONCAVECORNER ;
  SPACING 0.026  LAYER m6 CUTCLASS Via5_58Sx160 CONCAVECORNER ;
  SPACING 0.019  LAYER m6 CUTCLASS Via5_70x70   CONCAVECORNER ;
  SPACING 0.026  LAYER m6 CUTCLASS Via5_90x90   CONCAVECORNER ;
" ; 




 # ------------------------------------------------------------------
 # v5_Vxbxc_128
 # ------------------------------------------------------------------
 PROPERTY LEF58_KEEPOUTZONE "
  KEEPOUTZONE CUTCLASS Via5_58Sx44  TO Via5_58Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx44  TO Via5_58Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx44  TO Via5_58Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx44  TO Via5_58Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx44  TO Via5_58Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx44  TO Via5_58Sx160 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx44  TO Via5_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx44  TO Via5_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx56  TO Via5_58Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx56  TO Via5_58Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx56  TO Via5_58Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx56  TO Via5_58Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx56  TO Via5_58Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx56  TO Via5_58Sx160 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx56  TO Via5_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx56  TO Via5_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.12 SIDEEXTENSION 0.0 0.0 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx76  TO Via5_58Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx76  TO Via5_58Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx76  TO Via5_58Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx76  TO Via5_58Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx76  TO Via5_58Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx76  TO Via5_58Sx160 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx76  TO Via5_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx76  TO Via5_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx90  TO Via5_58Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx90  TO Via5_58Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx90  TO Via5_58Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx90  TO Via5_58Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx90  TO Via5_58Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx90  TO Via5_58Sx160 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx90  TO Via5_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx90  TO Via5_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx108 TO Via5_58Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx108 TO Via5_58Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx108 TO Via5_58Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx108 TO Via5_58Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx108 TO Via5_58Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx108 TO Via5_58Sx160 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx108 TO Via5_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx108 TO Via5_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx160 TO Via5_58Sx44  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx160 TO Via5_58Sx56  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx160 TO Via5_58Sx76  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx160 TO Via5_58Sx90  EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx160 TO Via5_58Sx108 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx160 TO Via5_58Sx160 EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx160 TO Via5_70x70   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
  KEEPOUTZONE CUTCLASS Via5_58Sx160 TO Via5_90x90   EXCEPTEXACTALIGNED 0.046 ENDEXTENSION 0.0 0.0 SIDEEXTENSION 0.0 0.12 SPIRALEXTENSION 0.0 ;
" ;


 
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 420 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 420 ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 420 ;

END v5








#################################################
# Layer definition : m6
#################################################
LAYER m6
 TYPE ROUTING ;
 DIRECTION HORIZONTAL ;
 # ------------------------------------------------------------------
 # Width 
 # ------------------------------------------------------------------
 WIDTH    0.0440 ;
 MINWIDTH 0.044 ; # m6_Mxc_01 ;
 MAXWIDTH 0.4 ; # m6_Mxc_08 ;
 PROPERTY LEF58_WIDTHTABLE "
  WIDTHTABLE 0.044 0.056 0.076 0.09 0.108 0.16 0.2 0.4 ;
 " ;
 # ------------------------------------------------------------------
 # Spacing
 # ------------------------------------------------------------------
 SPACING  0.046 ; # m6_Mxc_24 ;
 PITCH    0.0900 ; # WIDTH + SPACING 
 # ------------------------------------------------------------
 # |                Width Based Spacing Table                 |
 # ------------------------------------------------------------
 # | M6 Width | 44/56/76  | 90/108    | 160/200   | 400       |
 # ------------------------------------------------------------
 # | 44/56/76 | 46+, 46+  | 46+, 46+  | 60+, 46+  | 100+, 46+ |
 # | 90/108   | 46+, 46+  | 60+, 46+  | 60+, 46+  | 100+, 46+ |
 # | 160/200  | 60+, 46+  | 60+, 46+  | 60+, 46+  | 100+, 46+ |
 # | 400      | 100+, 46+ | 100+, 46+ | 100+, 46+ | 100+, 46+ |
 # ------------------------------------------------------------
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE TWOWIDTHS
   WIDTH  0.0000 0.0460 0.0460 0.0460 0.0460 0.0460 0.0600 0.0600 0.1000
   WIDTH  0.0440 0.0460 0.0460 0.0460 0.0460 0.0460 0.0600 0.0600 0.1000
   WIDTH  0.0560 0.0460 0.0460 0.0460 0.0460 0.0460 0.0600 0.0600 0.1000
   WIDTH  0.0760 0.0460 0.0460 0.0460 0.0600 0.0600 0.0600 0.0600 0.1000
   WIDTH  0.0900 0.0460 0.0460 0.0460 0.0600 0.0600 0.0600 0.0600 0.1000
   WIDTH  0.1080 0.0600 0.0600 0.0600 0.0600 0.0600 0.0600 0.0600 0.1000
   WIDTH  0.1600 0.0600 0.0600 0.0600 0.0600 0.0600 0.0600 0.0600 0.1000
   WIDTH  0.2000 0.1000 0.1000 0.1000 0.1000 0.1000 0.1000 0.1000 0.1000
  ; " ; 
 
 # +-----------+------------+------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                         |
 # +-----------+------------+------------------------------------------------------------------------------------------+
 # | m6_Mxc_38 | 0.0600     | width_01 OGD to width >= width_04 OGD space on one side, when width_01 OGD is sandwiched |
 # |           |            | between width >= width_04 OGD on both sides (min)                                        |
 # +-----------+------------+------------------------------------------------------------------------------------------+
 PROPERTY LEF58_FORBIDDENSPACING "
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.0890 WITHIN 0.1640 ;
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.1070 WITHIN 0.1640 ;
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.1590 WITHIN 0.1640 ;
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.1990 WITHIN 0.1640 ;
  FORBIDDENSPACING 0.000 0.0590 WIDTHRANGE 0.000 0.0450 PRL 0.0  OTHERWIDTH 0.3990 WITHIN 0.1640 ;
 " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                     Metal end-to-end spacing for aligned lines                                      |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m6_Mxc_41 | 0.0800     | m6 end-to-end space (min)                                                                  |
 # | m6_Mxc_08 | 0.4000     | width_08 value (OGD/PGD)                                                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.0800 ENDOFLINE  0.4010 WRONGDIRSPACING 0.001  WITHIN 0.0010  ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m6_Mxc_44 | 0.1600     | Width_01 to any width end-to-end space (min) if overlap between facing ends is < m6_Mxc_45 |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.0800 ENDOFLINE 0.0450 WITHIN 0.0010 ENDPRLSPACING 0.1600 PRL 0.0290 ; " ;
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # |                                  Metal end-to-end spacing for misaligned lines                                   |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                        |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 # | m6_Mxc_47 | 0.1000     | Min ETE space between a <=m6_Mxc_01 line and a <=m6_Mxc_02 line, when the line ends are |
 # |           |            | not facing each other (The line ends of the <=m6_Mxc_01 wide lines are extended by      |
 # |           |            | m6_Mxc_48 prior to this check)                                                          |
 # +-----------+------------+-----------------------------------------------------------------------------------------+
 PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.0570 EXTENSION 0.000 0.0125 0.1000 EXCEPTWITHIN -0.010 -0.001 CLASS M6_C2C ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m6_Mxc_80 | 0.0560     | Min Corner-to-corner space, when corners have no overlap                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.0560 ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                        Metal concave and convex corner rules                                        |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m6_Mxc_70 | 0.0180     | Minimum segment length                                                                     |
 # | m6_Mxc_71 | 0.1000     | Minimum length of at least one segment, when two segments are adjacent at a corner         |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 MINSTEP 0.0180 MAXEDGES 0 ;
 PROPERTY LEF58_MINSTEP "
  MINSTEP 0.1000 MAXEDGES 1 MINADJACENTLENGTH 0.1400 CONCAVECORNER ;
 " ;

 # ------------------------------------------------------------------
 # Area and size
 # ------------------------------------------------------------------
 AREA     0.00704000 ; # m6_Mxc_01 * m6_Mxc_60 ;
 PROPERTY LEF58_AREA "
  AREA 0.00704 RECTWIDTH 0.044 ;
  AREA 0.00896 RECTWIDTH 0.056 ;
  AREA 0.01216 RECTWIDTH 0.076 ;
  AREA 0.0144 RECTWIDTH 0.09 ;
  AREA 0.01728 RECTWIDTH 0.108 ;
  AREA 0.0256 RECTWIDTH 0.16 ;
  AREA 0.04 RECTWIDTH 0.2 ;
  AREA 0.16 RECTWIDTH 0.4 ;
 " ;
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 5000 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 3000  ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 10000 ;

END m6



#################################################
# Layer definition : v6
#################################################
LAYER v6
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS Via6_200x120 WIDTH 0.1200 LENGTH 0.2000 ;
  CUTCLASS Via6_400x120 WIDTH 0.1200 LENGTH 0.4000 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_ENCLOSURETABLE "
  ENCLOSURETABLE CUTCLASS Via6_200x120 
  WIDTH 0.181 ABOVE  0.0300 0.0300 0.0600 0.0600 INCLUDEABUTTED  ;
 " ;

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 0.24 ; # v6_Vxcyb_33 ;
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # |                           Via spacing table for vias on the same metal segment (SAMEMETAL)                            |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name   | Rule Value | Rule Description                                                                           |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | v6_Vxcyb_33 | 0.2400     | v6-to-v6 spacing (edges), minimum, all-directional check                                   |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.2400 
   CUTCLASS                 Via6_200x120 SIDE      Via6_200x120 END         Via6_400x120 SIDE      Via6_400x120 END       
   Via6_200x120 SIDE        -       -              -       -                -       -              -       -              
   Via6_200x120 END         -       -              -       -                -       -              -       -              
   Via6_400x120 SIDE        -       -              -       -                -       -              -       -              
   Via6_400x120 END         -       -              -       -                -       -              -       -              
  ; " ;
 # -----------------------------------------------------------
 # No clr table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No clr_samenet table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No stack table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 550 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 550 ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 550 ;

END v6








#################################################
# Layer definition : m7
#################################################
LAYER m7
 TYPE ROUTING ;
 DIRECTION VERTICAL ;
 # ------------------------------------------------------------------
 # Width 
 # ------------------------------------------------------------------
 WIDTH    0.1800 ;
 MINWIDTH 0.18 ; # m7_Myb_01 ;
 MAXWIDTH 0.9 ; # m7_Myb_21 ;
 PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
 # ------------------------------------------------------------------
 # Spacing
 # ------------------------------------------------------------------
 SPACING  0.18 ; # m7_Myb_02 ;
 PITCH    0.3600 ; # WIDTH + SPACING 
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                     Metal end-to-end spacing for aligned lines                                      |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m7_Myb_03 | 0.2400     | Min m7 space (end-to-end, attacker). Applies to segments identified as line ends.          |
 # | m7_Myb_21 | 0.9000     | m7 width allowed range, maximum                                                            |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.2400 ENDOFLINE  0.9010 WRONGDIRSPACING 0.001  WITHIN 0.0010  ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                        Metal concave and convex corner rules                                        |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m7_Myb_27 | 0.3080     | Minimum length of at least one segment, when two segments are adjacent at a corner         |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_MINSTEP "
  MINSTEP 0.3080 MAXEDGES 1 MINADJACENTLENGTH 0.3080 CONCAVECORNER ;
  MINSTEP 0.3080 MAXEDGES 1 MINBETWEENLENGTH 0.3080 ;
 " ;

 # ------------------------------------------------------------------
 # Area and size
 # ------------------------------------------------------------------
 AREA     0.09000000 ; # m7_Myb_24 ;
 PROPERTY LEF58_AREA "
  AREA 0.09 RECTWIDTH 0.18 ;
  AREA 0.1074 RECTWIDTH 0.24 ;
  AREA 0.1195 RECTWIDTH 0.27 ;
  AREA 0.1317 RECTWIDTH 0.23 ;
  AREA 0.1438 RECTWIDTH 0.33 ;
  AREA 0.1518 RECTWIDTH 0.36 ;
  AREA 0.1641 RECTWIDTH 0.38 ;
  AREA 0.1681 RECTWIDTH 0.41 ;
 " ;
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 5000 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 3000  ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 10000 ;

END m7



#################################################
# Layer definition : v7
#################################################
LAYER v7
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS Via7_120Ux200 WIDTH 0.1200 LENGTH 0.2000 ;
  CUTCLASS Via7_120x400 WIDTH 0.1200 LENGTH 0.4000 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------
PROPERTY LEF58_ENCLOSURETABLE "
  ENCLOSURETABLE CUTCLASS Via7_120Ux200 
  WIDTH 0.181 ABOVE  0.0300 0.0300 0.0600 0.0600 INCLUDEABUTTED  ;
 " ;

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 0.24 ; # v7_Vyb_33 ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                          Via spacing table for vias on the same metal segment (SAMEMETAL)                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | v7_Vyb_33 | 0.2400     | v7-to-v7 spacing (edges), minimum, all-directional check                                   |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.2400 
   CUTCLASS                 Via7_120Ux200 SIDE     Via7_120Ux200 END         Via7_120x400 SIDE      Via7_120x400 END       
   Via7_120Ux200 SIDE       -       -              -       -                 -       -              -       -              
   Via7_120Ux200 END        -       -              -       -                 -       -              -       -              
   Via7_120x400 SIDE        -       -              -       -                 -       -              -       -              
   Via7_120x400 END         -       -              -       -                 -       -              -       -              
  ; " ;
 # -----------------------------------------------------------
 # No clr table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No clr_samenet table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No stack table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 550 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 550 ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 550 ;

END v7








#################################################
# Layer definition : m8
#################################################
LAYER m8
 TYPE ROUTING ;
 DIRECTION HORIZONTAL ;
 # ------------------------------------------------------------------
 # Width 
 # ------------------------------------------------------------------
 WIDTH    0.1800 ;
 MINWIDTH 0.18 ; # m8_Myb_01 ;
 MAXWIDTH 0.9 ; # m8_Myb_21 ;
 PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
 # ------------------------------------------------------------------
 # Spacing
 # ------------------------------------------------------------------
 SPACING  0.18 ; # m8_Myb_02 ;
 PITCH    0.3600 ; # WIDTH + SPACING 
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                     Metal end-to-end spacing for aligned lines                                      |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m8_Myb_03 | 0.2400     | Min m8 space (end-to-end, attacker). Applies to segments identified as line ends.          |
 # | m8_Myb_21 | 0.9000     | m8 width allowed range, maximum                                                            |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.2400 ENDOFLINE  0.9010 WRONGDIRSPACING 0.001  WITHIN 0.0010  ; " ;
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # |                                        Metal concave and convex corner rules                                        |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name | Rule Value | Rule Description                                                                           |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 # | m8_Myb_27 | 0.3080     | Minimum length of at least one segment, when two segments are adjacent at a corner         |
 # +-----------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_MINSTEP "
  MINSTEP 0.3080 MAXEDGES 1 MINADJACENTLENGTH 0.3080 CONCAVECORNER ;
  MINSTEP 0.3080 MAXEDGES 1 MINBETWEENLENGTH 0.3080   ;
 " ;

 # ------------------------------------------------------------------
 # Area and size
 # ------------------------------------------------------------------
 AREA     0.09000000 ; # m8_Myb_24 ;
 PROPERTY LEF58_AREA "
  AREA 0.09 RECTWIDTH 0.18 ;
  AREA 0.1074 RECTWIDTH 0.24 ;
  AREA 0.1195 RECTWIDTH 0.27 ;
  AREA 0.1317 RECTWIDTH 0.23 ;
  AREA 0.1438 RECTWIDTH 0.33 ;
  AREA 0.1518 RECTWIDTH 0.36 ;
  AREA 0.1641 RECTWIDTH 0.38 ;
  AREA 0.1681 RECTWIDTH 0.41 ;
 " ;
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 5000 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 3000  ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 10000 ;

END m8



#################################################
# Layer definition : v8
#################################################
LAYER v8
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS Via8_200x120 WIDTH 0.1200 LENGTH 0.2000 ;
  CUTCLASS Via8_400x120 WIDTH 0.1200 LENGTH 0.4000 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 0.24 ; # v8_Vybga_33 ;
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # |                           Via spacing table for vias on the same metal segment (SAMEMETAL)                            |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name   | Rule Value | Rule Description                                                                           |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 # | v8_Vybga_33 | 0.2400     | v8-to-v8 spacing (edges), minimum, all-directional check                                   |
 # +-------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.2400 
   CUTCLASS                Via8_200x120 SIDE     Via8_200x120 END      Via8_400x120 SIDE     Via8_400x120 END      
   Via8_200x120 SIDE       -       -             -       -             -       -             -       -             
   Via8_200x120 END        -       -             -       -             -       -             -       -             
   Via8_400x120 SIDE       -       -             -       -             -       -             -       -             
   Via8_400x120 END        -       -             -       -             -       -             -       -             
  ; " ;
 # -----------------------------------------------------------
 # No clr table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No clr_samenet table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No stack table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 550 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 550 ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 550 ;

END v8



 



#################################################
# Layer definition : gmz
#################################################
LAYER gmz
 TYPE ROUTING ;
 DIRECTION VERTICAL ;
 # ------------------------------------------------------------------
 # Width 
 # ------------------------------------------------------------------
 WIDTH    0.5400 ;
 MINWIDTH 0.54 ; # gmz_Mga_01 ;
 MAXWIDTH 7 ; # gmz_Mga_21 ;
 # ------------------------------------------------------------------
 # Spacing
 # ------------------------------------------------------------------
 SPACING  0.54 ; # gmz_Mga_02 ;
 PITCH    1.0800 ; # WIDTH + SPACING 
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # |                                      Metal end-to-end spacing for aligned lines                                      |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name  | Rule Value | Rule Description                                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | gmz_Mga_02 | 0.5400     | Min gmz space (side-to-side, end-to-end, attacker, all types)                              |
 # | gmz_Mga_21 | 7.0000     | gmz width allowed range, maximum                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.5400 ENDOFLINE  7.0010 WRONGDIRSPACING 0.001  WITHIN 0.0010  ; " ;
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # |                                        Metal concave and convex corner rules                                         |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name  | Rule Value | Rule Description                                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | gmz_Mga_27 | 0.5400     | Minimum length of at least one segment, when two segments are adjacent at a corner         |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_MINSTEP "
  MINSTEP 0.5400 MAXEDGES 1 MINADJACENTLENGTH 0.5400 CONCAVECORNER ;
 " ;

 # ------------------------------------------------------------------
 # Area and size
 # ------------------------------------------------------------------
 AREA     1.15020000 ; # gmz_Mga_01 * gmz_Mga_23 ;
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 5000 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 3000  ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 10000 ;

END gmz



#################################################
# Layer definition : vmz
#################################################
LAYER vmz
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS VMZ_120x200  WIDTH 0.1200 LENGTH 0.2000 ;
  CUTCLASS VMZ_120x400  WIDTH 0.1200 LENGTH 0.4000 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 0.24 ; # vmz_Vga_33 ;
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # |                           Via spacing table for vias on the same metal segment (SAMEMETAL)                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name  | Rule Value | Rule Description                                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | vmz_Vga_33 | 0.2400     | vmz-to-vmz spacing (edges), minimum, all-directional check                                 |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 0.2400 
   CUTCLASS               VMZ_120x200 SIDE     VMZ_120x200 END      VMZ_120x400 SIDE     VMZ_120x400 END      
   VMZ_120x200 SIDE       -       -            -       -            -       -            -       -            
   VMZ_120x200 END        -       -            -       -            -       -            -       -            
   VMZ_120x400 SIDE       -       -            -       -            -       -            -       -            
   VMZ_120x400 END        -       -            -       -            -       -            -       -            
  ; " ;
 # -----------------------------------------------------------
 # No clr table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No clr_samenet table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No stack table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 550 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 550 ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 550 ;

END vmz








#################################################
# Layer definition : gm0
#################################################
LAYER gm0
 TYPE ROUTING ;
 DIRECTION HORIZONTAL ;
 # ------------------------------------------------------------------
 # Width 
 # ------------------------------------------------------------------
 WIDTH    0.5400 ;
 MINWIDTH 0.54 ; # gm0_Mga_01 ;
 MAXWIDTH 7 ; # gm0_Mga_21 ;
 # ------------------------------------------------------------------
 # Spacing
 # ------------------------------------------------------------------
 SPACING  0.54 ; # gm0_Mga_02 ;
 PITCH    1.0800 ; # WIDTH + SPACING 
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # |                                      Metal end-to-end spacing for aligned lines                                      |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name  | Rule Value | Rule Description                                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | gm0_Mga_02 | 0.5400     | Min gmz space (side-to-side, end-to-end, attacker, all types)                              |
 # | gm0_Mga_21 | 7.0000     | gmz width allowed range, maximum                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 0.5400 ENDOFLINE  7.0010 WRONGDIRSPACING 0.001  WITHIN 0.0010  ; " ;
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # |                                        Metal concave and convex corner rules                                         |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name  | Rule Value | Rule Description                                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | gm0_Mga_27 | 0.5400     | Minimum length of at least one segment, when two segments are adjacent at a corner         |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_MINSTEP "
  MINSTEP 0.5400 MAXEDGES 1 MINADJACENTLENGTH 0.5400 CONCAVECORNER ;
 " ;

 # ------------------------------------------------------------------
 # Area and size
 # ------------------------------------------------------------------
 AREA     1.15020000 ; # gm0_Mga_01 * gm0_Mga_23 ;
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 5000 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 3000  ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 10000 ;

END gm0



#################################################
# Layer definition : gv0
#################################################
LAYER gv0
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS GV0_1850x800 WIDTH 0.8000 LENGTH 1.8500 ;
  CUTCLASS GV0_3700x800 WIDTH 0.8000 LENGTH 3.7000 ;
  CUTCLASS GV0_7400x800 WIDTH 0.8000 LENGTH 7.4000 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 2 ; # gv0_Vgagb_40 ;
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # |                            Via spacing table for vias on the same metal segment (SAMEMETAL)                            |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name    | Rule Value | Rule Description                                                                           |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 # | gv0_Vgagb_40 | 2.0000     | gv0-to-gv0 spacing between facing edges                                                    |
 # | gv0_Vgagb_41 | 2.5000     | gv0-to-gv0 corner-to-corner space (no facing edges)                                        |
 # +--------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 2.5000 
   CUTCLASS                GV0_1850x800 SIDE     GV0_1850x800 END      GV0_3700x800 SIDE     GV0_3700x800 END      GV0_7400x800 SIDE     GV0_7400x800 END      
   GV0_1850x800 SIDE       -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        
   GV0_1850x800 END        -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        
   GV0_3700x800 SIDE       -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        
   GV0_3700x800 END        -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        
   GV0_7400x800 SIDE       -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        
   GV0_7400x800 END        -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        -       2.0000        
  ; " ;
 # -----------------------------------------------------------
 # No clr table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No clr_samenet table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No stack table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------
 ANTENNAMODEL OXIDE1 ;
 ANTENNAAREARATIO 550 ;
 ANTENNAMODEL OXIDE2 ;
 ANTENNAAREARATIO 550 ;
 ANTENNAMODEL OXIDE3 ;
 ANTENNAAREARATIO 550 ;

END gv0




#################################################
# Layer definition : CE1
#################################################
LAYER CE1
 TYPE ROUTING ;
 PROPERTY LEF58_TYPE "TYPE STACKEDMIMCAP ;" ;
 DIRECTION VERTICAL ;
 PITCH 3 ; # MIM_01 + MIM_02 ;
 WIDTH 2 ; # MIM_01 ;
 MINWIDTH 2 ; # MIM_01 ;
 SPACING 1 ; # MIM_02 ;
END CE1



 

#################################################
# Layer definition : CE2
#################################################
LAYER CE2
 TYPE ROUTING ;
 PROPERTY LEF58_TYPE "TYPE STACKEDMIMCAP ;" ;
 DIRECTION VERTICAL ;
 PITCH 3 ; # MIM_01 + MIM_02 ;
 WIDTH 2 ; # MIM_01 ;
 MINWIDTH 2 ; # MIM_01 ;
 SPACING 1 ; # MIM_02 ;
END CE2





#################################################
# Layer definition : gmb
#################################################
LAYER gmb
 TYPE ROUTING ;
 DIRECTION VERTICAL ;
 # ------------------------------------------------------------------
 # Width 
 # ------------------------------------------------------------------
 WIDTH    1.0000 ;
 MINWIDTH 1 ; # gmb_Mgb_01 ;
 MAXWIDTH 12 ; # gmb_Mgb_21 ;
 # ------------------------------------------------------------------
 # Spacing
 # ------------------------------------------------------------------
 SPACING  1 ; # gmb_Mgb_02 ;
 PITCH    2.0000 ; # WIDTH + SPACING 
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # |                                      Metal end-to-end spacing for aligned lines                                      |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name  | Rule Value | Rule Description                                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | gmb_Mgb_02 | 1.0000     | gmb space (all directions), minimum                                                        |
 # | gmb_Mgb_21 | 12.0000    | gmb width allowed range, maximum                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACING "SPACING 1.0000 ENDOFLINE  12.0010 WRONGDIRSPACING 0.001  WITHIN 0.0010  ; " ;
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # |                                        Metal concave and convex corner rules                                         |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name  | Rule Value | Rule Description                                                                           |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 # | gmb_Mgb_27 | 0.5400     | Minimum length of at least one segment, when two segments are adjacent at a corner         |
 # +------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_MINSTEP "
  MINSTEP 0.5400 MAXEDGES 1 MINADJACENTLENGTH 0.5400 CONCAVECORNER ;
 " ;

 # ------------------------------------------------------------------
 # Area and size
 # ------------------------------------------------------------------
 AREA     4.84000000 ; # gmb_Mgb_01 * gmb_Mgb_23 ;
 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------


END gmb



#################################################
# Layer definition : gv1
#################################################
LAYER gv1
 TYPE CUT ;
 # ------------------------------------------------------------------
 # Cutclass definitions
 # ------------------------------------------------------------------
 PROPERTY LEF58_CUTCLASS "
  CUTCLASS GV1_6000x10000 WIDTH 6.0000 LENGTH 10.0000 ;
  CUTCLASS GV1_6000x18000 WIDTH 6.0000 LENGTH 18.0000 ;
  CUTCLASS GV1_6000x30000 WIDTH 6.0000 LENGTH 30.0000 ;
 " ;
 # ------------------------------------------------------------------
 # Enclosure definitions
 # ------------------------------------------------------------------

 # ------------------------------------------------------------------
 # Spacing definitions
 # ------------------------------------------------------------------
 SPACING 37 ; # c4_Bumpp55_102 - xSize/2 of GV1_18000x6000 - xSize/2 of GV1_18000x6000 ;
 # +--------------------------------------------------------------------------------+------------+--------------------------------------------------------------------------------------------+
 # |                                                             Via spacing table for vias on the same metal segment (SAMEMETAL)                                                             |
 # +--------------------------------------------------------------------------------+------------+--------------------------------------------------------------------------------------------+
 # | Rule Name                                                                      | Rule Value | Rule Description                                                                           |
 # +--------------------------------------------------------------------------------+------------+--------------------------------------------------------------------------------------------+
 # | c4_Bumpp55_102 - sqrt((v1.x/2)^2 + (v1.y/2)^2) - sqrt((v2.x/2)^2 + (v2.y/2)^2) | 43.3381    |                                                                                            |
 # | c4_Bumpp55_102 - xSize/2 of GV1_6000x10000 - xSize/2 of GV1_6000x10000         | 49.0000    |                                                                                            |
 # | c4_Bumpp55_102 - xSize/2 of GV1_6000x10000 - xSize/2 of GV1_6000x18000         | 49.0000    |                                                                                            |
 # | c4_Bumpp55_102 - xSize/2 of GV1_6000x18000 - xSize/2 of GV1_6000x10000         | 49.0000    |                                                                                            |
 # | c4_Bumpp55_102 - xSize/2 of GV1_6000x18000 - xSize/2 of GV1_6000x18000         | 49.0000    |                                                                                            |
 # | c4_Bumpp55_102 - ySize/2 of GV1_6000x10000 - ySize/2 of GV1_6000x10000         | 45.0000    |                                                                                            |
 # | c4_Bumpp55_102 - ySize/2 of GV1_6000x10000 - ySize/2 of GV1_6000x18000         | 41.0000    |                                                                                            |
 # | c4_Bumpp55_102 - ySize/2 of GV1_6000x18000 - ySize/2 of GV1_6000x10000         | 41.0000    |                                                                                            |
 # | c4_Bumpp55_102 - ySize/2 of GV1_6000x18000 - ySize/2 of GV1_6000x18000         | 37.0000    |                                                                                            |
 # | c4_Bumpp_406 - sqrt((v1.x/2)^2 + (v1.y/2)^2) - sqrt((v2.x/2)^2 + (v2.y/2)^2)   | 79.1720    |                                                                                            |
 # | c4_Bumpp_406 - xSize/2 of GV1_6000x10000 - xSize/2 of GV1_6000x30000           | 94.3000    |                                                                                            |
 # | c4_Bumpp_406 - xSize/2 of GV1_6000x18000 - xSize/2 of GV1_6000x30000           | 94.3000    |                                                                                            |
 # | c4_Bumpp_406 - xSize/2 of GV1_6000x30000 - xSize/2 of GV1_6000x10000           | 94.3000    |                                                                                            |
 # | c4_Bumpp_406 - xSize/2 of GV1_6000x30000 - xSize/2 of GV1_6000x18000           | 94.3000    |                                                                                            |
 # | c4_Bumpp_406 - xSize/2 of GV1_6000x30000 - xSize/2 of GV1_6000x30000           | 94.3000    |                                                                                            |
 # | c4_Bumpp_406 - ySize/2 of GV1_6000x10000 - ySize/2 of GV1_6000x30000           | 80.3000    |                                                                                            |
 # | c4_Bumpp_406 - ySize/2 of GV1_6000x18000 - ySize/2 of GV1_6000x30000           | 76.3000    |                                                                                            |
 # | c4_Bumpp_406 - ySize/2 of GV1_6000x30000 - ySize/2 of GV1_6000x10000           | 80.3000    |                                                                                            |
 # | c4_Bumpp_406 - ySize/2 of GV1_6000x30000 - ySize/2 of GV1_6000x18000           | 76.3000    |                                                                                            |
 # | c4_Bumpp_406 - ySize/2 of GV1_6000x30000 - ySize/2 of GV1_6000x30000           | 70.3000    |                                                                                            |
 # +--------------------------------------------------------------------------------+------------+--------------------------------------------------------------------------------------------+
 PROPERTY LEF58_SPACINGTABLE "
  SPACINGTABLE DEFAULT 69.7059 
   CUTCLASS                  GV1_6000x10000 SIDE     GV1_6000x10000 END      GV1_6000x18000 SIDE     GV1_6000x18000 END      GV1_6000x30000 SIDE     GV1_6000x30000 END      
   GV1_6000x10000 SIDE       43.3381 49.0000         43.3381 -               39.6822 49.0000         39.6822 -               -       94.3000         -       -               
   GV1_6000x10000 END        43.3381 -               43.3381 45.0000         39.6822 -               39.6822 41.0000         -       -               -       80.3000         
   GV1_6000x18000 SIDE       39.6822 49.0000         39.6822 -               36.0263 49.0000         36.0263 -               -       94.3000         -       -               
   GV1_6000x18000 END        39.6822 -               39.6822 41.0000         36.0263 -               36.0263 37.0000         -       -               -       76.3000         
   GV1_6000x30000 SIDE       -       94.3000         -       -               -       94.3000         -       -               -       94.3000         -       -               
   GV1_6000x30000 END        -       -               -       80.3000         -       -               -       76.3000         -       -               -       70.3000         
  ; " ;
 # -----------------------------------------------------------
 # No clr table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No clr_samenet table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # -----------------------------------------------------------
 # No stack table (Vn to Vn-1) required 
 # -----------------------------------------------------------

 # ------------------------------------------------------------------
 # Antenna definitions
 # ------------------------------------------------------------------


END gv1





#################################################
# Layer definition : c4
#################################################
LAYER c4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PROPERTY LEF58_WIDTHTABLE "WIDTHTABLE 51.0 54.0 85.0 ;" ;
  PITCH 100.3 ; # c4_Bumpp45_412 + c4_Bumpp_406 - c4_Bumpp45_412 ;
  WIDTH 51 ; # c4_Bumpp45_412 ;
  MINWIDTH 51 ; # c4_Bumpp45_412 ;
  SPACING 49.3 ; # c4_Bumpp_406 - c4_Bumpp45_412 ;
END c4

#################################################
# Layer definition : c4emib
#################################################
LAYER c4emib
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PROPERTY LEF58_WIDTHTABLE "WIDTHTABLE 20.0 28.0 ;" ;
  PROPERTY LEF58_TYPE "TYPE MIMCAP ;" ;
  PITCH 55 ; # c4_Bumpp45_101 + c4_Bumpp55_102 - c4_Bumpp45_101 ;
  WIDTH 20 ; # c4_Bumpp45_101 ;
  MINWIDTH 20 ; # c4_Bumpp45_101 ;
  SPACING 35 ; # c4_Bumpp55_102 - c4_Bumpp45_101 ;
END c4emib


##################################################
# Via Definitions
##################################################

# |-------------------------------------------------------------------------------------------|
# | Via Naming Convention: [viaLayer]_[cutSize]_[lowerMetal]_[UpperMetal]                     |
# |-------------------------------------------------------------------------------------------|
# |  viaLayer   | viaL      | Via cut layer with lowercase "via" and integer (ex: via1, via2) |
# |             |           |    via = lowercase "via" string indicating via definition       |
# |             |           |    L = via cut layer                                            |
# |-------------|-----------|-----------------------------------------------------------------|
# |  cutSize    | N{S}xM{S} | Via cutclass size N by M with lowercase "x" and                 |
# |             |           | including self aligned "S" on one side                          |
# |             |           |    N = via cut N dimension                                      |
# |             |           |    M = via cut M dimension                                      |
# |             |           |    x = lowercase "x" separating N and M                         |
# |             |           |    S = self aligned side on either the N or M side              |
# |-------------|-----------|-----------------------------------------------------------------|
# |  lowerMetal | W{HV}     | Lower metal layer width and uppercase direction indication      |
# |             |           |    W = integer width in nm                                      |
# |             |           |    H = horizontal metal direction                               |
# |             |           |    V = vertical metal direction                                 |
# |-------------|-----------|-----------------------------------------------------------------|
# |  upperMetal | W{HV}     | Upper metal layer width and uppercase direction indication      |
# |             |           |    W = integer width in nm                                      |
# |             |           |    H = horizontal                                               |
# |             |           |    V = vertical                                                 |
# |-------------------------------------------------------------------------------------------|
# |  NOTES                                                                                    |
# |-------------------------------------------------------------------------------------------|
# |  1.  Vias connecting preferred direction layers to each other and will                    |
# |      have an "H" width and a "V" width in the name (via1_60Sx44_68V_44H)                  |
# |-------------------------------------------------------------------------------------------|
# |  2.  Vias connecting non-preferred direction metal layers can have a name with            |
# |      two "H" widths (via7_68Sx60_68H_60H) or two "V" widths (via7_68Sx60_60V_68V)         |
# |                                                                                           |
# |-------------------------------------------------------------------------------------------|
# | Example     | via1_60Sx44_68V_44H                                                         |
# |-------------|-----------------------------------------------------------------------------|
# |  via1       | Via cut layer 1                                                             |
# |  60Sx44     | Via cut specified Via1_60Sx44                                               |
# |  68V        | 68nm vertical metal width (M1 in this case)                                 |
# |  44H        | 44nm horizontal metal width (M2 in this case)                               |
# |-------------------------------------------------------------------------------------------|

VIA VIA1_60SX44_68V_44H
  # v1   size: x=0.0600 y=0.0440
  # m1   size: x=0.0680 y=0.0440   enclosure: x=0.0040 y=0.0000
  # m2   size: x=0.1040 y=0.0440   enclosure: x=0.0220 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.0340 -0.0220 0.0340 0.0220 ;
  LAYER v1   ; RECT -0.0300 -0.0220 0.0300 0.0220 ;
  LAYER m2   ; RECT -0.0520 -0.0220 0.0520 0.0220 ;
END VIA1_60SX44_68V_44H

VIA VIA1_60SX56_68V_56H
  # v1   size: x=0.0600 y=0.0560
  # m1   size: x=0.0680 y=0.0760   enclosure: x=0.0040 y=0.0100
  # m2   size: x=0.1040 y=0.0560   enclosure: x=0.0220 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.0340 -0.0380 0.0340 0.0380 ;
  LAYER v1   ; RECT -0.0300 -0.0280 0.0300 0.0280 ;
  LAYER m2   ; RECT -0.0520 -0.0280 0.0520 0.0280 ;
END VIA1_60SX56_68V_56H

VIA VIA1_60SX76_68V_76H
  # v1   size: x=0.0600 y=0.0760
  # m1   size: x=0.0680 y=0.0960   enclosure: x=0.0040 y=0.0100
  # m2   size: x=0.1040 y=0.0760   enclosure: x=0.0220 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.0340 -0.0480 0.0340 0.0480 ;
  LAYER v1   ; RECT -0.0300 -0.0380 0.0300 0.0380 ;
  LAYER m2   ; RECT -0.0520 -0.0380 0.0520 0.0380 ;
END VIA1_60SX76_68V_76H

VIA VIA1_60SX90_68V_90H
  # v1   size: x=0.0600 y=0.0900
  # m1   size: x=0.0680 y=0.1100   enclosure: x=0.0040 y=0.0100
  # m2   size: x=0.1040 y=0.0900   enclosure: x=0.0220 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.0340 -0.0550 0.0340 0.0550 ;
  LAYER v1   ; RECT -0.0300 -0.0450 0.0300 0.0450 ;
  LAYER m2   ; RECT -0.0520 -0.0450 0.0520 0.0450 ;
END VIA1_60SX90_68V_90H

VIA VIA1_60SX108_68V_108H
  # v1   size: x=0.0600 y=0.1080
  # m1   size: x=0.0680 y=0.1280   enclosure: x=0.0040 y=0.0100
  # m2   size: x=0.1040 y=0.1080   enclosure: x=0.0220 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.0340 -0.0640 0.0340 0.0640 ;
  LAYER v1   ; RECT -0.0300 -0.0540 0.0300 0.0540 ;
  LAYER m2   ; RECT -0.0520 -0.0540 0.0520 0.0540 ;
END VIA1_60SX108_68V_108H

VIA VIA1_60SX44_100V_44H
  # v1   size: x=0.0600 y=0.0440
  # m1   size: x=0.1000 y=0.0640   enclosure: x=0.0200 y=0.0100
  # m2   size: x=0.1040 y=0.0440   enclosure: x=0.0220 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.0500 -0.0320 0.0500 0.0320 ;
  LAYER v1   ; RECT -0.0300 -0.0220 0.0300 0.0220 ;
  LAYER m2   ; RECT -0.0520 -0.0220 0.0520 0.0220 ;
END VIA1_60SX44_100V_44H

VIA VIA1_60SX56_100V_56H
  # v1   size: x=0.0600 y=0.0560
  # m1   size: x=0.1000 y=0.0760   enclosure: x=0.0200 y=0.0100
  # m2   size: x=0.1040 y=0.0560   enclosure: x=0.0220 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
  LAYER v1   ; RECT -0.0300 -0.0280 0.0300 0.0280 ;
  LAYER m2   ; RECT -0.0520 -0.0280 0.0520 0.0280 ;
END VIA1_60SX56_100V_56H

VIA VIA1_60SX76_100V_76H
  # v1   size: x=0.0600 y=0.0760
  # m1   size: x=0.1000 y=0.0960   enclosure: x=0.0200 y=0.0100
  # m2   size: x=0.1040 y=0.0760   enclosure: x=0.0220 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.0500 -0.0480 0.0500 0.0480 ;
  LAYER v1   ; RECT -0.0300 -0.0380 0.0300 0.0380 ;
  LAYER m2   ; RECT -0.0520 -0.0380 0.0520 0.0380 ;
END VIA1_60SX76_100V_76H

VIA VIA1_60SX90_100V_90H
  # v1   size: x=0.0600 y=0.0900
  # m1   size: x=0.1000 y=0.1100   enclosure: x=0.0200 y=0.0100
  # m2   size: x=0.1040 y=0.0900   enclosure: x=0.0220 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.0500 -0.0550 0.0500 0.0550 ;
  LAYER v1   ; RECT -0.0300 -0.0450 0.0300 0.0450 ;
  LAYER m2   ; RECT -0.0520 -0.0450 0.0520 0.0450 ;
END VIA1_60SX90_100V_90H

VIA VIA1_60SX108_100V_108H
  # v1   size: x=0.0600 y=0.1080
  # m1   size: x=0.1000 y=0.1280   enclosure: x=0.0200 y=0.0100
  # m2   size: x=0.1040 y=0.1080   enclosure: x=0.0220 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.0500 -0.0640 0.0500 0.0640 ;
  LAYER v1   ; RECT -0.0300 -0.0540 0.0300 0.0540 ;
  LAYER m2   ; RECT -0.0520 -0.0540 0.0520 0.0540 ;
END VIA1_60SX108_100V_108H

VIA VIA2_44X58S_44H_44V
  # v2   size: x=0.0440 y=0.0580
  # m2   size: x=0.0680 y=0.0440   enclosure: x=0.0120 y=-0.0070
  # m3   size: x=0.0440 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0340 -0.0220 0.0340 0.0220 ;
  LAYER v2   ; RECT -0.0220 -0.0290 0.0220 0.0290 ;
  LAYER m3   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
END VIA2_44X58S_44H_44V

VIA VIA2_56X58S_44H_56V
  # v2   size: x=0.0560 y=0.0580
  # m2   size: x=0.0800 y=0.0440   enclosure: x=0.0120 y=-0.0070
  # m3   size: x=0.0560 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0400 -0.0220 0.0400 0.0220 ;
  LAYER v2   ; RECT -0.0280 -0.0290 0.0280 0.0290 ;
  LAYER m3   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
END VIA2_56X58S_44H_56V

VIA VIA2_76X58S_44H_76V
  # v2   size: x=0.0760 y=0.0580
  # m2   size: x=0.1000 y=0.0440   enclosure: x=0.0120 y=-0.0070
  # m3   size: x=0.0760 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
  LAYER v2   ; RECT -0.0380 -0.0290 0.0380 0.0290 ;
  LAYER m3   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
END VIA2_76X58S_44H_76V

VIA VIA2_90X58S_44H_90V
  # v2   size: x=0.0900 y=0.0580
  # m2   size: x=0.1140 y=0.0440   enclosure: x=0.0120 y=-0.0070
  # m3   size: x=0.0900 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0570 -0.0220 0.0570 0.0220 ;
  LAYER v2   ; RECT -0.0450 -0.0290 0.0450 0.0290 ;
  LAYER m3   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
END VIA2_90X58S_44H_90V

VIA VIA2_108X58S_44H_108V
  # v2   size: x=0.1080 y=0.0580
  # m2   size: x=0.1320 y=0.0440   enclosure: x=0.0120 y=-0.0070
  # m3   size: x=0.1080 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0660 -0.0220 0.0660 0.0220 ;
  LAYER v2   ; RECT -0.0540 -0.0290 0.0540 0.0290 ;
  LAYER m3   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
END VIA2_108X58S_44H_108V

VIA VIA2_44X58S_56H_44V
  # v2   size: x=0.0440 y=0.0580
  # m2   size: x=0.0680 y=0.0560   enclosure: x=0.0120 y=-0.0010
  # m3   size: x=0.0440 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0340 -0.0280 0.0340 0.0280 ;
  LAYER v2   ; RECT -0.0220 -0.0290 0.0220 0.0290 ;
  LAYER m3   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
END VIA2_44X58S_56H_44V

VIA VIA2_56X58S_56H_56V
  # v2   size: x=0.0560 y=0.0580
  # m2   size: x=0.0800 y=0.0560   enclosure: x=0.0120 y=-0.0010
  # m3   size: x=0.0560 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0400 -0.0280 0.0400 0.0280 ;
  LAYER v2   ; RECT -0.0280 -0.0290 0.0280 0.0290 ;
  LAYER m3   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
END VIA2_56X58S_56H_56V

VIA VIA2_76X58S_56H_76V
  # v2   size: x=0.0760 y=0.0580
  # m2   size: x=0.1000 y=0.0560   enclosure: x=0.0120 y=-0.0010
  # m3   size: x=0.0760 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
  LAYER v2   ; RECT -0.0380 -0.0290 0.0380 0.0290 ;
  LAYER m3   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
END VIA2_76X58S_56H_76V

VIA VIA2_90X58S_56H_90V
  # v2   size: x=0.0900 y=0.0580
  # m2   size: x=0.1140 y=0.0560   enclosure: x=0.0120 y=-0.0010
  # m3   size: x=0.0900 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0570 -0.0280 0.0570 0.0280 ;
  LAYER v2   ; RECT -0.0450 -0.0290 0.0450 0.0290 ;
  LAYER m3   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
END VIA2_90X58S_56H_90V

VIA VIA2_108X58S_56H_108V
  # v2   size: x=0.1080 y=0.0580
  # m2   size: x=0.1320 y=0.0560   enclosure: x=0.0120 y=-0.0010
  # m3   size: x=0.1080 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0660 -0.0280 0.0660 0.0280 ;
  LAYER v2   ; RECT -0.0540 -0.0290 0.0540 0.0290 ;
  LAYER m3   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
END VIA2_108X58S_56H_108V

VIA VIA2_44X58S_76H_44V
  # v2   size: x=0.0440 y=0.0580
  # m2   size: x=0.0680 y=0.0760   enclosure: x=0.0120 y=0.0090
  # m3   size: x=0.0440 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0340 -0.0380 0.0340 0.0380 ;
  LAYER v2   ; RECT -0.0220 -0.0290 0.0220 0.0290 ;
  LAYER m3   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
END VIA2_44X58S_76H_44V

VIA VIA2_56X58S_76H_56V
  # v2   size: x=0.0560 y=0.0580
  # m2   size: x=0.0800 y=0.0760   enclosure: x=0.0120 y=0.0090
  # m3   size: x=0.0560 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0400 -0.0380 0.0400 0.0380 ;
  LAYER v2   ; RECT -0.0280 -0.0290 0.0280 0.0290 ;
  LAYER m3   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
END VIA2_56X58S_76H_56V

VIA VIA2_76X58S_76H_76V
  # v2   size: x=0.0760 y=0.0580
  # m2   size: x=0.1000 y=0.0760   enclosure: x=0.0120 y=0.0090
  # m3   size: x=0.0760 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
  LAYER v2   ; RECT -0.0380 -0.0290 0.0380 0.0290 ;
  LAYER m3   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
END VIA2_76X58S_76H_76V

VIA VIA2_90X58S_76H_90V
  # v2   size: x=0.0900 y=0.0580
  # m2   size: x=0.1140 y=0.0760   enclosure: x=0.0120 y=0.0090
  # m3   size: x=0.0900 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0570 -0.0380 0.0570 0.0380 ;
  LAYER v2   ; RECT -0.0450 -0.0290 0.0450 0.0290 ;
  LAYER m3   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
END VIA2_90X58S_76H_90V

VIA VIA2_108X58S_76H_108V
  # v2   size: x=0.1080 y=0.0580
  # m2   size: x=0.1320 y=0.0760   enclosure: x=0.0120 y=0.0090
  # m3   size: x=0.1080 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0660 -0.0380 0.0660 0.0380 ;
  LAYER v2   ; RECT -0.0540 -0.0290 0.0540 0.0290 ;
  LAYER m3   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
END VIA2_108X58S_76H_108V

VIA VIA2_44X58S_90H_44V
  # v2   size: x=0.0440 y=0.0580
  # m2   size: x=0.0680 y=0.0900   enclosure: x=0.0120 y=0.0160
  # m3   size: x=0.0440 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0340 -0.0450 0.0340 0.0450 ;
  LAYER v2   ; RECT -0.0220 -0.0290 0.0220 0.0290 ;
  LAYER m3   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
END VIA2_44X58S_90H_44V

VIA VIA2_56X58S_90H_56V
  # v2   size: x=0.0560 y=0.0580
  # m2   size: x=0.0800 y=0.0900   enclosure: x=0.0120 y=0.0160
  # m3   size: x=0.0560 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0400 -0.0450 0.0400 0.0450 ;
  LAYER v2   ; RECT -0.0280 -0.0290 0.0280 0.0290 ;
  LAYER m3   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
END VIA2_56X58S_90H_56V

VIA VIA2_76X58S_90H_76V
  # v2   size: x=0.0760 y=0.0580
  # m2   size: x=0.1000 y=0.0900   enclosure: x=0.0120 y=0.0160
  # m3   size: x=0.0760 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
  LAYER v2   ; RECT -0.0380 -0.0290 0.0380 0.0290 ;
  LAYER m3   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
END VIA2_76X58S_90H_76V

VIA VIA2_90X58S_90H_90V
  # v2   size: x=0.0900 y=0.0580
  # m2   size: x=0.1140 y=0.0900   enclosure: x=0.0120 y=0.0160
  # m3   size: x=0.0900 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0570 -0.0450 0.0570 0.0450 ;
  LAYER v2   ; RECT -0.0450 -0.0290 0.0450 0.0290 ;
  LAYER m3   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
END VIA2_90X58S_90H_90V

VIA VIA2_108X58S_90H_108V
  # v2   size: x=0.1080 y=0.0580
  # m2   size: x=0.1320 y=0.0900   enclosure: x=0.0120 y=0.0160
  # m3   size: x=0.1080 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0660 -0.0450 0.0660 0.0450 ;
  LAYER v2   ; RECT -0.0540 -0.0290 0.0540 0.0290 ;
  LAYER m3   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
END VIA2_108X58S_90H_108V

VIA VIA2_44X58S_108H_44V
  # v2   size: x=0.0440 y=0.0580
  # m2   size: x=0.0680 y=0.1080   enclosure: x=0.0120 y=0.0250
  # m3   size: x=0.0440 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0340 -0.0540 0.0340 0.0540 ;
  LAYER v2   ; RECT -0.0220 -0.0290 0.0220 0.0290 ;
  LAYER m3   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
END VIA2_44X58S_108H_44V

VIA VIA2_56X58S_108H_56V
  # v2   size: x=0.0560 y=0.0580
  # m2   size: x=0.0800 y=0.1080   enclosure: x=0.0120 y=0.0250
  # m3   size: x=0.0560 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0400 -0.0540 0.0400 0.0540 ;
  LAYER v2   ; RECT -0.0280 -0.0290 0.0280 0.0290 ;
  LAYER m3   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
END VIA2_56X58S_108H_56V

VIA VIA2_76X58S_108H_76V
  # v2   size: x=0.0760 y=0.0580
  # m2   size: x=0.1000 y=0.1080   enclosure: x=0.0120 y=0.0250
  # m3   size: x=0.0760 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
  LAYER v2   ; RECT -0.0380 -0.0290 0.0380 0.0290 ;
  LAYER m3   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
END VIA2_76X58S_108H_76V

VIA VIA2_90X58S_108H_90V
  # v2   size: x=0.0900 y=0.0580
  # m2   size: x=0.1140 y=0.1080   enclosure: x=0.0120 y=0.0250
  # m3   size: x=0.0900 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0570 -0.0540 0.0570 0.0540 ;
  LAYER v2   ; RECT -0.0450 -0.0290 0.0450 0.0290 ;
  LAYER m3   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
END VIA2_90X58S_108H_90V

VIA VIA2_108X58S_108H_108V
  # v2   size: x=0.1080 y=0.0580
  # m2   size: x=0.1320 y=0.1080   enclosure: x=0.0120 y=0.0250
  # m3   size: x=0.1080 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.0660 -0.0540 0.0660 0.0540 ;
  LAYER v2   ; RECT -0.0540 -0.0290 0.0540 0.0290 ;
  LAYER m3   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
END VIA2_108X58S_108H_108V

VIA VIA3_58SX44_44V_44H
  # v3   size: x=0.0580 y=0.0440
  # m3   size: x=0.0440 y=0.0680   enclosure: x=-0.0070 y=0.0120
  # m4   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0220 -0.0340 0.0220 0.0340 ;
  LAYER v3   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m4   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA3_58SX44_44V_44H

VIA VIA3_58SX56_44V_56H
  # v3   size: x=0.0580 y=0.0560
  # m3   size: x=0.0440 y=0.0800   enclosure: x=-0.0070 y=0.0120
  # m4   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0220 -0.0400 0.0220 0.0400 ;
  LAYER v3   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m4   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA3_58SX56_44V_56H

VIA VIA3_58SX76_44V_76H
  # v3   size: x=0.0580 y=0.0760
  # m3   size: x=0.0440 y=0.1000   enclosure: x=-0.0070 y=0.0120
  # m4   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
  LAYER v3   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m4   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA3_58SX76_44V_76H

VIA VIA3_58SX90_44V_90H
  # v3   size: x=0.0580 y=0.0900
  # m3   size: x=0.0440 y=0.1140   enclosure: x=-0.0070 y=0.0120
  # m4   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0220 -0.0570 0.0220 0.0570 ;
  LAYER v3   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m4   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA3_58SX90_44V_90H

VIA VIA3_58SX108_44V_108H
  # v3   size: x=0.0580 y=0.1080
  # m3   size: x=0.0440 y=0.1320   enclosure: x=-0.0070 y=0.0120
  # m4   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0220 -0.0660 0.0220 0.0660 ;
  LAYER v3   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m4   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA3_58SX108_44V_108H

VIA VIA3_58SX44_56V_44H
  # v3   size: x=0.0580 y=0.0440
  # m3   size: x=0.0560 y=0.0680   enclosure: x=-0.0010 y=0.0120
  # m4   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0280 -0.0340 0.0280 0.0340 ;
  LAYER v3   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m4   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA3_58SX44_56V_44H

VIA VIA3_58SX56_56V_56H
  # v3   size: x=0.0580 y=0.0560
  # m3   size: x=0.0560 y=0.0800   enclosure: x=-0.0010 y=0.0120
  # m4   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0280 -0.0400 0.0280 0.0400 ;
  LAYER v3   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m4   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA3_58SX56_56V_56H

VIA VIA3_58SX76_56V_76H
  # v3   size: x=0.0580 y=0.0760
  # m3   size: x=0.0560 y=0.1000   enclosure: x=-0.0010 y=0.0120
  # m4   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
  LAYER v3   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m4   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA3_58SX76_56V_76H

VIA VIA3_58SX90_56V_90H
  # v3   size: x=0.0580 y=0.0900
  # m3   size: x=0.0560 y=0.1140   enclosure: x=-0.0010 y=0.0120
  # m4   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0280 -0.0570 0.0280 0.0570 ;
  LAYER v3   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m4   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA3_58SX90_56V_90H

VIA VIA3_58SX108_56V_108H
  # v3   size: x=0.0580 y=0.1080
  # m3   size: x=0.0560 y=0.1320   enclosure: x=-0.0010 y=0.0120
  # m4   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0280 -0.0660 0.0280 0.0660 ;
  LAYER v3   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m4   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA3_58SX108_56V_108H

VIA VIA3_58SX44_76V_44H
  # v3   size: x=0.0580 y=0.0440
  # m3   size: x=0.0760 y=0.0680   enclosure: x=0.0090 y=0.0120
  # m4   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0380 -0.0340 0.0380 0.0340 ;
  LAYER v3   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m4   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA3_58SX44_76V_44H

VIA VIA3_58SX56_76V_56H
  # v3   size: x=0.0580 y=0.0560
  # m3   size: x=0.0760 y=0.0800   enclosure: x=0.0090 y=0.0120
  # m4   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0380 -0.0400 0.0380 0.0400 ;
  LAYER v3   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m4   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA3_58SX56_76V_56H

VIA VIA3_58SX76_76V_76H
  # v3   size: x=0.0580 y=0.0760
  # m3   size: x=0.0760 y=0.1000   enclosure: x=0.0090 y=0.0120
  # m4   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
  LAYER v3   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m4   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA3_58SX76_76V_76H

VIA VIA3_58SX90_76V_90H
  # v3   size: x=0.0580 y=0.0900
  # m3   size: x=0.0760 y=0.1140   enclosure: x=0.0090 y=0.0120
  # m4   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0380 -0.0570 0.0380 0.0570 ;
  LAYER v3   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m4   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA3_58SX90_76V_90H

VIA VIA3_58SX108_76V_108H
  # v3   size: x=0.0580 y=0.1080
  # m3   size: x=0.0760 y=0.1320   enclosure: x=0.0090 y=0.0120
  # m4   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0380 -0.0660 0.0380 0.0660 ;
  LAYER v3   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m4   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA3_58SX108_76V_108H

VIA VIA3_58SX44_90V_44H
  # v3   size: x=0.0580 y=0.0440
  # m3   size: x=0.0900 y=0.0680   enclosure: x=0.0160 y=0.0120
  # m4   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0450 -0.0340 0.0450 0.0340 ;
  LAYER v3   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m4   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA3_58SX44_90V_44H

VIA VIA3_58SX56_90V_56H
  # v3   size: x=0.0580 y=0.0560
  # m3   size: x=0.0900 y=0.0800   enclosure: x=0.0160 y=0.0120
  # m4   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0450 -0.0400 0.0450 0.0400 ;
  LAYER v3   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m4   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA3_58SX56_90V_56H

VIA VIA3_58SX76_90V_76H
  # v3   size: x=0.0580 y=0.0760
  # m3   size: x=0.0900 y=0.1000   enclosure: x=0.0160 y=0.0120
  # m4   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
  LAYER v3   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m4   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA3_58SX76_90V_76H

VIA VIA3_58SX90_90V_90H
  # v3   size: x=0.0580 y=0.0900
  # m3   size: x=0.0900 y=0.1140   enclosure: x=0.0160 y=0.0120
  # m4   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0450 -0.0570 0.0450 0.0570 ;
  LAYER v3   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m4   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA3_58SX90_90V_90H

VIA VIA3_58SX108_90V_108H
  # v3   size: x=0.0580 y=0.1080
  # m3   size: x=0.0900 y=0.1320   enclosure: x=0.0160 y=0.0120
  # m4   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0450 -0.0660 0.0450 0.0660 ;
  LAYER v3   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m4   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA3_58SX108_90V_108H

VIA VIA3_58SX44_108V_44H
  # v3   size: x=0.0580 y=0.0440
  # m3   size: x=0.1080 y=0.0680   enclosure: x=0.0250 y=0.0120
  # m4   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0540 -0.0340 0.0540 0.0340 ;
  LAYER v3   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m4   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA3_58SX44_108V_44H

VIA VIA3_58SX56_108V_56H
  # v3   size: x=0.0580 y=0.0560
  # m3   size: x=0.1080 y=0.0800   enclosure: x=0.0250 y=0.0120
  # m4   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0540 -0.0400 0.0540 0.0400 ;
  LAYER v3   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m4   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA3_58SX56_108V_56H

VIA VIA3_58SX76_108V_76H
  # v3   size: x=0.0580 y=0.0760
  # m3   size: x=0.1080 y=0.1000   enclosure: x=0.0250 y=0.0120
  # m4   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
  LAYER v3   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m4   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA3_58SX76_108V_76H

VIA VIA3_58SX90_108V_90H
  # v3   size: x=0.0580 y=0.0900
  # m3   size: x=0.1080 y=0.1140   enclosure: x=0.0250 y=0.0120
  # m4   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0540 -0.0570 0.0540 0.0570 ;
  LAYER v3   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m4   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA3_58SX90_108V_90H

VIA VIA3_58SX108_108V_108H
  # v3   size: x=0.0580 y=0.1080
  # m3   size: x=0.1080 y=0.1320   enclosure: x=0.0250 y=0.0120
  # m4   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.0540 -0.0660 0.0540 0.0660 ;
  LAYER v3   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m4   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA3_58SX108_108V_108H

VIA VIA4_44X58S_44H_44V
  # v4   size: x=0.0440 y=0.0580
  # m4   size: x=0.0680 y=0.0440   enclosure: x=0.0120 y=-0.0070
  # m5   size: x=0.0440 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0340 -0.0220 0.0340 0.0220 ;
  LAYER v4   ; RECT -0.0220 -0.0290 0.0220 0.0290 ;
  LAYER m5   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
END VIA4_44X58S_44H_44V

VIA VIA4_56X58S_44H_56V
  # v4   size: x=0.0560 y=0.0580
  # m4   size: x=0.0800 y=0.0440   enclosure: x=0.0120 y=-0.0070
  # m5   size: x=0.0560 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0400 -0.0220 0.0400 0.0220 ;
  LAYER v4   ; RECT -0.0280 -0.0290 0.0280 0.0290 ;
  LAYER m5   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
END VIA4_56X58S_44H_56V

VIA VIA4_76X58S_44H_76V
  # v4   size: x=0.0760 y=0.0580
  # m4   size: x=0.1000 y=0.0440   enclosure: x=0.0120 y=-0.0070
  # m5   size: x=0.0760 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
  LAYER v4   ; RECT -0.0380 -0.0290 0.0380 0.0290 ;
  LAYER m5   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
END VIA4_76X58S_44H_76V

VIA VIA4_90X58S_44H_90V
  # v4   size: x=0.0900 y=0.0580
  # m4   size: x=0.1140 y=0.0440   enclosure: x=0.0120 y=-0.0070
  # m5   size: x=0.0900 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0570 -0.0220 0.0570 0.0220 ;
  LAYER v4   ; RECT -0.0450 -0.0290 0.0450 0.0290 ;
  LAYER m5   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
END VIA4_90X58S_44H_90V

VIA VIA4_108X58S_44H_108V
  # v4   size: x=0.1080 y=0.0580
  # m4   size: x=0.1320 y=0.0440   enclosure: x=0.0120 y=-0.0070
  # m5   size: x=0.1080 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0660 -0.0220 0.0660 0.0220 ;
  LAYER v4   ; RECT -0.0540 -0.0290 0.0540 0.0290 ;
  LAYER m5   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
END VIA4_108X58S_44H_108V

VIA VIA4_160X58S_44H_160V
  # v4   size: x=0.1600 y=0.0580
  # m4   size: x=0.1840 y=0.0440   enclosure: x=0.0120 y=-0.0070
  # m5   size: x=0.1600 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0920 -0.0220 0.0920 0.0220 ;
  LAYER v4   ; RECT -0.0800 -0.0290 0.0800 0.0290 ;
  LAYER m5   ; RECT -0.0800 -0.0500 0.0800 0.0500 ;
END VIA4_160X58S_44H_160V

VIA VIA4_70X70_56H_200V
  # v4   size: x=0.0700 y=0.0700
  # m4   size: x=0.0940 y=0.0560   enclosure: x=0.0120 y=-0.0070
  # m5   size: x=0.2000 y=0.1120   enclosure: x=0.0650 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0470 -0.0280 0.0470 0.0280 ;
  LAYER v4   ; RECT -0.0350 -0.0350 0.0350 0.0350 ;
  LAYER m5   ; RECT -0.1000 -0.0560 0.1000 0.0560 ;
END VIA4_70X70_56H_200V

VIA VIA4_44X58S_56H_44V
  # v4   size: x=0.0440 y=0.0580
  # m4   size: x=0.0680 y=0.0560   enclosure: x=0.0120 y=-0.0010
  # m5   size: x=0.0440 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0340 -0.0280 0.0340 0.0280 ;
  LAYER v4   ; RECT -0.0220 -0.0290 0.0220 0.0290 ;
  LAYER m5   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
END VIA4_44X58S_56H_44V

VIA VIA4_56X58S_56H_56V
  # v4   size: x=0.0560 y=0.0580
  # m4   size: x=0.0800 y=0.0560   enclosure: x=0.0120 y=-0.0010
  # m5   size: x=0.0560 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0400 -0.0280 0.0400 0.0280 ;
  LAYER v4   ; RECT -0.0280 -0.0290 0.0280 0.0290 ;
  LAYER m5   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
END VIA4_56X58S_56H_56V

VIA VIA4_76X58S_56H_76V
  # v4   size: x=0.0760 y=0.0580
  # m4   size: x=0.1000 y=0.0560   enclosure: x=0.0120 y=-0.0010
  # m5   size: x=0.0760 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
  LAYER v4   ; RECT -0.0380 -0.0290 0.0380 0.0290 ;
  LAYER m5   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
END VIA4_76X58S_56H_76V

VIA VIA4_90X58S_56H_90V
  # v4   size: x=0.0900 y=0.0580
  # m4   size: x=0.1140 y=0.0560   enclosure: x=0.0120 y=-0.0010
  # m5   size: x=0.0900 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0570 -0.0280 0.0570 0.0280 ;
  LAYER v4   ; RECT -0.0450 -0.0290 0.0450 0.0290 ;
  LAYER m5   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
END VIA4_90X58S_56H_90V

VIA VIA4_108X58S_56H_108V
  # v4   size: x=0.1080 y=0.0580
  # m4   size: x=0.1320 y=0.0560   enclosure: x=0.0120 y=-0.0010
  # m5   size: x=0.1080 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0660 -0.0280 0.0660 0.0280 ;
  LAYER v4   ; RECT -0.0540 -0.0290 0.0540 0.0290 ;
  LAYER m5   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
END VIA4_108X58S_56H_108V

VIA VIA4_160X58S_56H_160V
  # v4   size: x=0.1600 y=0.0580
  # m4   size: x=0.1840 y=0.0560   enclosure: x=0.0120 y=-0.0010
  # m5   size: x=0.1600 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0920 -0.0280 0.0920 0.0280 ;
  LAYER v4   ; RECT -0.0800 -0.0290 0.0800 0.0290 ;
  LAYER m5   ; RECT -0.0800 -0.0500 0.0800 0.0500 ;
END VIA4_160X58S_56H_160V

VIA VIA4_44X58S_76H_44V
  # v4   size: x=0.0440 y=0.0580
  # m4   size: x=0.0680 y=0.0760   enclosure: x=0.0120 y=0.0090
  # m5   size: x=0.0440 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0340 -0.0380 0.0340 0.0380 ;
  LAYER v4   ; RECT -0.0220 -0.0290 0.0220 0.0290 ;
  LAYER m5   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
END VIA4_44X58S_76H_44V

VIA VIA4_56X58S_76H_56V
  # v4   size: x=0.0560 y=0.0580
  # m4   size: x=0.0800 y=0.0760   enclosure: x=0.0120 y=0.0090
  # m5   size: x=0.0560 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0400 -0.0380 0.0400 0.0380 ;
  LAYER v4   ; RECT -0.0280 -0.0290 0.0280 0.0290 ;
  LAYER m5   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
END VIA4_56X58S_76H_56V

VIA VIA4_76X58S_76H_76V
  # v4   size: x=0.0760 y=0.0580
  # m4   size: x=0.1000 y=0.0760   enclosure: x=0.0120 y=0.0090
  # m5   size: x=0.0760 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
  LAYER v4   ; RECT -0.0380 -0.0290 0.0380 0.0290 ;
  LAYER m5   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
END VIA4_76X58S_76H_76V

VIA VIA4_90X58S_76H_90V
  # v4   size: x=0.0900 y=0.0580
  # m4   size: x=0.1140 y=0.0760   enclosure: x=0.0120 y=0.0090
  # m5   size: x=0.0900 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0570 -0.0380 0.0570 0.0380 ;
  LAYER v4   ; RECT -0.0450 -0.0290 0.0450 0.0290 ;
  LAYER m5   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
END VIA4_90X58S_76H_90V

VIA VIA4_108X58S_76H_108V
  # v4   size: x=0.1080 y=0.0580
  # m4   size: x=0.1320 y=0.0760   enclosure: x=0.0120 y=0.0090
  # m5   size: x=0.1080 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0660 -0.0380 0.0660 0.0380 ;
  LAYER v4   ; RECT -0.0540 -0.0290 0.0540 0.0290 ;
  LAYER m5   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
END VIA4_108X58S_76H_108V

VIA VIA4_160X58S_76H_160V
  # v4   size: x=0.1600 y=0.0580
  # m4   size: x=0.1840 y=0.0760   enclosure: x=0.0120 y=0.0090
  # m5   size: x=0.1600 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0920 -0.0380 0.0920 0.0380 ;
  LAYER v4   ; RECT -0.0800 -0.0290 0.0800 0.0290 ;
  LAYER m5   ; RECT -0.0800 -0.0500 0.0800 0.0500 ;
END VIA4_160X58S_76H_160V

VIA VIA4_70X70_76H_200V
  # v4   size: x=0.0700 y=0.0700
  # m4   size: x=0.0940 y=0.0760   enclosure: x=0.0120 y=0.0030
  # m5   size: x=0.2000 y=0.1120   enclosure: x=0.0650 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0470 -0.0380 0.0470 0.0380 ;
  LAYER v4   ; RECT -0.0350 -0.0350 0.0350 0.0350 ;
  LAYER m5   ; RECT -0.1000 -0.0560 0.1000 0.0560 ;
END VIA4_70X70_76H_200V

VIA VIA4_44X58S_90H_44V
  # v4   size: x=0.0440 y=0.0580
  # m4   size: x=0.0680 y=0.0900   enclosure: x=0.0120 y=0.0160
  # m5   size: x=0.0440 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0340 -0.0450 0.0340 0.0450 ;
  LAYER v4   ; RECT -0.0220 -0.0290 0.0220 0.0290 ;
  LAYER m5   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
END VIA4_44X58S_90H_44V

VIA VIA4_56X58S_90H_56V
  # v4   size: x=0.0560 y=0.0580
  # m4   size: x=0.0800 y=0.0900   enclosure: x=0.0120 y=0.0160
  # m5   size: x=0.0560 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0400 -0.0450 0.0400 0.0450 ;
  LAYER v4   ; RECT -0.0280 -0.0290 0.0280 0.0290 ;
  LAYER m5   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
END VIA4_56X58S_90H_56V

VIA VIA4_76X58S_90H_76V
  # v4   size: x=0.0760 y=0.0580
  # m4   size: x=0.1000 y=0.0900   enclosure: x=0.0120 y=0.0160
  # m5   size: x=0.0760 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
  LAYER v4   ; RECT -0.0380 -0.0290 0.0380 0.0290 ;
  LAYER m5   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
END VIA4_76X58S_90H_76V

VIA VIA4_90X58S_90H_90V
  # v4   size: x=0.0900 y=0.0580
  # m4   size: x=0.1140 y=0.0900   enclosure: x=0.0120 y=0.0160
  # m5   size: x=0.0900 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0570 -0.0450 0.0570 0.0450 ;
  LAYER v4   ; RECT -0.0450 -0.0290 0.0450 0.0290 ;
  LAYER m5   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
END VIA4_90X58S_90H_90V

VIA VIA4_108X58S_90H_108V
  # v4   size: x=0.1080 y=0.0580
  # m4   size: x=0.1320 y=0.0900   enclosure: x=0.0120 y=0.0160
  # m5   size: x=0.1080 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0660 -0.0450 0.0660 0.0450 ;
  LAYER v4   ; RECT -0.0540 -0.0290 0.0540 0.0290 ;
  LAYER m5   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
END VIA4_108X58S_90H_108V

VIA VIA4_160X58S_90H_160V
  # v4   size: x=0.1600 y=0.0580
  # m4   size: x=0.1840 y=0.0900   enclosure: x=0.0120 y=0.0160
  # m5   size: x=0.1600 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0920 -0.0450 0.0920 0.0450 ;
  LAYER v4   ; RECT -0.0800 -0.0290 0.0800 0.0290 ;
  LAYER m5   ; RECT -0.0800 -0.0500 0.0800 0.0500 ;
END VIA4_160X58S_90H_160V

VIA VIA4_70X70_90H_200V
  # v4   size: x=0.0700 y=0.0700
  # m4   size: x=0.0940 y=0.0900   enclosure: x=0.0120 y=0.0100
  # m5   size: x=0.2000 y=0.1120   enclosure: x=0.0650 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0470 -0.0450 0.0470 0.0450 ;
  LAYER v4   ; RECT -0.0350 -0.0350 0.0350 0.0350 ;
  LAYER m5   ; RECT -0.1000 -0.0560 0.1000 0.0560 ;
END VIA4_70X70_90H_200V

VIA VIA4_44X58S_108H_44V
  # v4   size: x=0.0440 y=0.0580
  # m4   size: x=0.0680 y=0.1080   enclosure: x=0.0120 y=0.0250
  # m5   size: x=0.0440 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0340 -0.0540 0.0340 0.0540 ;
  LAYER v4   ; RECT -0.0220 -0.0290 0.0220 0.0290 ;
  LAYER m5   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
END VIA4_44X58S_108H_44V

VIA VIA4_56X58S_108H_56V
  # v4   size: x=0.0560 y=0.0580
  # m4   size: x=0.0800 y=0.1080   enclosure: x=0.0120 y=0.0250
  # m5   size: x=0.0560 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0400 -0.0540 0.0400 0.0540 ;
  LAYER v4   ; RECT -0.0280 -0.0290 0.0280 0.0290 ;
  LAYER m5   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
END VIA4_56X58S_108H_56V

VIA VIA4_76X58S_108H_76V
  # v4   size: x=0.0760 y=0.0580
  # m4   size: x=0.1000 y=0.1080   enclosure: x=0.0120 y=0.0250
  # m5   size: x=0.0760 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
  LAYER v4   ; RECT -0.0380 -0.0290 0.0380 0.0290 ;
  LAYER m5   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
END VIA4_76X58S_108H_76V

VIA VIA4_90X58S_108H_90V
  # v4   size: x=0.0900 y=0.0580
  # m4   size: x=0.1140 y=0.1080   enclosure: x=0.0120 y=0.0250
  # m5   size: x=0.0900 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0570 -0.0540 0.0570 0.0540 ;
  LAYER v4   ; RECT -0.0450 -0.0290 0.0450 0.0290 ;
  LAYER m5   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
END VIA4_90X58S_108H_90V

VIA VIA4_108X58S_108H_108V
  # v4   size: x=0.1080 y=0.0580
  # m4   size: x=0.1320 y=0.1080   enclosure: x=0.0120 y=0.0250
  # m5   size: x=0.1080 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0660 -0.0540 0.0660 0.0540 ;
  LAYER v4   ; RECT -0.0540 -0.0290 0.0540 0.0290 ;
  LAYER m5   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
END VIA4_108X58S_108H_108V

VIA VIA4_160X58S_108H_160V
  # v4   size: x=0.1600 y=0.0580
  # m4   size: x=0.1840 y=0.1080   enclosure: x=0.0120 y=0.0250
  # m5   size: x=0.1600 y=0.1000   enclosure: x=0.0000 y=0.0210
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0920 -0.0540 0.0920 0.0540 ;
  LAYER v4   ; RECT -0.0800 -0.0290 0.0800 0.0290 ;
  LAYER m5   ; RECT -0.0800 -0.0500 0.0800 0.0500 ;
END VIA4_160X58S_108H_160V

VIA VIA4_90X90_108H_200V
  # v4   size: x=0.0900 y=0.0900
  # m4   size: x=0.1140 y=0.1080   enclosure: x=0.0120 y=0.0090
  # m5   size: x=0.2000 y=0.1700   enclosure: x=0.0550 y=0.0400
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.0570 -0.0540 0.0570 0.0540 ;
  LAYER v4   ; RECT -0.0450 -0.0450 0.0450 0.0450 ;
  LAYER m5   ; RECT -0.1000 -0.0850 0.1000 0.0850 ;
END VIA4_90X90_108H_200V

VIA VIA5_58SX44_44V_44H
  # v5   size: x=0.0580 y=0.0440
  # m5   size: x=0.0440 y=0.0680   enclosure: x=-0.0070 y=0.0120
  # m6   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0220 -0.0340 0.0220 0.0340 ;
  LAYER v5   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m6   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA5_58SX44_44V_44H

VIA VIA5_58SX56_44V_56H
  # v5   size: x=0.0580 y=0.0560
  # m5   size: x=0.0440 y=0.0800   enclosure: x=-0.0070 y=0.0120
  # m6   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0220 -0.0400 0.0220 0.0400 ;
  LAYER v5   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m6   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA5_58SX56_44V_56H

VIA VIA5_58SX76_44V_76H
  # v5   size: x=0.0580 y=0.0760
  # m5   size: x=0.0440 y=0.1000   enclosure: x=-0.0070 y=0.0120
  # m6   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0220 -0.0500 0.0220 0.0500 ;
  LAYER v5   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m6   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA5_58SX76_44V_76H

VIA VIA5_58SX90_44V_90H
  # v5   size: x=0.0580 y=0.0900
  # m5   size: x=0.0440 y=0.1140   enclosure: x=-0.0070 y=0.0120
  # m6   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0220 -0.0570 0.0220 0.0570 ;
  LAYER v5   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m6   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA5_58SX90_44V_90H

VIA VIA5_58SX108_44V_108H
  # v5   size: x=0.0580 y=0.1080
  # m5   size: x=0.0440 y=0.1320   enclosure: x=-0.0070 y=0.0120
  # m6   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0220 -0.0660 0.0220 0.0660 ;
  LAYER v5   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m6   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA5_58SX108_44V_108H

VIA VIA5_58SX160_44V_160H
  # v5   size: x=0.0580 y=0.1600
  # m5   size: x=0.0440 y=0.1840   enclosure: x=-0.0070 y=0.0120
  # m6   size: x=0.1000 y=0.1600   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0220 -0.0920 0.0220 0.0920 ;
  LAYER v5   ; RECT -0.0290 -0.0800 0.0290 0.0800 ;
  LAYER m6   ; RECT -0.0500 -0.0800 0.0500 0.0800 ;
END VIA5_58SX160_44V_160H

VIA VIA5_70X70_56V_200H
  # v5   size: x=0.0700 y=0.0700
  # m5   size: x=0.0560 y=0.0940   enclosure: x=-0.0070 y=0.0120
  # m6   size: x=0.1120 y=0.2000   enclosure: x=0.0210 y=0.0650
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0280 -0.0470 0.0280 0.0470 ;
  LAYER v5   ; RECT -0.0350 -0.0350 0.0350 0.0350 ;
  LAYER m6   ; RECT -0.0560 -0.1000 0.0560 0.1000 ;
END VIA5_70X70_56V_200H

VIA VIA5_70X70_56V_400H
  # v5   size: x=0.0700 y=0.0700
  # m5   size: x=0.0560 y=0.0940   enclosure: x=-0.0070 y=0.0120
  # m6   size: x=0.1120 y=0.4000   enclosure: x=0.0210 y=0.1650
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0280 -0.0470 0.0280 0.0470 ;
  LAYER v5   ; RECT -0.0350 -0.0350 0.0350 0.0350 ;
  LAYER m6   ; RECT -0.0560 -0.2000 0.0560 0.2000 ;
END VIA5_70X70_56V_400H

VIA VIA5_58SX44_56V_44H
  # v5   size: x=0.0580 y=0.0440
  # m5   size: x=0.0560 y=0.0680   enclosure: x=-0.0010 y=0.0120
  # m6   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0280 -0.0340 0.0280 0.0340 ;
  LAYER v5   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m6   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA5_58SX44_56V_44H

VIA VIA5_58SX56_56V_56H
  # v5   size: x=0.0580 y=0.0560
  # m5   size: x=0.0560 y=0.0800   enclosure: x=-0.0010 y=0.0120
  # m6   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0280 -0.0400 0.0280 0.0400 ;
  LAYER v5   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m6   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA5_58SX56_56V_56H

VIA VIA5_58SX76_56V_76H
  # v5   size: x=0.0580 y=0.0760
  # m5   size: x=0.0560 y=0.1000   enclosure: x=-0.0010 y=0.0120
  # m6   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0280 -0.0500 0.0280 0.0500 ;
  LAYER v5   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m6   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA5_58SX76_56V_76H

VIA VIA5_58SX90_56V_90H
  # v5   size: x=0.0580 y=0.0900
  # m5   size: x=0.0560 y=0.1140   enclosure: x=-0.0010 y=0.0120
  # m6   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0280 -0.0570 0.0280 0.0570 ;
  LAYER v5   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m6   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA5_58SX90_56V_90H

VIA VIA5_58SX108_56V_108H
  # v5   size: x=0.0580 y=0.1080
  # m5   size: x=0.0560 y=0.1320   enclosure: x=-0.0010 y=0.0120
  # m6   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0280 -0.0660 0.0280 0.0660 ;
  LAYER v5   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m6   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA5_58SX108_56V_108H

VIA VIA5_58SX160_56V_160H
  # v5   size: x=0.0580 y=0.1600
  # m5   size: x=0.0560 y=0.1840   enclosure: x=-0.0010 y=0.0120
  # m6   size: x=0.1000 y=0.1600   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0280 -0.0920 0.0280 0.0920 ;
  LAYER v5   ; RECT -0.0290 -0.0800 0.0290 0.0800 ;
  LAYER m6   ; RECT -0.0500 -0.0800 0.0500 0.0800 ;
END VIA5_58SX160_56V_160H

VIA VIA5_58SX44_76V_44H
  # v5   size: x=0.0580 y=0.0440
  # m5   size: x=0.0760 y=0.0680   enclosure: x=0.0090 y=0.0120
  # m6   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0380 -0.0340 0.0380 0.0340 ;
  LAYER v5   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m6   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA5_58SX44_76V_44H

VIA VIA5_58SX56_76V_56H
  # v5   size: x=0.0580 y=0.0560
  # m5   size: x=0.0760 y=0.0800   enclosure: x=0.0090 y=0.0120
  # m6   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0380 -0.0400 0.0380 0.0400 ;
  LAYER v5   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m6   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA5_58SX56_76V_56H

VIA VIA5_58SX76_76V_76H
  # v5   size: x=0.0580 y=0.0760
  # m5   size: x=0.0760 y=0.1000   enclosure: x=0.0090 y=0.0120
  # m6   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0380 -0.0500 0.0380 0.0500 ;
  LAYER v5   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m6   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA5_58SX76_76V_76H

VIA VIA5_58SX90_76V_90H
  # v5   size: x=0.0580 y=0.0900
  # m5   size: x=0.0760 y=0.1140   enclosure: x=0.0090 y=0.0120
  # m6   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0380 -0.0570 0.0380 0.0570 ;
  LAYER v5   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m6   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA5_58SX90_76V_90H

VIA VIA5_58SX108_76V_108H
  # v5   size: x=0.0580 y=0.1080
  # m5   size: x=0.0760 y=0.1320   enclosure: x=0.0090 y=0.0120
  # m6   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0380 -0.0660 0.0380 0.0660 ;
  LAYER v5   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m6   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA5_58SX108_76V_108H

VIA VIA5_58SX160_76V_160H
  # v5   size: x=0.0580 y=0.1600
  # m5   size: x=0.0760 y=0.1840   enclosure: x=0.0090 y=0.0120
  # m6   size: x=0.1000 y=0.1600   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0380 -0.0920 0.0380 0.0920 ;
  LAYER v5   ; RECT -0.0290 -0.0800 0.0290 0.0800 ;
  LAYER m6   ; RECT -0.0500 -0.0800 0.0500 0.0800 ;
END VIA5_58SX160_76V_160H

VIA VIA5_70X70_76V_200H
  # v5   size: x=0.0700 y=0.0700
  # m5   size: x=0.0760 y=0.0940   enclosure: x=0.0030 y=0.0120
  # m6   size: x=0.1120 y=0.2000   enclosure: x=0.0210 y=0.0650
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0380 -0.0470 0.0380 0.0470 ;
  LAYER v5   ; RECT -0.0350 -0.0350 0.0350 0.0350 ;
  LAYER m6   ; RECT -0.0560 -0.1000 0.0560 0.1000 ;
END VIA5_70X70_76V_200H

VIA VIA5_70X70_76V_400H
  # v5   size: x=0.0700 y=0.0700
  # m5   size: x=0.0760 y=0.0940   enclosure: x=0.0030 y=0.0120
  # m6   size: x=0.1120 y=0.4000   enclosure: x=0.0210 y=0.1650
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0380 -0.0470 0.0380 0.0470 ;
  LAYER v5   ; RECT -0.0350 -0.0350 0.0350 0.0350 ;
  LAYER m6   ; RECT -0.0560 -0.2000 0.0560 0.2000 ;
END VIA5_70X70_76V_400H

VIA VIA5_58SX44_90V_44H
  # v5   size: x=0.0580 y=0.0440
  # m5   size: x=0.0900 y=0.0680   enclosure: x=0.0160 y=0.0120
  # m6   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0450 -0.0340 0.0450 0.0340 ;
  LAYER v5   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m6   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA5_58SX44_90V_44H

VIA VIA5_58SX56_90V_56H
  # v5   size: x=0.0580 y=0.0560
  # m5   size: x=0.0900 y=0.0800   enclosure: x=0.0160 y=0.0120
  # m6   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0450 -0.0400 0.0450 0.0400 ;
  LAYER v5   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m6   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA5_58SX56_90V_56H

VIA VIA5_58SX76_90V_76H
  # v5   size: x=0.0580 y=0.0760
  # m5   size: x=0.0900 y=0.1000   enclosure: x=0.0160 y=0.0120
  # m6   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0450 -0.0500 0.0450 0.0500 ;
  LAYER v5   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m6   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA5_58SX76_90V_76H

VIA VIA5_58SX90_90V_90H
  # v5   size: x=0.0580 y=0.0900
  # m5   size: x=0.0900 y=0.1140   enclosure: x=0.0160 y=0.0120
  # m6   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0450 -0.0570 0.0450 0.0570 ;
  LAYER v5   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m6   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA5_58SX90_90V_90H

VIA VIA5_58SX108_90V_108H
  # v5   size: x=0.0580 y=0.1080
  # m5   size: x=0.0900 y=0.1320   enclosure: x=0.0160 y=0.0120
  # m6   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0450 -0.0660 0.0450 0.0660 ;
  LAYER v5   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m6   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA5_58SX108_90V_108H

VIA VIA5_58SX160_90V_160H
  # v5   size: x=0.0580 y=0.1600
  # m5   size: x=0.0900 y=0.1840   enclosure: x=0.0160 y=0.0120
  # m6   size: x=0.1000 y=0.1600   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0450 -0.0920 0.0450 0.0920 ;
  LAYER v5   ; RECT -0.0290 -0.0800 0.0290 0.0800 ;
  LAYER m6   ; RECT -0.0500 -0.0800 0.0500 0.0800 ;
END VIA5_58SX160_90V_160H

VIA VIA5_70X70_90V_200H
  # v5   size: x=0.0700 y=0.0700
  # m5   size: x=0.0900 y=0.0940   enclosure: x=0.0100 y=0.0120
  # m6   size: x=0.1120 y=0.2000   enclosure: x=0.0210 y=0.0650
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0450 -0.0470 0.0450 0.0470 ;
  LAYER v5   ; RECT -0.0350 -0.0350 0.0350 0.0350 ;
  LAYER m6   ; RECT -0.0560 -0.1000 0.0560 0.1000 ;
END VIA5_70X70_90V_200H

VIA VIA5_70X70_90V_400H
  # v5   size: x=0.0700 y=0.0700
  # m5   size: x=0.0900 y=0.0940   enclosure: x=0.0100 y=0.0120
  # m6   size: x=0.1120 y=0.4000   enclosure: x=0.0210 y=0.1650
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0450 -0.0470 0.0450 0.0470 ;
  LAYER v5   ; RECT -0.0350 -0.0350 0.0350 0.0350 ;
  LAYER m6   ; RECT -0.0560 -0.2000 0.0560 0.2000 ;
END VIA5_70X70_90V_400H

VIA VIA5_58SX44_108V_44H
  # v5   size: x=0.0580 y=0.0440
  # m5   size: x=0.1080 y=0.0680   enclosure: x=0.0250 y=0.0120
  # m6   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0540 -0.0340 0.0540 0.0340 ;
  LAYER v5   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m6   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA5_58SX44_108V_44H

VIA VIA5_58SX56_108V_56H
  # v5   size: x=0.0580 y=0.0560
  # m5   size: x=0.1080 y=0.0800   enclosure: x=0.0250 y=0.0120
  # m6   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0540 -0.0400 0.0540 0.0400 ;
  LAYER v5   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m6   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA5_58SX56_108V_56H

VIA VIA5_58SX76_108V_76H
  # v5   size: x=0.0580 y=0.0760
  # m5   size: x=0.1080 y=0.1000   enclosure: x=0.0250 y=0.0120
  # m6   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0540 -0.0500 0.0540 0.0500 ;
  LAYER v5   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m6   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA5_58SX76_108V_76H

VIA VIA5_58SX90_108V_90H
  # v5   size: x=0.0580 y=0.0900
  # m5   size: x=0.1080 y=0.1140   enclosure: x=0.0250 y=0.0120
  # m6   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0540 -0.0570 0.0540 0.0570 ;
  LAYER v5   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m6   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA5_58SX90_108V_90H

VIA VIA5_58SX108_108V_108H
  # v5   size: x=0.0580 y=0.1080
  # m5   size: x=0.1080 y=0.1320   enclosure: x=0.0250 y=0.0120
  # m6   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0540 -0.0660 0.0540 0.0660 ;
  LAYER v5   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m6   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA5_58SX108_108V_108H

VIA VIA5_58SX160_108V_160H
  # v5   size: x=0.0580 y=0.1600
  # m5   size: x=0.1080 y=0.1840   enclosure: x=0.0250 y=0.0120
  # m6   size: x=0.1000 y=0.1600   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0540 -0.0920 0.0540 0.0920 ;
  LAYER v5   ; RECT -0.0290 -0.0800 0.0290 0.0800 ;
  LAYER m6   ; RECT -0.0500 -0.0800 0.0500 0.0800 ;
END VIA5_58SX160_108V_160H

VIA VIA5_90X90_108V_200H
  # v5   size: x=0.0900 y=0.0900
  # m5   size: x=0.1080 y=0.1140   enclosure: x=0.0090 y=0.0120
  # m6   size: x=0.1700 y=0.2000   enclosure: x=0.0400 y=0.0550
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0540 -0.0570 0.0540 0.0570 ;
  LAYER v5   ; RECT -0.0450 -0.0450 0.0450 0.0450 ;
  LAYER m6   ; RECT -0.0850 -0.1000 0.0850 0.1000 ;
END VIA5_90X90_108V_200H

VIA VIA5_90X90_108V_400H
  # v5   size: x=0.0900 y=0.0900
  # m5   size: x=0.1080 y=0.1140   enclosure: x=0.0090 y=0.0120
  # m6   size: x=0.1700 y=0.4000   enclosure: x=0.0400 y=0.1550
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0540 -0.0570 0.0540 0.0570 ;
  LAYER v5   ; RECT -0.0450 -0.0450 0.0450 0.0450 ;
  LAYER m6   ; RECT -0.0850 -0.2000 0.0850 0.2000 ;
END VIA5_90X90_108V_400H

VIA VIA5_58SX44_160V_44H
  # v5   size: x=0.0580 y=0.0440
  # m5   size: x=0.1600 y=0.0680   enclosure: x=0.0510 y=0.0120
  # m6   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0800 -0.0340 0.0800 0.0340 ;
  LAYER v5   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m6   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA5_58SX44_160V_44H

VIA VIA5_58SX56_160V_56H
  # v5   size: x=0.0580 y=0.0560
  # m5   size: x=0.1600 y=0.0800   enclosure: x=0.0510 y=0.0120
  # m6   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0800 -0.0400 0.0800 0.0400 ;
  LAYER v5   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m6   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA5_58SX56_160V_56H

VIA VIA5_58SX76_160V_76H
  # v5   size: x=0.0580 y=0.0760
  # m5   size: x=0.1600 y=0.1000   enclosure: x=0.0510 y=0.0120
  # m6   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0800 -0.0500 0.0800 0.0500 ;
  LAYER v5   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m6   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA5_58SX76_160V_76H

VIA VIA5_58SX90_160V_90H
  # v5   size: x=0.0580 y=0.0900
  # m5   size: x=0.1600 y=0.1140   enclosure: x=0.0510 y=0.0120
  # m6   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0800 -0.0570 0.0800 0.0570 ;
  LAYER v5   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m6   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA5_58SX90_160V_90H

VIA VIA5_58SX108_160V_108H
  # v5   size: x=0.0580 y=0.1080
  # m5   size: x=0.1600 y=0.1320   enclosure: x=0.0510 y=0.0120
  # m6   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0800 -0.0660 0.0800 0.0660 ;
  LAYER v5   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m6   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA5_58SX108_160V_108H

VIA VIA5_58SX160_160V_160H
  # v5   size: x=0.0580 y=0.1600
  # m5   size: x=0.1600 y=0.1840   enclosure: x=0.0510 y=0.0120
  # m6   size: x=0.1000 y=0.1600   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0800 -0.0920 0.0800 0.0920 ;
  LAYER v5   ; RECT -0.0290 -0.0800 0.0290 0.0800 ;
  LAYER m6   ; RECT -0.0500 -0.0800 0.0500 0.0800 ;
END VIA5_58SX160_160V_160H

VIA VIA5_90X90_160V_200H
  # v5   size: x=0.0900 y=0.0900
  # m5   size: x=0.1600 y=0.1140   enclosure: x=0.0350 y=0.0120
  # m6   size: x=0.1700 y=0.2000   enclosure: x=0.0400 y=0.0550
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0800 -0.0570 0.0800 0.0570 ;
  LAYER v5   ; RECT -0.0450 -0.0450 0.0450 0.0450 ;
  LAYER m6   ; RECT -0.0850 -0.1000 0.0850 0.1000 ;
END VIA5_90X90_160V_200H

VIA VIA5_90X90_160V_400H
  # v5   size: x=0.0900 y=0.0900
  # m5   size: x=0.1600 y=0.1140   enclosure: x=0.0350 y=0.0120
  # m6   size: x=0.1700 y=0.4000   enclosure: x=0.0400 y=0.1550
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.0800 -0.0570 0.0800 0.0570 ;
  LAYER v5   ; RECT -0.0450 -0.0450 0.0450 0.0450 ;
  LAYER m6   ; RECT -0.0850 -0.2000 0.0850 0.2000 ;
END VIA5_90X90_160V_400H

VIA VIA5_58SX44_200V_44H
  # v5   size: x=0.0580 y=0.0440
  # m5   size: x=0.2000 y=0.0680   enclosure: x=0.0710 y=0.0120
  # m6   size: x=0.1000 y=0.0440   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.1000 -0.0340 0.1000 0.0340 ;
  LAYER v5   ; RECT -0.0290 -0.0220 0.0290 0.0220 ;
  LAYER m6   ; RECT -0.0500 -0.0220 0.0500 0.0220 ;
END VIA5_58SX44_200V_44H

VIA VIA5_58SX56_200V_56H
  # v5   size: x=0.0580 y=0.0560
  # m5   size: x=0.2000 y=0.0800   enclosure: x=0.0710 y=0.0120
  # m6   size: x=0.1000 y=0.0560   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.1000 -0.0400 0.1000 0.0400 ;
  LAYER v5   ; RECT -0.0290 -0.0280 0.0290 0.0280 ;
  LAYER m6   ; RECT -0.0500 -0.0280 0.0500 0.0280 ;
END VIA5_58SX56_200V_56H

VIA VIA5_58SX76_200V_76H
  # v5   size: x=0.0580 y=0.0760
  # m5   size: x=0.2000 y=0.1000   enclosure: x=0.0710 y=0.0120
  # m6   size: x=0.1000 y=0.0760   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.1000 -0.0500 0.1000 0.0500 ;
  LAYER v5   ; RECT -0.0290 -0.0380 0.0290 0.0380 ;
  LAYER m6   ; RECT -0.0500 -0.0380 0.0500 0.0380 ;
END VIA5_58SX76_200V_76H

VIA VIA5_58SX90_200V_90H
  # v5   size: x=0.0580 y=0.0900
  # m5   size: x=0.2000 y=0.1140   enclosure: x=0.0710 y=0.0120
  # m6   size: x=0.1000 y=0.0900   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.1000 -0.0570 0.1000 0.0570 ;
  LAYER v5   ; RECT -0.0290 -0.0450 0.0290 0.0450 ;
  LAYER m6   ; RECT -0.0500 -0.0450 0.0500 0.0450 ;
END VIA5_58SX90_200V_90H

VIA VIA5_58SX108_200V_108H
  # v5   size: x=0.0580 y=0.1080
  # m5   size: x=0.2000 y=0.1320   enclosure: x=0.0710 y=0.0120
  # m6   size: x=0.1000 y=0.1080   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.1000 -0.0660 0.1000 0.0660 ;
  LAYER v5   ; RECT -0.0290 -0.0540 0.0290 0.0540 ;
  LAYER m6   ; RECT -0.0500 -0.0540 0.0500 0.0540 ;
END VIA5_58SX108_200V_108H

VIA VIA5_58SX160_200V_160H
  # v5   size: x=0.0580 y=0.1600
  # m5   size: x=0.2000 y=0.1840   enclosure: x=0.0710 y=0.0120
  # m6   size: x=0.1000 y=0.1600   enclosure: x=0.0210 y=0.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.1000 -0.0920 0.1000 0.0920 ;
  LAYER v5   ; RECT -0.0290 -0.0800 0.0290 0.0800 ;
  LAYER m6   ; RECT -0.0500 -0.0800 0.0500 0.0800 ;
END VIA5_58SX160_200V_160H

VIA VIA5_90X90_200V_200H
  # v5   size: x=0.0900 y=0.0900
  # m5   size: x=0.2000 y=0.1140   enclosure: x=0.0550 y=0.0120
  # m6   size: x=0.1700 y=0.2000   enclosure: x=0.0400 y=0.0550
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.1000 -0.0570 0.1000 0.0570 ;
  LAYER v5   ; RECT -0.0450 -0.0450 0.0450 0.0450 ;
  LAYER m6   ; RECT -0.0850 -0.1000 0.0850 0.1000 ;
END VIA5_90X90_200V_200H

VIA VIA5_90X90_200V_400H
  # v5   size: x=0.0900 y=0.0900
  # m5   size: x=0.2000 y=0.1140   enclosure: x=0.0550 y=0.0120
  # m6   size: x=0.1700 y=0.4000   enclosure: x=0.0400 y=0.1550
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.1000 -0.0570 0.1000 0.0570 ;
  LAYER v5   ; RECT -0.0450 -0.0450 0.0450 0.0450 ;
  LAYER m6   ; RECT -0.0850 -0.2000 0.0850 0.2000 ;
END VIA5_90X90_200V_400H

VIA VIA6_200X120U_160H_180V
  # v6   size: x=0.2000 y=0.1200
  # m6   size: x=0.3200 y=0.1600   enclosure: x=0.0600 y=0.0200
  # m7   size: x=0.1800 y=0.2400   enclosure: x=-0.0100 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.1600 -0.0800 0.1600 0.0800 ;
  LAYER v6   ; RECT -0.1000 -0.0600 0.1000 0.0600 ;
  LAYER m7   ; RECT -0.0900 -0.1200 0.0900 0.1200 ;
END VIA6_200X120U_160H_180V

VIA VIA6_120X200_400H_180V
  # v6   size: x=0.1200 y=0.2000
  # m6   size: x=0.2400 y=0.4000   enclosure: x=0.0600 y=0.1000
  # m7   size: x=0.1800 y=0.3200   enclosure: x=0.0300 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.1200 -0.2000 0.1200 0.2000 ;
  LAYER v6   ; RECT -0.0600 -0.1000 0.0600 0.1000 ;
  LAYER m7   ; RECT -0.0900 -0.1600 0.0900 0.1600 ;
END VIA6_120X200_400H_180V

VIA VIA6_200X120_160H_260V
  # v6   size: x=0.2000 y=0.1200
  # m6   size: x=0.3200 y=0.1600   enclosure: x=0.0600 y=0.0200
  # m7   size: x=0.2600 y=0.2400   enclosure: x=0.0300 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.1600 -0.0800 0.1600 0.0800 ;
  LAYER v6   ; RECT -0.1000 -0.0600 0.1000 0.0600 ;
  LAYER m7   ; RECT -0.1300 -0.1200 0.1300 0.1200 ;
END VIA6_200X120_160H_260V

VIA VIA6_400X120_160H_460V
  # v6   size: x=0.4000 y=0.1200
  # m6   size: x=0.5200 y=0.1600   enclosure: x=0.0600 y=0.0200
  # m7   size: x=0.4600 y=0.2400   enclosure: x=0.0300 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.2600 -0.0800 0.2600 0.0800 ;
  LAYER v6   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER m7   ; RECT -0.2300 -0.1200 0.2300 0.1200 ;
END VIA6_400X120_160H_460V

VIA VIA6_200X120U_200H_180V
  # v6   size: x=0.2000 y=0.1200
  # m6   size: x=0.3200 y=0.2000   enclosure: x=0.0600 y=0.0400
  # m7   size: x=0.1800 y=0.2400   enclosure: x=-0.0100 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.1600 -0.1000 0.1600 0.1000 ;
  LAYER v6   ; RECT -0.1000 -0.0600 0.1000 0.0600 ;
  LAYER m7   ; RECT -0.0900 -0.1200 0.0900 0.1200 ;
END VIA6_200X120U_200H_180V

VIA VIA6_200X120_200H_260V
  # v6   size: x=0.2000 y=0.1200
  # m6   size: x=0.3200 y=0.2000   enclosure: x=0.0600 y=0.0400
  # m7   size: x=0.2600 y=0.2400   enclosure: x=0.0300 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.1600 -0.1000 0.1600 0.1000 ;
  LAYER v6   ; RECT -0.1000 -0.0600 0.1000 0.0600 ;
  LAYER m7   ; RECT -0.1300 -0.1200 0.1300 0.1200 ;
END VIA6_200X120_200H_260V

VIA VIA6_400X120_200H_460V
  # v6   size: x=0.4000 y=0.1200
  # m6   size: x=0.5200 y=0.2000   enclosure: x=0.0600 y=0.0400
  # m7   size: x=0.4600 y=0.2400   enclosure: x=0.0300 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.2600 -0.1000 0.2600 0.1000 ;
  LAYER v6   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER m7   ; RECT -0.2300 -0.1200 0.2300 0.1200 ;
END VIA6_400X120_200H_460V

VIA VIA6_400X120_400H_460V
  # v6   size: x=0.4000 y=0.1200
  # m6   size: x=0.5200 y=0.4000   enclosure: x=0.0600 y=0.1400
  # m7   size: x=0.4600 y=0.2400   enclosure: x=0.0300 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.2600 -0.2000 0.2600 0.2000 ;
  LAYER v6   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER m7   ; RECT -0.2300 -0.1200 0.2300 0.1200 ;
END VIA6_400X120_400H_460V

VIA VIA7_120UX200_180V_180H
  # v7   size: x=0.1200 y=0.2000
  # m7   size: x=0.1800 y=0.3200   enclosure: x=0.0300 y=0.0600
  # m8   size: x=0.2400 y=0.1800   enclosure: x=0.0600 y=-0.0100
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.0900 -0.1600 0.0900 0.1600 ;
  LAYER v7   ; RECT -0.0600 -0.1000 0.0600 0.1000 ;
  LAYER m8   ; RECT -0.1200 -0.0900 0.1200 0.0900 ;
END VIA7_120UX200_180V_180H

VIA VIA7_200X120_240V_180H
  # v7   size: x=0.2000 y=0.1200
  # m7   size: x=0.2400 y=0.2400   enclosure: x=0.0200 y=0.0600
  # m8   size: x=0.3200 y=0.1800   enclosure: x=0.0600 y=0.0300
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.1200 -0.1200 0.1200 0.1200 ;
  LAYER v7   ; RECT -0.1000 -0.0600 0.1000 0.0600 ;
  LAYER m8   ; RECT -0.1600 -0.0900 0.1600 0.0900 ;
END VIA7_200X120_240V_180H

VIA VIA7_120X200_180V_260H
  # v7   size: x=0.1200 y=0.2000
  # m7   size: x=0.1800 y=0.3200   enclosure: x=0.0300 y=0.0600
  # m8   size: x=0.2400 y=0.2600   enclosure: x=0.0600 y=0.0300
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.0900 -0.1600 0.0900 0.1600 ;
  LAYER v7   ; RECT -0.0600 -0.1000 0.0600 0.1000 ;
  LAYER m8   ; RECT -0.1200 -0.1300 0.1200 0.1300 ;
END VIA7_120X200_180V_260H

VIA VIA7_120X400_180V_460H
  # v7   size: x=0.1200 y=0.4000
  # m7   size: x=0.1800 y=0.5200   enclosure: x=0.0300 y=0.0600
  # m8   size: x=0.2400 y=0.4600   enclosure: x=0.0600 y=0.0300
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.0900 -0.2600 0.0900 0.2600 ;
  LAYER v7   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER m8   ; RECT -0.1200 -0.2300 0.1200 0.2300 ;
END VIA7_120X400_180V_460H

VIA VIA7_400X120_440V_180H
  # v7   size: x=0.4000 y=0.1200
  # m7   size: x=0.4400 y=0.2400   enclosure: x=0.0200 y=0.0600
  # m8   size: x=0.5200 y=0.1800   enclosure: x=0.0600 y=0.0300
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.2200 -0.1200 0.2200 0.1200 ;
  LAYER v7   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER m8   ; RECT -0.2600 -0.0900 0.2600 0.0900 ;
END VIA7_400X120_440V_180H

VIA via7_120x400_600V_460H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3000 -0.2300 0.3000 0.2300 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3000 -0.2300 0.3000 0.2300 ;
END via7_120x400_600V_460H_ARRAY_2x1

VIA via7_120x400_600V_500H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3000 -0.2500 0.3000 0.2500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3000 -0.2500 0.3000 0.2500 ;
END via7_120x400_600V_500H_ARRAY_2x1

VIA via7_120x400_600V_600H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3000 -0.3000 0.3000 0.3000 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3000 -0.3000 0.3000 0.3000 ;
END via7_120x400_600V_600H_ARRAY_2x1

VIA via7_120x400_600V_700H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3000 -0.3500 0.3000 0.3500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3000 -0.3500 0.3000 0.3500 ;
END via7_120x400_600V_700H_ARRAY_2x1

VIA via7_120x400_600V_800H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3000 -0.4000 0.3000 0.4000 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3000 -0.4000 0.3000 0.4000 ;
END via7_120x400_600V_800H_ARRAY_2x1

VIA via7_120x400_600V_900H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3000 -0.4500 0.3000 0.4500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3000 -0.4500 0.3000 0.4500 ;
END via7_120x400_600V_900H_ARRAY_2x1

VIA via7_120x400_700V_460H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3500 -0.2300 0.3500 0.2300 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3500 -0.2300 0.3500 0.2300 ;
END via7_120x400_700V_460H_ARRAY_2x1

VIA via7_120x400_700V_500H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3500 -0.2500 0.3500 0.2500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3500 -0.2500 0.3500 0.2500 ;
END via7_120x400_700V_500H_ARRAY_2x1

VIA via7_120x400_700V_600H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3500 -0.3000 0.3500 0.3000 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3500 -0.3000 0.3500 0.3000 ;
END via7_120x400_700V_600H_ARRAY_2x1

VIA via7_120x400_700V_700H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3500 -0.3500 0.3500 0.3500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3500 -0.3500 0.3500 0.3500 ;
END via7_120x400_700V_700H_ARRAY_2x1

VIA via7_120x400_700V_800H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3500 -0.4000 0.3500 0.4000 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3500 -0.4000 0.3500 0.4000 ;
END via7_120x400_700V_800H_ARRAY_2x1

VIA via7_120x400_700V_900H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.3500 -0.4500 0.3500 0.4500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.3500 -0.4500 0.3500 0.4500 ;
END via7_120x400_700V_900H_ARRAY_2x1

VIA via7_120x400_800V_460H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4000 -0.2300 0.4000 0.2300 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4000 -0.2300 0.4000 0.2300 ;
END via7_120x400_800V_460H_ARRAY_2x1

VIA via7_120x400_800V_500H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4000 -0.2500 0.4000 0.2500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4000 -0.2500 0.4000 0.2500 ;
END via7_120x400_800V_500H_ARRAY_2x1

VIA via7_120x400_800V_600H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4000 -0.3000 0.4000 0.3000 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4000 -0.3000 0.4000 0.3000 ;
END via7_120x400_800V_600H_ARRAY_2x1

VIA via7_120x400_800V_700H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4000 -0.3500 0.4000 0.3500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4000 -0.3500 0.4000 0.3500 ;
END via7_120x400_800V_700H_ARRAY_2x1

VIA via7_120x400_800V_800H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4000 -0.4000 0.4000 0.4000 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4000 -0.4000 0.4000 0.4000 ;
END via7_120x400_800V_800H_ARRAY_2x1

VIA via7_120x400_800V_900H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4000 -0.4500 0.4000 0.4500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4000 -0.4500 0.4000 0.4500 ;
END via7_120x400_800V_900H_ARRAY_2x1

VIA via7_120x400_900V_460H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4500 -0.2300 0.4500 0.2300 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4500 -0.2300 0.4500 0.2300 ;
END via7_120x400_900V_460H_ARRAY_2x1

VIA via7_120x400_900V_500H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4500 -0.2500 0.4500 0.2500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4500 -0.2500 0.4500 0.2500 ;
END via7_120x400_900V_500H_ARRAY_2x1

VIA via7_120x400_900V_600H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4500 -0.3000 0.4500 0.3000 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4500 -0.3000 0.4500 0.3000 ;
END via7_120x400_900V_600H_ARRAY_2x1

VIA via7_120x400_900V_700H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4500 -0.3500 0.4500 0.3500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4500 -0.3500 0.4500 0.3500 ;
END via7_120x400_900V_700H_ARRAY_2x1

VIA via7_120x400_900V_800H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4500 -0.4000 0.4500 0.4000 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4500 -0.4000 0.4500 0.4000 ;
END via7_120x400_900V_800H_ARRAY_2x1

VIA via7_120x400_900V_900H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.4500 -0.4500 0.4500 0.4500 ;
  LAYER v7   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v7   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER m8   ; RECT -0.4500 -0.4500 0.4500 0.4500 ;
END via7_120x400_900V_900H_ARRAY_2x1

VIA VIA8_400X120_180H_540V
  # v8   size: x=0.4000 y=0.1200
  # m8   size: x=0.5200 y=0.1800   enclosure: x=0.0600 y=0.0300
  # gmz   size: x=0.5400 y=0.2400   enclosure: x=0.0700 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.2600 -0.0900 0.2600 0.0900 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER gmz  ; RECT -0.2700 -0.1200 0.2700 0.1200 ;
END VIA8_400X120_180H_540V

VIA VIA8_400X120_180H_721V
  # v8   size: x=0.4000 y=0.1200
  # m8   size: x=0.5200 y=0.1800   enclosure: x=0.0600 y=0.0300
  # gmz   size: x=0.7210 y=0.2900   enclosure: x=0.1605 y=0.0850
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.2600 -0.0900 0.2600 0.0900 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER gmz  ; RECT -0.3605 -0.1450 0.3605 0.1450 ;
END VIA8_400X120_180H_721V

VIA VIA8_400X120_180H_1201V
  # v8   size: x=0.4000 y=0.1200
  # m8   size: x=0.5200 y=0.1800   enclosure: x=0.0600 y=0.0300
  # gmz   size: x=1.2010 y=0.3600   enclosure: x=0.4005 y=0.1200
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.2600 -0.0900 0.2600 0.0900 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER gmz  ; RECT -0.6005 -0.1800 0.6005 0.1800 ;
END VIA8_400X120_180H_1201V

VIA VIA8_400X120_180H_2401V
  # v8   size: x=0.4000 y=0.1200
  # m8   size: x=0.5200 y=0.1800   enclosure: x=0.0600 y=0.0300
  # gmz   size: x=2.4010 y=0.4600   enclosure: x=1.0005 y=0.1700
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.2600 -0.0900 0.2600 0.0900 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER gmz  ; RECT -1.2005 -0.2300 1.2005 0.2300 ;
END VIA8_400X120_180H_2401V

VIA VIA8_120X400_440H_540V
  # v8   size: x=0.1200 y=0.4000
  # m8   size: x=0.2400 y=0.4400   enclosure: x=0.0600 y=0.0200
  # gmz   size: x=0.5400 y=0.5200   enclosure: x=0.2100 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.1200 -0.2200 0.1200 0.2200 ;
  LAYER v8   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gmz  ; RECT -0.2700 -0.2600 0.2700 0.2600 ;
END VIA8_120X400_440H_540V

VIA VIA8_120X400_440H_721V
  # v8   size: x=0.1200 y=0.4000
  # m8   size: x=0.2400 y=0.4400   enclosure: x=0.0600 y=0.0200
  # gmz   size: x=0.7210 y=0.5700   enclosure: x=0.3005 y=0.0850
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.1200 -0.2200 0.1200 0.2200 ;
  LAYER v8   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gmz  ; RECT -0.3605 -0.2850 0.3605 0.2850 ;
END VIA8_120X400_440H_721V

VIA VIA8_120X400_440H_1201V
  # v8   size: x=0.1200 y=0.4000
  # m8   size: x=0.2400 y=0.4400   enclosure: x=0.0600 y=0.0200
  # gmz   size: x=1.2010 y=0.6400   enclosure: x=0.5405 y=0.1200
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.1200 -0.2200 0.1200 0.2200 ;
  LAYER v8   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gmz  ; RECT -0.6005 -0.3200 0.6005 0.3200 ;
END VIA8_120X400_440H_1201V

VIA VIA8_120X400_440H_2401V
  # v8   size: x=0.1200 y=0.4000
  # m8   size: x=0.2400 y=0.4400   enclosure: x=0.0600 y=0.0200
  # gmz   size: x=2.4010 y=0.7400   enclosure: x=1.1405 y=0.1700
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.1200 -0.2200 0.1200 0.2200 ;
  LAYER v8   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gmz  ; RECT -1.2005 -0.3700 1.2005 0.3700 ;
END VIA8_120X400_440H_2401V

VIA VMZ_120X400_540V_540H
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.5400 y=0.5400   enclosure: x=0.2100 y=0.0700
  # gm0   size: x=0.2400 y=0.5400   enclosure: x=0.0600 y=0.0700
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -0.2700 0.2700 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -0.1200 -0.2700 0.1200 0.2700 ;
END VMZ_120X400_540V_540H

VIA VMZ_120X400_540V_721H
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.5400 y=0.5400   enclosure: x=0.2100 y=0.0700
  # gm0   size: x=0.2900 y=0.7210   enclosure: x=0.0850 y=0.1605
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -0.2700 0.2700 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -0.1450 -0.3605 0.1450 0.3605 ;
END VMZ_120X400_540V_721H

VIA VMZ_120X400_540V_1201H
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.5400 y=0.5400   enclosure: x=0.2100 y=0.0700
  # gm0   size: x=0.3600 y=1.2010   enclosure: x=0.1200 y=0.4005
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -0.2700 0.2700 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -0.1800 -0.6005 0.1800 0.6005 ;
END VMZ_120X400_540V_1201H

VIA VMZ_120x400_540V_2130H_ARRAY_1x2
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -1.0650 0.2700 1.0650 ;
  LAYER vmz  ; RECT -0.0600 -0.5200 0.0600 -0.1200 ;
  LAYER vmz  ; RECT -0.0600 0.1200 0.0600 0.5200 ;
  LAYER gm0  ; RECT -0.2700 -1.0650 0.2700 1.0650 ;
END VMZ_120x400_540V_2130H_ARRAY_1x2

VIA VMZ_120X400_540V_2401H
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.5400 y=0.5400   enclosure: x=0.2100 y=0.0700
  # gm0   size: x=0.4600 y=2.4010   enclosure: x=0.1700 y=1.0005
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -0.2700 0.2700 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -0.2300 -1.2005 0.2300 1.2005 ;
END VMZ_120X400_540V_2401H

VIA VMZ_120x400_540V_3980H_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -1.9900 0.2700 1.9900 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -0.2700 -1.9900 0.2700 1.9900 ;
END VMZ_120x400_540V_3980H_ARRAY_1x3

VIA VMZ_120x400_721V_2130H_ARRAY_1x2
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.3610 -1.0650 0.3610 1.0650 ;
  LAYER vmz  ; RECT -0.0600 -0.5200 0.0600 -0.1200 ;
  LAYER vmz  ; RECT -0.0600 0.1200 0.0600 0.5200 ;
  LAYER gm0  ; RECT -0.3610 -1.0650 0.3610 1.0650 ;
END VMZ_120x400_721V_2130H_ARRAY_1x2

VIA VMZ_120x400_721V_3980H_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.3610 -1.9900 0.3610 1.9900 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -0.3610 -1.9900 0.3610 1.9900 ;
END VMZ_120x400_721V_3980H_ARRAY_1x3

VIA VMZ_120x400_1201V_540H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -0.2700 0.6010 0.2700 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gm0  ; RECT -0.6010 -0.2700 0.6010 0.2700 ;
END VMZ_120x400_1201V_540H_ARRAY_2x1

VIA VMZ_120x400_1201V_721H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -0.3610 0.6010 0.3610 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gm0  ; RECT -0.6010 -0.3610 0.6010 0.3610 ;
END VMZ_120x400_1201V_721H_ARRAY_2x1

VIA VMZ_120x400_1201V_1080H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -0.5400 0.6010 0.5400 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gm0  ; RECT -0.6010 -0.5400 0.6010 0.5400 ;
END VMZ_120x400_1201V_1080H_ARRAY_2x1

VIA VMZ_120x400_1201V_1201H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -0.6010 0.6010 0.6010 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gm0  ; RECT -0.6010 -0.6010 0.6010 0.6010 ;
END VMZ_120x400_1201V_1201H_ARRAY_2x1

VIA VMZ_120x400_1201V_2130H_ARRAY_2x2
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -1.0650 0.6010 1.0650 ;
  LAYER vmz  ; RECT -0.2400 -0.5200 -0.1200 -0.1200 ;
  LAYER vmz  ; RECT -0.2400 0.1200 -0.1200 0.5200 ;
  LAYER vmz  ; RECT 0.1200 -0.5200 0.2400 -0.1200 ;
  LAYER vmz  ; RECT 0.1200 0.1200 0.2400 0.5200 ;
  LAYER gm0  ; RECT -0.6010 -1.0650 0.6010 1.0650 ;
END VMZ_120x400_1201V_2130H_ARRAY_2x2

VIA VMZ_120x400_1201V_2401H_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -1.2010 0.6010 1.2010 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gm0  ; RECT -0.6010 -1.2010 0.6010 1.2010 ;
END VMZ_120x400_1201V_2401H_ARRAY_2x1

VIA VMZ_120x400_1201V_3980H_ARRAY_2x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -1.9900 0.6010 1.9900 ;
  LAYER vmz  ; RECT -0.2400 -0.8400 -0.1200 -0.4400 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT -0.2400 0.4400 -0.1200 0.8400 ;
  LAYER vmz  ; RECT 0.1200 -0.8400 0.2400 -0.4400 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.1200 0.4400 0.2400 0.8400 ;
  LAYER gm0  ; RECT -0.6010 -1.9900 0.6010 1.9900 ;
END VMZ_120x400_1201V_3980H_ARRAY_2x3

VIA VMZ_120x400_2401V_540H_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -0.2700 1.2010 0.2700 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -0.2700 1.2010 0.2700 ;
END VMZ_120x400_2401V_540H_ARRAY_6x1

VIA VMZ_120x400_2401V_721H_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -0.3610 1.2010 0.3610 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -0.3610 1.2010 0.3610 ;
END VMZ_120x400_2401V_721H_ARRAY_6x1

VIA VMZ_120x400_2401V_1080H_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -0.5400 1.2010 0.5400 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -0.5400 1.2010 0.5400 ;
END VMZ_120x400_2401V_1080H_ARRAY_6x1

VIA VMZ_120x400_2401V_1201H_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -0.6010 1.2010 0.6010 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -0.6010 1.2010 0.6010 ;
END VMZ_120x400_2401V_1201H_ARRAY_6x1

VIA VMZ_120x400_2401V_2130H_ARRAY_6x2
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -1.0650 1.2010 1.0650 ;
  LAYER vmz  ; RECT -0.9600 -0.5200 -0.8400 -0.1200 ;
  LAYER vmz  ; RECT -0.9600 0.1200 -0.8400 0.5200 ;
  LAYER vmz  ; RECT -0.6000 -0.5200 -0.4800 -0.1200 ;
  LAYER vmz  ; RECT -0.6000 0.1200 -0.4800 0.5200 ;
  LAYER vmz  ; RECT -0.2400 -0.5200 -0.1200 -0.1200 ;
  LAYER vmz  ; RECT -0.2400 0.1200 -0.1200 0.5200 ;
  LAYER vmz  ; RECT 0.1200 -0.5200 0.2400 -0.1200 ;
  LAYER vmz  ; RECT 0.1200 0.1200 0.2400 0.5200 ;
  LAYER vmz  ; RECT 0.4800 -0.5200 0.6000 -0.1200 ;
  LAYER vmz  ; RECT 0.4800 0.1200 0.6000 0.5200 ;
  LAYER vmz  ; RECT 0.8400 -0.5200 0.9600 -0.1200 ;
  LAYER vmz  ; RECT 0.8400 0.1200 0.9600 0.5200 ;
  LAYER gm0  ; RECT -1.2010 -1.0650 1.2010 1.0650 ;
END VMZ_120x400_2401V_2130H_ARRAY_6x2

VIA VMZ_120x400_2401V_2401H_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -1.2010 1.2010 1.2010 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -1.2010 1.2010 1.2010 ;
END VMZ_120x400_2401V_2401H_ARRAY_6x1

VIA VMZ_120x400_2401V_3980H_ARRAY_6x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -1.9900 1.2010 1.9900 ;
  LAYER vmz  ; RECT -0.9600 -0.8400 -0.8400 -0.4400 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.9600 0.4400 -0.8400 0.8400 ;
  LAYER vmz  ; RECT -0.6000 -0.8400 -0.4800 -0.4400 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.6000 0.4400 -0.4800 0.8400 ;
  LAYER vmz  ; RECT -0.2400 -0.8400 -0.1200 -0.4400 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT -0.2400 0.4400 -0.1200 0.8400 ;
  LAYER vmz  ; RECT 0.1200 -0.8400 0.2400 -0.4400 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.1200 0.4400 0.2400 0.8400 ;
  LAYER vmz  ; RECT 0.4800 -0.8400 0.6000 -0.4400 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.4800 0.4400 0.6000 0.8400 ;
  LAYER vmz  ; RECT 0.8400 -0.8400 0.9600 -0.4400 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER vmz  ; RECT 0.8400 0.4400 0.9600 0.8400 ;
  LAYER gm0  ; RECT -1.2010 -1.9900 1.2010 1.9900 ;
END VMZ_120x400_2401V_3980H_ARRAY_6x3

VIA GV0_800X1850_2130H_2000V
  # gv0   size: x=0.8000 y=1.8500
  # gm0   size: x=1.0800 y=2.1300   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=2.0000 y=3.0500   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5400 -1.0650 0.5400 1.0650 ;
  LAYER gv0  ; RECT -0.4000 -0.9250 0.4000 0.9250 ;
  LAYER gmb  ; RECT -1.0000 -1.5250 1.0000 1.5250 ;
END GV0_800X1850_2130H_2000V

VIA GV0_1850X800_1080H_3050V
  # gv0   size: x=1.8500 y=0.8000
  # gm0   size: x=2.1300 y=1.0800   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=3.0500 y=2.0000   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.0650 -0.5400 1.0650 0.5400 ;
  LAYER gv0  ; RECT -0.9250 -0.4000 0.9250 0.4000 ;
  LAYER gmb  ; RECT -1.5250 -1.0000 1.5250 1.0000 ;
END GV0_1850X800_1080H_3050V

VIA GV0_3700X800_1080H_4900V
  # gv0   size: x=3.7000 y=0.8000
  # gm0   size: x=3.9800 y=1.0800   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=4.9000 y=2.0000   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.9900 -0.5400 1.9900 0.5400 ;
  LAYER gv0  ; RECT -1.8500 -0.4000 1.8500 0.4000 ;
  LAYER gmb  ; RECT -2.4500 -1.0000 2.4500 1.0000 ;
END GV0_3700X800_1080H_4900V

VIA GV0_7400X800_1080H_8600V
  # gv0   size: x=7.4000 y=0.8000
  # gm0   size: x=7.6800 y=1.0800   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=8.6000 y=2.0000   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -3.8400 -0.5400 3.8400 0.5400 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -4.3000 -1.0000 4.3000 1.0000 ;
END GV0_7400X800_1080H_8600V

VIA GV0_800X3700_3980H_2000V
  # gv0   size: x=0.8000 y=3.7000
  # gm0   size: x=1.0800 y=3.9800   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=2.0000 y=4.9000   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5400 -1.9900 0.5400 1.9900 ;
  LAYER gv0  ; RECT -0.4000 -1.8500 0.4000 1.8500 ;
  LAYER gmb  ; RECT -1.0000 -2.4500 1.0000 2.4500 ;
END GV0_800X3700_3980H_2000V

VIA GV1_6000X18000_12000V_20000H
  # gv1   size: x=6.0000 y=18.0000
  # gmb   size: x=12.0000 y=24.0000   enclosure: x=3.0000 y=3.0000
  # c4emib   size: x=20.0000 y=20.0000   enclosure: x=7.0000 y=1.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -6.0000 -12.0000 6.0000 12.0000 ;
  LAYER gv1  ; RECT -3.0000 -9.0000 3.0000 9.0000 ;
  LAYER c4emib ; RECT -10.0000 -10.0000 10.0000 10.0000 ;
END GV1_6000X18000_12000V_20000H

VIA GV1_6000X10000_12000V_28000H
  # gv1   size: x=6.0000 y=10.0000
  # gmb   size: x=12.0000 y=16.0000   enclosure: x=3.0000 y=3.0000
  # c4emib   size: x=28.0000 y=28.0000   enclosure: x=11.0000 y=9.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -6.0000 -8.0000 6.0000 8.0000 ;
  LAYER gv1  ; RECT -3.0000 -5.0000 3.0000 5.0000 ;
  LAYER c4emib ; RECT -14.0000 -14.0000 14.0000 14.0000 ;
END GV1_6000X10000_12000V_28000H

VIA GV1_6000X30000_12000V_51000H
  # gv1   size: x=6.0000 y=30.0000
  # gmb   size: x=12.0000 y=36.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=51.0000 y=51.0000   enclosure: x=22.5000 y=10.5000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -6.0000 -18.0000 6.0000 18.0000 ;
  LAYER gv1  ; RECT -3.0000 -15.0000 3.0000 15.0000 ;
  LAYER c4   ; RECT -25.5000 -25.5000 25.5000 25.5000 ;
END GV1_6000X30000_12000V_51000H

VIA GV1_6000X30000_12000V_54000H
  # gv1   size: x=6.0000 y=30.0000
  # gmb   size: x=12.0000 y=36.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=51.0000 y=54.0000   enclosure: x=22.5000 y=12.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -6.0000 -18.0000 6.0000 18.0000 ;
  LAYER gv1  ; RECT -3.0000 -15.0000 3.0000 15.0000 ;
  LAYER c4   ; RECT -25.5000 -27.0000 25.5000 27.0000 ;
END GV1_6000X30000_12000V_54000H

VIA GV1_6000X30000_12000V_85000H
  # gv1   size: x=6.0000 y=30.0000
  # gmb   size: x=12.0000 y=36.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=51.0000 y=85.0000   enclosure: x=22.5000 y=27.5000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -6.0000 -18.0000 6.0000 18.0000 ;
  LAYER gv1  ; RECT -3.0000 -15.0000 3.0000 15.0000 ;
  LAYER c4   ; RECT -25.5000 -42.5000 25.5000 42.5000 ;
END GV1_6000X30000_12000V_85000H

VIA GV0_7400X800_540H_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -0.2700 0.5000 0.2700 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -0.2700 -0.5000 0.2700 0.5000 ;
END GV0_7400X800_540H_1000V_illegal

VIA GV0_7400X800_721H_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -0.3610 0.5000 0.3610 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -0.3610 -0.5000 0.3610 0.5000 ;
END GV0_7400X800_721H_1000V_illegal

VIA GV0_7400X800_1080H_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -0.5400 0.5000 0.5400 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -0.5400 -0.5000 0.5400 0.5000 ;
END GV0_7400X800_1080H_1000V_illegal

VIA GV0_7400X800_1201H_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -0.6010 0.5000 0.6010 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -0.6010 -0.5000 0.6010 0.5000 ;
END GV0_7400X800_1201H_1000V_illegal

VIA GV0_7400X800_2130H_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -1.0650 0.5000 1.0650 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -1.0650 -0.5000 1.0650 0.5000 ;
END GV0_7400X800_2130H_1000V_illegal

VIA GV0_7400X800_2401H_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -1.2010 0.5000 1.2010 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -1.2010 -0.5000 1.2010 0.5000 ;
END GV0_7400X800_2401H_1000V_illegal

VIA GV0_7400X800_3980H_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -1.9900 0.5000 1.9900 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -1.9900 -0.5000 1.9900 0.5000 ;
END GV0_7400X800_3980H_1000V_illegal

##################################################
# Adding extra via which had PGVIA Construct in map table
##################################################
VIA VIA8_400X120_180H_540H
  # v8   size: x=0.4000 y=0.1200
  # m8   size: x=0.5200 y=0.1800   enclosure: x=0.0600 y=0.0300
  # gmz   size: x=0.5200 y=0.5400   enclosure: x=0.0600 y=0.2100
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.2600 -0.0900 0.2600 0.0900 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER gmz  ; RECT -0.2600 -0.2700 0.2600 0.2700 ;
END VIA8_400X120_180H_540H
VIA VIA8_400X120_180H_721H
  # v8   size: x=0.4000 y=0.1200
  # m8   size: x=0.5200 y=0.1800   enclosure: x=0.0600 y=0.0300
  # gmz   size: x=0.5700 y=0.7210   enclosure: x=0.0850 y=0.3005
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.2600 -0.0900 0.2600 0.0900 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER gmz  ; RECT -0.2850 -0.3605 0.2850 0.3605 ;
END VIA8_400X120_180H_721H
VIA VIA8_400X120_180H_1201H
  # v8   size: x=0.4000 y=0.1200
  # m8   size: x=0.5200 y=0.1800   enclosure: x=0.0600 y=0.0300
  # gmz   size: x=0.6400 y=1.2010   enclosure: x=0.1200 y=0.5405
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.2600 -0.0900 0.2600 0.0900 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER gmz  ; RECT -0.3200 -0.6005 0.3200 0.6005 ;
END VIA8_400X120_180H_1201H
VIA via8_400x120_180H_2401V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.0900 1.2010 0.0900 ;
  LAYER v8   ; RECT -0.8400 -0.0600 -0.4400 0.0600 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER v8   ; RECT 0.4400 -0.0600 0.8400 0.0600 ;
  LAYER gmz  ; RECT -1.2010 -0.0900 1.2010 0.0900 ;
END via8_400x120_180H_2401V_ARRAY_3x1
VIA via8_400x120_181H_2401V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.0910 1.2010 0.0910 ;
  LAYER v8   ; RECT -0.8400 -0.0600 -0.4400 0.0600 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER v8   ; RECT 0.4400 -0.0600 0.8400 0.0600 ;
  LAYER gmz  ; RECT -1.2010 -0.0910 1.2010 0.0910 ;
END via8_400x120_181H_2401V_ARRAY_3x1
VIA via8_400x120_190H_2401V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.0950 1.2010 0.0950 ;
  LAYER v8   ; RECT -0.8400 -0.0600 -0.4400 0.0600 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER v8   ; RECT 0.4400 -0.0600 0.8400 0.0600 ;
  LAYER gmz  ; RECT -1.2010 -0.0950 1.2010 0.0950 ;
END via8_400x120_190H_2401V_ARRAY_3x1
VIA via8_400x120_260H_2401V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.1300 1.2010 0.1300 ;
  LAYER v8   ; RECT -0.8400 -0.0600 -0.4400 0.0600 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER v8   ; RECT 0.4400 -0.0600 0.8400 0.0600 ;
  LAYER gmz  ; RECT -1.2010 -0.1300 1.2010 0.1300 ;
END via8_400x120_260H_2401V_ARRAY_3x1
VIA via8_400x120_300H_2401V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.1500 1.2010 0.1500 ;
  LAYER v8   ; RECT -0.8400 -0.0600 -0.4400 0.0600 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER v8   ; RECT 0.4400 -0.0600 0.8400 0.0600 ;
  LAYER gmz  ; RECT -1.2010 -0.1500 1.2010 0.1500 ;
END via8_400x120_300H_2401V_ARRAY_3x1
VIA via8_400x120_400H_2401V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.2000 1.2010 0.2000 ;
  LAYER v8   ; RECT -0.8400 -0.0600 -0.4400 0.0600 ;
  LAYER v8   ; RECT -0.2000 -0.0600 0.2000 0.0600 ;
  LAYER v8   ; RECT 0.4400 -0.0600 0.8400 0.0600 ;
  LAYER gmz  ; RECT -1.2010 -0.2000 1.2010 0.2000 ;
END via8_400x120_400H_2401V_ARRAY_3x1
VIA VIA8_120X400_440H_540H
  # v8   size: x=0.1200 y=0.4000
  # m8   size: x=0.2400 y=0.4400   enclosure: x=0.0600 y=0.0200
  # gmz   size: x=0.2400 y=0.5400   enclosure: x=0.0600 y=0.0700
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.1200 -0.2200 0.1200 0.2200 ;
  LAYER v8   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gmz  ; RECT -0.1200 -0.2700 0.1200 0.2700 ;
END VIA8_120X400_440H_540H
VIA via8_120x400_460H_721V_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.3610 -0.2300 0.3610 0.2300 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gmz  ; RECT -0.3610 -0.2300 0.3610 0.2300 ;
END via8_120x400_460H_721V_ARRAY_2x1
VIA via8_120x400_460H_1201V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.6010 -0.2300 0.6010 0.2300 ;
  LAYER v8   ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER v8   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER v8   ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gmz  ; RECT -0.6010 -0.2300 0.6010 0.2300 ;
END via8_120x400_460H_1201V_ARRAY_3x1
VIA via8_120x400_460H_2401V_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.2300 1.2010 0.2300 ;
  LAYER v8   ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER v8   ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER v8   ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER v8   ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gmz  ; RECT -1.2010 -0.2300 1.2010 0.2300 ;
END via8_120x400_460H_2401V_ARRAY_6x1
VIA via8_120x400_500H_721V_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.3610 -0.2500 0.3610 0.2500 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gmz  ; RECT -0.3610 -0.2500 0.3610 0.2500 ;
END via8_120x400_500H_721V_ARRAY_2x1
VIA via8_120x400_500H_1201V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.6010 -0.2500 0.6010 0.2500 ;
  LAYER v8   ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER v8   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER v8   ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gmz  ; RECT -0.6010 -0.2500 0.6010 0.2500 ;
END via8_120x400_500H_1201V_ARRAY_3x1
VIA via8_120x400_500H_2401V_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.2500 1.2010 0.2500 ;
  LAYER v8   ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER v8   ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER v8   ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER v8   ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gmz  ; RECT -1.2010 -0.2500 1.2010 0.2500 ;
END via8_120x400_500H_2401V_ARRAY_6x1
VIA via8_120x400_600H_721V_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.3610 -0.3000 0.3610 0.3000 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gmz  ; RECT -0.3610 -0.3000 0.3610 0.3000 ;
END via8_120x400_600H_721V_ARRAY_2x1
VIA via8_120x400_600H_1201V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.6010 -0.3000 0.6010 0.3000 ;
  LAYER v8   ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER v8   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER v8   ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gmz  ; RECT -0.6010 -0.3000 0.6010 0.3000 ;
END via8_120x400_600H_1201V_ARRAY_3x1
VIA via8_120x400_600H_2401V_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.3000 1.2010 0.3000 ;
  LAYER v8   ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER v8   ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER v8   ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER v8   ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gmz  ; RECT -1.2010 -0.3000 1.2010 0.3000 ;
END via8_120x400_600H_2401V_ARRAY_6x1
VIA via8_120x400_700H_721V_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.3610 -0.3500 0.3610 0.3500 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gmz  ; RECT -0.3610 -0.3500 0.3610 0.3500 ;
END via8_120x400_700H_721V_ARRAY_2x1
VIA via8_120x400_700H_1201V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.6010 -0.3500 0.6010 0.3500 ;
  LAYER v8   ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER v8   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER v8   ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gmz  ; RECT -0.6010 -0.3500 0.6010 0.3500 ;
END via8_120x400_700H_1201V_ARRAY_3x1
VIA via8_120x400_700H_2401V_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.3500 1.2010 0.3500 ;
  LAYER v8   ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER v8   ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER v8   ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER v8   ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gmz  ; RECT -1.2010 -0.3500 1.2010 0.3500 ;
END via8_120x400_700H_2401V_ARRAY_6x1
VIA via8_120x400_800H_721V_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.3610 -0.4000 0.3610 0.4000 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gmz  ; RECT -0.3610 -0.4000 0.3610 0.4000 ;
END via8_120x400_800H_721V_ARRAY_2x1
VIA via8_120x400_800H_1201V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.6010 -0.4000 0.6010 0.4000 ;
  LAYER v8   ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER v8   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER v8   ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gmz  ; RECT -0.6010 -0.4000 0.6010 0.4000 ;
END via8_120x400_800H_1201V_ARRAY_3x1
VIA via8_120x400_800H_2401V_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.4000 1.2010 0.4000 ;
  LAYER v8   ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER v8   ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER v8   ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER v8   ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gmz  ; RECT -1.2010 -0.4000 1.2010 0.4000 ;
END via8_120x400_800H_2401V_ARRAY_6x1
VIA via8_120x400_900H_721V_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.3610 -0.4500 0.3610 0.4500 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gmz  ; RECT -0.3610 -0.4500 0.3610 0.4500 ;
END via8_120x400_900H_721V_ARRAY_2x1
VIA via8_120x400_900H_1201V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.6010 -0.4500 0.6010 0.4500 ;
  LAYER v8   ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER v8   ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER v8   ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gmz  ; RECT -0.6010 -0.4500 0.6010 0.4500 ;
END via8_120x400_900H_1201V_ARRAY_3x1
VIA via8_120x400_900H_2401V_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -1.2010 -0.4500 1.2010 0.4500 ;
  LAYER v8   ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER v8   ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER v8   ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER v8   ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER v8   ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER v8   ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gmz  ; RECT -1.2010 -0.4500 1.2010 0.4500 ;
END via8_120x400_900H_2401V_ARRAY_6x1
VIA VMZ_120X400_540H_540V
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.3200 y=0.5400   enclosure: x=0.1000 y=0.0700
  # gm0   size: x=0.5400 y=0.5200   enclosure: x=0.2100 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.1600 -0.2700 0.1600 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -0.2700 -0.2600 0.2700 0.2600 ;
END VMZ_120X400_540H_540V
VIA VMZ_120X400_540H_721V
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.3200 y=0.5400   enclosure: x=0.1000 y=0.0700
  # gm0   size: x=0.7210 y=0.5700   enclosure: x=0.3005 y=0.0850
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.1600 -0.2700 0.1600 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -0.3605 -0.2850 0.3605 0.2850 ;
END VMZ_120X400_540H_721V
VIA VMZ_120X400_540H_1201V
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.3200 y=0.5400   enclosure: x=0.1000 y=0.0700
  # gm0   size: x=1.2010 y=0.6400   enclosure: x=0.5405 y=0.1200
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.1600 -0.2700 0.1600 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -0.6005 -0.3200 0.6005 0.3200 ;
END VMZ_120X400_540H_1201V
VIA VMZ_120x400_540H_2130V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.0650 -0.2700 1.0650 0.2700 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gm0  ; RECT -1.0650 -0.2700 1.0650 0.2700 ;
END VMZ_120x400_540H_2130V_ARRAY_3x1
VIA VMZ_120X400_540H_2401V
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.3200 y=0.5400   enclosure: x=0.1000 y=0.0700
  # gm0   size: x=2.4010 y=0.7400   enclosure: x=1.1405 y=0.1700
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.1600 -0.2700 0.1600 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -1.2005 -0.3700 1.2005 0.3700 ;
END VMZ_120X400_540H_2401V
VIA VMZ_120x400_540H_3980V_ARRAY_5x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.9900 -0.2700 1.9900 0.2700 ;
  LAYER vmz  ; RECT -0.7800 -0.2000 -0.6600 0.2000 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER vmz  ; RECT 0.6600 -0.2000 0.7800 0.2000 ;
  LAYER gm0  ; RECT -1.9900 -0.2700 1.9900 0.2700 ;
END VMZ_120x400_540H_3980V_ARRAY_5x1
VIA VMZ_120x400_721H_2130V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.0650 -0.3610 1.0650 0.3610 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gm0  ; RECT -1.0650 -0.3610 1.0650 0.3610 ;
END VMZ_120x400_721H_2130V_ARRAY_3x1
VIA VMZ_120x400_721H_3980V_ARRAY_5x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.9900 -0.3610 1.9900 0.3610 ;
  LAYER vmz  ; RECT -0.7800 -0.2000 -0.6600 0.2000 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER vmz  ; RECT 0.6600 -0.2000 0.7800 0.2000 ;
  LAYER gm0  ; RECT -1.9900 -0.3610 1.9900 0.3610 ;
END VMZ_120x400_721H_3980V_ARRAY_5x1
VIA VMZ_120x400_1201H_540V_ARRAY_1x2
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -0.6010 0.2700 0.6010 ;
  LAYER vmz  ; RECT -0.0600 -0.5200 0.0600 -0.1200 ;
  LAYER vmz  ; RECT -0.0600 0.1200 0.0600 0.5200 ;
  LAYER gm0  ; RECT -0.2700 -0.6010 0.2700 0.6010 ;
END VMZ_120x400_1201H_540V_ARRAY_1x2
VIA VMZ_120x400_1201H_2130V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.0650 -0.6010 1.0650 0.6010 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gm0  ; RECT -1.0650 -0.6010 1.0650 0.6010 ;
END VMZ_120x400_1201H_2130V_ARRAY_3x1
VIA VMZ_120x400_1201H_3980V_ARRAY_5x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.9900 -0.6010 1.9900 0.6010 ;
  LAYER vmz  ; RECT -0.7800 -0.2000 -0.6600 0.2000 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER vmz  ; RECT 0.6600 -0.2000 0.7800 0.2000 ;
  LAYER gm0  ; RECT -1.9900 -0.6010 1.9900 0.6010 ;
END VMZ_120x400_1201H_3980V_ARRAY_5x1
VIA VMZ_120x400_2401H_540V_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -1.2010 0.2700 1.2010 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -0.2700 -1.2010 0.2700 1.2010 ;
END VMZ_120x400_2401H_540V_ARRAY_1x3
VIA VMZ_120x400_2401H_721V_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.3610 -1.2010 0.3610 1.2010 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -0.3610 -1.2010 0.3610 1.2010 ;
END VMZ_120x400_2401H_721V_ARRAY_1x3
VIA VMZ_120x400_2401H_1080V_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.5400 -1.2010 0.5400 1.2010 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -0.5400 -1.2010 0.5400 1.2010 ;
END VMZ_120x400_2401H_1080V_ARRAY_1x3
VIA VMZ_120x400_2401H_1201V_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -1.2010 0.6010 1.2010 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -0.6010 -1.2010 0.6010 1.2010 ;
END VMZ_120x400_2401H_1201V_ARRAY_1x3
VIA VMZ_120x400_2401H_2130V_ARRAY_3x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.0650 -1.2010 1.0650 1.2010 ;
  LAYER vmz  ; RECT -0.4200 -0.8400 -0.3000 -0.4400 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.4200 0.4400 -0.3000 0.8400 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER vmz  ; RECT 0.3000 -0.8400 0.4200 -0.4400 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER vmz  ; RECT 0.3000 0.4400 0.4200 0.8400 ;
  LAYER gm0  ; RECT -1.0650 -1.2010 1.0650 1.2010 ;
END VMZ_120x400_2401H_2130V_ARRAY_3x3
VIA VMZ_120x400_2401H_2401V_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -1.2010 1.2010 1.2010 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -1.2010 -1.2010 1.2010 1.2010 ;
END VMZ_120x400_2401H_2401V_ARRAY_1x3
VIA VMZ_120x400_2401H_3980V_ARRAY_5x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.9900 -1.2010 1.9900 1.2010 ;
  LAYER vmz  ; RECT -0.7800 -0.8400 -0.6600 -0.4400 ;
  LAYER vmz  ; RECT -0.7800 -0.2000 -0.6600 0.2000 ;
  LAYER vmz  ; RECT -0.7800 0.4400 -0.6600 0.8400 ;
  LAYER vmz  ; RECT -0.4200 -0.8400 -0.3000 -0.4400 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.4200 0.4400 -0.3000 0.8400 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER vmz  ; RECT 0.3000 -0.8400 0.4200 -0.4400 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER vmz  ; RECT 0.3000 0.4400 0.4200 0.8400 ;
  LAYER vmz  ; RECT 0.6600 -0.8400 0.7800 -0.4400 ;
  LAYER vmz  ; RECT 0.6600 -0.2000 0.7800 0.2000 ;
  LAYER vmz  ; RECT 0.6600 0.4400 0.7800 0.8400 ;
  LAYER gm0  ; RECT -1.9900 -1.2010 1.9900 1.2010 ;
END VMZ_120x400_2401H_3980V_ARRAY_5x3
VIA GV0_1850X800_2130V_2000H
  # gv0   size: x=1.8500 y=0.8000
  # gm0   size: x=2.1300 y=1.0800   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=3.0500 y=2.0000   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.0650 -0.5400 1.0650 0.5400 ;
  LAYER gv0  ; RECT -0.9250 -0.4000 0.9250 0.4000 ;
  LAYER gmb  ; RECT -1.5250 -1.0000 1.5250 1.0000 ;
END GV0_1850X800_2130V_2000H
VIA GV0_800X1850_1080V_3050H
  # gv0   size: x=0.8000 y=1.8500
  # gm0   size: x=1.0800 y=2.1300   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=2.0000 y=3.0500   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5400 -1.0650 0.5400 1.0650 ;
  LAYER gv0  ; RECT -0.4000 -0.9250 0.4000 0.9250 ;
  LAYER gmb  ; RECT -1.0000 -1.5250 1.0000 1.5250 ;
END GV0_800X1850_1080V_3050H
VIA GV0_800X3700_1080V_4900H
  # gv0   size: x=0.8000 y=3.7000
  # gm0   size: x=1.0800 y=3.9800   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=2.0000 y=4.9000   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5400 -1.9900 0.5400 1.9900 ;
  LAYER gv0  ; RECT -0.4000 -1.8500 0.4000 1.8500 ;
  LAYER gmb  ; RECT -1.0000 -2.4500 1.0000 2.4500 ;
END GV0_800X3700_1080V_4900H
VIA GV0_800X7400_1080V_8600H
  # gv0   size: x=0.8000 y=7.4000
  # gm0   size: x=1.0800 y=7.6800   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=2.0000 y=8.6000   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5400 -3.8400 0.5400 3.8400 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -1.0000 -4.3000 1.0000 4.3000 ;
END GV0_800X7400_1080V_8600H
VIA GV0_3700X800_3980V_2000H
  # gv0   size: x=3.7000 y=0.8000
  # gm0   size: x=3.9800 y=1.0800   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=4.9000 y=2.0000   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.9900 -0.5400 1.9900 0.5400 ;
  LAYER gv0  ; RECT -1.8500 -0.4000 1.8500 0.4000 ;
  LAYER gmb  ; RECT -2.4500 -1.0000 2.4500 1.0000 ;
END GV0_3700X800_3980V_2000H
VIA GV0_3700x800_3980V_4900H_ARRAY_1x2
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.9900 -2.4500 1.9900 2.4500 ;
  LAYER gv0  ; RECT -1.8500 -1.8000 1.8500 -1.0000 ;
  LAYER gv0  ; RECT -1.8500 1.0000 1.8500 1.8000 ;
  LAYER gmb  ; RECT -1.9900 -2.4500 1.9900 2.4500 ;
END GV0_3700x800_3980V_4900H_ARRAY_1x2
VIA GV1_18000X6000_12000H_20000V
  # gv1   size: x=18.0000 y=6.0000
  # gmb   size: x=24.0000 y=12.0000   enclosure: x=3.0000 y=3.0000
  # c4emib   size: x=20.0000 y=20.0000   enclosure: x=1.0000 y=7.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -12.0000 -6.0000 12.0000 6.0000 ;
  LAYER gv1  ; RECT -9.0000 -3.0000 9.0000 3.0000 ;
  LAYER c4emib ; RECT -10.0000 -10.0000 10.0000 10.0000 ;
END GV1_18000X6000_12000H_20000V
VIA GV1_10000X6000_12000H_28000V
  # gv1   size: x=10.0000 y=6.0000
  # gmb   size: x=16.0000 y=12.0000   enclosure: x=3.0000 y=3.0000
  # c4emib   size: x=28.0000 y=28.0000   enclosure: x=9.0000 y=11.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -8.0000 -6.0000 8.0000 6.0000 ;
  LAYER gv1  ; RECT -5.0000 -3.0000 5.0000 3.0000 ;
  LAYER c4emib ; RECT -14.0000 -14.0000 14.0000 14.0000 ;
END GV1_10000X6000_12000H_28000V
VIA GV1_30000X6000_12000H_51000V
  # gv1   size: x=30.0000 y=6.0000
  # gmb   size: x=36.0000 y=12.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=51.0000 y=51.0000   enclosure: x=10.5000 y=22.5000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -18.0000 -6.0000 18.0000 6.0000 ;
  LAYER gv1  ; RECT -15.0000 -3.0000 15.0000 3.0000 ;
  LAYER c4   ; RECT -25.5000 -25.5000 25.5000 25.5000 ;
END GV1_30000X6000_12000H_51000V
VIA GV1_30000X6000_12000H_54000V
  # gv1   size: x=30.0000 y=6.0000
  # gmb   size: x=36.0000 y=12.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=54.0000 y=51.0000   enclosure: x=12.0000 y=22.5000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -18.0000 -6.0000 18.0000 6.0000 ;
  LAYER gv1  ; RECT -15.0000 -3.0000 15.0000 3.0000 ;
  LAYER c4   ; RECT -27.0000 -25.5000 27.0000 25.5000 ;
END GV1_30000X6000_12000H_54000V
VIA GV1_30000X6000_12000H_85000V
  # gv1   size: x=30.0000 y=6.0000
  # gmb   size: x=36.0000 y=12.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=85.0000 y=51.0000   enclosure: x=27.5000 y=22.5000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -18.0000 -6.0000 18.0000 6.0000 ;
  LAYER gv1  ; RECT -15.0000 -3.0000 15.0000 3.0000 ;
  LAYER c4   ; RECT -42.5000 -25.5000 42.5000 25.5000 ;
END GV1_30000X6000_12000H_85000V
VIA GV0_800X7400_540V_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.2700 -0.5000 0.2700 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -0.2700 0.5000 0.2700 ;
END GV0_800X7400_540V_1000H_illegal
VIA GV0_800X7400_721V_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.3610 -0.5000 0.3610 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -0.3610 0.5000 0.3610 ;
END GV0_800X7400_721V_1000H_illegal
VIA GV0_800X7400_1080V_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5400 -0.5000 0.5400 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -0.5400 0.5000 0.5400 ;
END GV0_800X7400_1080V_1000H_illegal
VIA GV0_800X7400_1201V_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.6010 -0.5000 0.6010 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -0.6010 0.5000 0.6010 ;
END GV0_800X7400_1201V_1000H_illegal
VIA GV0_800X7400_2130V_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.0650 -0.5000 1.0650 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -1.0650 0.5000 1.0650 ;
END GV0_800X7400_2130V_1000H_illegal
VIA GV0_800X7400_2401V_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.2010 -0.5000 1.2010 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -1.2010 0.5000 1.2010 ;
END GV0_800X7400_2401V_1000H_illegal
VIA GV0_800X7400_3980V_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.9900 -0.5000 1.9900 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -1.9900 0.5000 1.9900 ;
END GV0_800X7400_3980V_1000H_illegal
VIA VMZ_120X400_540H_540H
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.3200 y=0.5400   enclosure: x=0.1000 y=0.0700
  # gm0   size: x=0.2400 y=0.5400   enclosure: x=0.0600 y=0.0700
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.1600 -0.2700 0.1600 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -0.1200 -0.2700 0.1200 0.2700 ;
END VMZ_120X400_540H_540H
VIA VMZ_120x400_540H_721V_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.3610 -0.2700 0.3610 0.2700 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gm0  ; RECT -0.3610 -0.2700 0.3610 0.2700 ;
END VMZ_120x400_540H_721V_ARRAY_2x1
VIA VMZ_120x400_540H_1080V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.5400 -0.2700 0.5400 0.2700 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gm0  ; RECT -0.5400 -0.2700 0.5400 0.2700 ;
END VMZ_120x400_540H_1080V_ARRAY_3x1
VIA VMZ_120x400_540H_1201V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -0.2700 0.6010 0.2700 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gm0  ; RECT -0.6010 -0.2700 0.6010 0.2700 ;
END VMZ_120x400_540H_1201V_ARRAY_3x1
VIA VMZ_120x400_540H_2130V_ARRAY_5x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.0650 -0.2700 1.0650 0.2700 ;
  LAYER vmz  ; RECT -0.7800 -0.2000 -0.6600 0.2000 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER vmz  ; RECT 0.6600 -0.2000 0.7800 0.2000 ;
  LAYER gm0  ; RECT -1.0650 -0.2700 1.0650 0.2700 ;
END VMZ_120x400_540H_2130V_ARRAY_5x1
VIA VMZ_120x400_540H_2401V_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -0.2700 1.2010 0.2700 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -0.2700 1.2010 0.2700 ;
END VMZ_120x400_540H_2401V_ARRAY_6x1
VIA VMZ_120x400_540H_3980V_ARRAY_10x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.9900 -0.2700 1.9900 0.2700 ;
  LAYER vmz  ; RECT -1.6800 -0.2000 -1.5600 0.2000 ;
  LAYER vmz  ; RECT -1.3200 -0.2000 -1.2000 0.2000 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER vmz  ; RECT 1.2000 -0.2000 1.3200 0.2000 ;
  LAYER vmz  ; RECT 1.5600 -0.2000 1.6800 0.2000 ;
  LAYER gm0  ; RECT -1.9900 -0.2700 1.9900 0.2700 ;
END VMZ_120x400_540H_3980V_ARRAY_10x1
VIA VMZ_120x400_721H_721V_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.3610 -0.3610 0.3610 0.3610 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gm0  ; RECT -0.3610 -0.3610 0.3610 0.3610 ;
END VMZ_120x400_721H_721V_ARRAY_2x1
VIA VMZ_120x400_721H_1080V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.5400 -0.3610 0.5400 0.3610 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gm0  ; RECT -0.5400 -0.3610 0.5400 0.3610 ;
END VMZ_120x400_721H_1080V_ARRAY_3x1
VIA VMZ_120x400_721H_1201V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -0.3610 0.6010 0.3610 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gm0  ; RECT -0.6010 -0.3610 0.6010 0.3610 ;
END VMZ_120x400_721H_1201V_ARRAY_3x1
VIA VMZ_120x400_721H_2130V_ARRAY_5x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.0650 -0.3610 1.0650 0.3610 ;
  LAYER vmz  ; RECT -0.7800 -0.2000 -0.6600 0.2000 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER vmz  ; RECT 0.6600 -0.2000 0.7800 0.2000 ;
  LAYER gm0  ; RECT -1.0650 -0.3610 1.0650 0.3610 ;
END VMZ_120x400_721H_2130V_ARRAY_5x1
VIA VMZ_120x400_721H_2401V_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -0.3610 1.2010 0.3610 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -0.3610 1.2010 0.3610 ;
END VMZ_120x400_721H_2401V_ARRAY_6x1
VIA VMZ_120x400_721H_3980V_ARRAY_10x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.9900 -0.3610 1.9900 0.3610 ;
  LAYER vmz  ; RECT -1.6800 -0.2000 -1.5600 0.2000 ;
  LAYER vmz  ; RECT -1.3200 -0.2000 -1.2000 0.2000 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER vmz  ; RECT 1.2000 -0.2000 1.3200 0.2000 ;
  LAYER vmz  ; RECT 1.5600 -0.2000 1.6800 0.2000 ;
  LAYER gm0  ; RECT -1.9900 -0.3610 1.9900 0.3610 ;
END VMZ_120x400_721H_3980V_ARRAY_10x1
VIA VMZ_120x400_1201H_721V_ARRAY_2x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.3610 -0.6010 0.3610 0.6010 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER gm0  ; RECT -0.3610 -0.6010 0.3610 0.6010 ;
END VMZ_120x400_1201H_721V_ARRAY_2x1
VIA VMZ_120x400_1201H_1080V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.5400 -0.6010 0.5400 0.6010 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gm0  ; RECT -0.5400 -0.6010 0.5400 0.6010 ;
END VMZ_120x400_1201H_1080V_ARRAY_3x1
VIA VMZ_120x400_1201H_1201V_ARRAY_3x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -0.6010 0.6010 0.6010 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER gm0  ; RECT -0.6010 -0.6010 0.6010 0.6010 ;
END VMZ_120x400_1201H_1201V_ARRAY_3x1
VIA VMZ_120x400_1201H_2130V_ARRAY_5x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.0650 -0.6010 1.0650 0.6010 ;
  LAYER vmz  ; RECT -0.7800 -0.2000 -0.6600 0.2000 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER vmz  ; RECT 0.6600 -0.2000 0.7800 0.2000 ;
  LAYER gm0  ; RECT -1.0650 -0.6010 1.0650 0.6010 ;
END VMZ_120x400_1201H_2130V_ARRAY_5x1
VIA VMZ_120x400_1201H_2401V_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -0.6010 1.2010 0.6010 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -0.6010 1.2010 0.6010 ;
END VMZ_120x400_1201H_2401V_ARRAY_6x1
VIA VMZ_120x400_1201H_3980V_ARRAY_10x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.9900 -0.6010 1.9900 0.6010 ;
  LAYER vmz  ; RECT -1.6800 -0.2000 -1.5600 0.2000 ;
  LAYER vmz  ; RECT -1.3200 -0.2000 -1.2000 0.2000 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER vmz  ; RECT 1.2000 -0.2000 1.3200 0.2000 ;
  LAYER vmz  ; RECT 1.5600 -0.2000 1.6800 0.2000 ;
  LAYER gm0  ; RECT -1.9900 -0.6010 1.9900 0.6010 ;
END VMZ_120x400_1201H_3980V_ARRAY_10x1
VIA VMZ_120x400_2401H_721V_ARRAY_2x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.3610 -1.2010 0.3610 1.2010 ;
  LAYER vmz  ; RECT -0.2400 -0.8400 -0.1200 -0.4400 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT -0.2400 0.4400 -0.1200 0.8400 ;
  LAYER vmz  ; RECT 0.1200 -0.8400 0.2400 -0.4400 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.1200 0.4400 0.2400 0.8400 ;
  LAYER gm0  ; RECT -0.3610 -1.2010 0.3610 1.2010 ;
END VMZ_120x400_2401H_721V_ARRAY_2x3
VIA VMZ_120x400_2401H_1080V_ARRAY_3x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.5400 -1.2010 0.5400 1.2010 ;
  LAYER vmz  ; RECT -0.4200 -0.8400 -0.3000 -0.4400 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.4200 0.4400 -0.3000 0.8400 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER vmz  ; RECT 0.3000 -0.8400 0.4200 -0.4400 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER vmz  ; RECT 0.3000 0.4400 0.4200 0.8400 ;
  LAYER gm0  ; RECT -0.5400 -1.2010 0.5400 1.2010 ;
END VMZ_120x400_2401H_1080V_ARRAY_3x3
VIA VMZ_120x400_2401H_1201V_ARRAY_3x2
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -1.2010 0.6010 1.2010 ;
  LAYER vmz  ; RECT -0.4200 -0.5200 -0.3000 -0.1200 ;
  LAYER vmz  ; RECT -0.4200 0.1200 -0.3000 0.5200 ;
  LAYER vmz  ; RECT -0.0600 -0.5200 0.0600 -0.1200 ;
  LAYER vmz  ; RECT -0.0600 0.1200 0.0600 0.5200 ;
  LAYER vmz  ; RECT 0.3000 -0.5200 0.4200 -0.1200 ;
  LAYER vmz  ; RECT 0.3000 0.1200 0.4200 0.5200 ;
  LAYER gm0  ; RECT -0.6010 -1.2010 0.6010 1.2010 ;
END VMZ_120x400_2401H_1201V_ARRAY_3x2
VIA VMZ_120x400_2401H_2130V_ARRAY_5x2
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.0650 -1.2010 1.0650 1.2010 ;
  LAYER vmz  ; RECT -0.7800 -0.5200 -0.6600 -0.1200 ;
  LAYER vmz  ; RECT -0.7800 0.1200 -0.6600 0.5200 ;
  LAYER vmz  ; RECT -0.4200 -0.5200 -0.3000 -0.1200 ;
  LAYER vmz  ; RECT -0.4200 0.1200 -0.3000 0.5200 ;
  LAYER vmz  ; RECT -0.0600 -0.5200 0.0600 -0.1200 ;
  LAYER vmz  ; RECT -0.0600 0.1200 0.0600 0.5200 ;
  LAYER vmz  ; RECT 0.3000 -0.5200 0.4200 -0.1200 ;
  LAYER vmz  ; RECT 0.3000 0.1200 0.4200 0.5200 ;
  LAYER vmz  ; RECT 0.6600 -0.5200 0.7800 -0.1200 ;
  LAYER vmz  ; RECT 0.6600 0.1200 0.7800 0.5200 ;
  LAYER gm0  ; RECT -1.0650 -1.2010 1.0650 1.2010 ;
END VMZ_120x400_2401H_2130V_ARRAY_5x2
VIA VMZ_120x400_2401H_2401V_ARRAY_6x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -1.2010 1.2010 1.2010 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -1.2010 1.2010 1.2010 ;
END VMZ_120x400_2401H_2401V_ARRAY_6x1
VIA VMZ_120x400_2401H_3980V_ARRAY_10x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.9900 -1.2010 1.9900 1.2010 ;
  LAYER vmz  ; RECT -1.6800 -0.2000 -1.5600 0.2000 ;
  LAYER vmz  ; RECT -1.3200 -0.2000 -1.2000 0.2000 ;
  LAYER vmz  ; RECT -0.9600 -0.2000 -0.8400 0.2000 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.8400 -0.2000 0.9600 0.2000 ;
  LAYER vmz  ; RECT 1.2000 -0.2000 1.3200 0.2000 ;
  LAYER vmz  ; RECT 1.5600 -0.2000 1.6800 0.2000 ;
  LAYER gm0  ; RECT -1.9900 -1.2010 1.9900 1.2010 ;
END VMZ_120x400_2401H_3980V_ARRAY_10x1
VIA GV0_7400X800_1080H_2000H
  # gv0   size: x=7.4000 y=0.8000
  # gm0   size: x=7.6800 y=1.0800   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=8.6000 y=2.0000   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -3.8400 -0.5400 3.8400 0.5400 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -4.3000 -1.0000 4.3000 1.0000 ;
END GV0_7400X800_1080H_2000H
VIA GV1_18000X6000_12000H_20000H
  # gv1   size: x=18.0000 y=6.0000
  # gmb   size: x=24.0000 y=12.0000   enclosure: x=3.0000 y=3.0000
  # c4emib   size: x=20.0000 y=20.0000   enclosure: x=1.0000 y=7.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -12.0000 -6.0000 12.0000 6.0000 ;
  LAYER gv1  ; RECT -9.0000 -3.0000 9.0000 3.0000 ;
  LAYER c4emib ; RECT -10.0000 -10.0000 10.0000 10.0000 ;
END GV1_18000X6000_12000H_20000H
VIA GV1_10000X6000_12000H_28000H
  # gv1   size: x=10.0000 y=6.0000
  # gmb   size: x=16.0000 y=12.0000   enclosure: x=3.0000 y=3.0000
  # c4emib   size: x=28.0000 y=28.0000   enclosure: x=9.0000 y=11.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -8.0000 -6.0000 8.0000 6.0000 ;
  LAYER gv1  ; RECT -5.0000 -3.0000 5.0000 3.0000 ;
  LAYER c4emib ; RECT -14.0000 -14.0000 14.0000 14.0000 ;
END GV1_10000X6000_12000H_28000H
VIA GV1_30000X6000_12000H_51000H
  # gv1   size: x=30.0000 y=6.0000
  # gmb   size: x=36.0000 y=12.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=51.0000 y=51.0000   enclosure: x=10.5000 y=22.5000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -18.0000 -6.0000 18.0000 6.0000 ;
  LAYER gv1  ; RECT -15.0000 -3.0000 15.0000 3.0000 ;
  LAYER c4   ; RECT -25.5000 -25.5000 25.5000 25.5000 ;
END GV1_30000X6000_12000H_51000H
VIA GV1_30000X6000_12000H_54000H
  # gv1   size: x=30.0000 y=6.0000
  # gmb   size: x=36.0000 y=12.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=51.0000 y=54.0000   enclosure: x=10.5000 y=24.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -18.0000 -6.0000 18.0000 6.0000 ;
  LAYER gv1  ; RECT -15.0000 -3.0000 15.0000 3.0000 ;
  LAYER c4   ; RECT -25.5000 -27.0000 25.5000 27.0000 ;
END GV1_30000X6000_12000H_54000H
VIA GV1_30000X6000_12000H_85000H
  # gv1   size: x=30.0000 y=6.0000
  # gmb   size: x=36.0000 y=12.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=51.0000 y=85.0000   enclosure: x=10.5000 y=39.5000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -18.0000 -6.0000 18.0000 6.0000 ;
  LAYER gv1  ; RECT -15.0000 -3.0000 15.0000 3.0000 ;
  LAYER c4   ; RECT -25.5000 -42.5000 25.5000 42.5000 ;
END GV1_30000X6000_12000H_85000H
VIA GV0_7400X800_540H_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -0.2700 0.5000 0.2700 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -0.2700 -0.5000 0.2700 0.5000 ;
END GV0_7400X800_540H_1000H_illegal
VIA GV0_7400X800_721H_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -0.3610 0.5000 0.3610 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -0.3610 -0.5000 0.3610 0.5000 ;
END GV0_7400X800_721H_1000H_illegal
VIA GV0_7400X800_1080H_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -0.5400 0.5000 0.5400 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -0.5400 -0.5000 0.5400 0.5000 ;
END GV0_7400X800_1080H_1000H_illegal
VIA GV0_7400X800_1201H_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -0.6010 0.5000 0.6010 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -0.6010 -0.5000 0.6010 0.5000 ;
END GV0_7400X800_1201H_1000H_illegal
VIA GV0_7400X800_2130H_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -1.0650 0.5000 1.0650 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -1.0650 -0.5000 1.0650 0.5000 ;
END GV0_7400X800_2130H_1000H_illegal
VIA GV0_7400X800_2401H_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -1.2010 0.5000 1.2010 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -1.2010 -0.5000 1.2010 0.5000 ;
END GV0_7400X800_2401H_1000H_illegal
VIA GV0_7400X800_3980H_1000H_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5000 -1.9900 0.5000 1.9900 ;
  LAYER gv0  ; RECT -3.7000 -0.4000 3.7000 0.4000 ;
  LAYER gmb  ; RECT -1.9900 -0.5000 1.9900 0.5000 ;
END GV0_7400X800_3980H_1000H_illegal
VIA VMZ_120X400_540V_540V
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.5400 y=0.5400   enclosure: x=0.2100 y=0.0700
  # gm0   size: x=0.5400 y=0.5200   enclosure: x=0.2100 y=0.0600
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -0.2700 0.2700 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -0.2700 -0.2600 0.2700 0.2600 ;
END VMZ_120X400_540V_540V
VIA VMZ_120X400_540V_721V
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.5400 y=0.5400   enclosure: x=0.2100 y=0.0700
  # gm0   size: x=0.7210 y=0.5700   enclosure: x=0.3005 y=0.0850
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -0.2700 0.2700 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -0.3605 -0.2850 0.3605 0.2850 ;
END VMZ_120X400_540V_721V
VIA VMZ_120X400_540V_1201V
  # vmz   size: x=0.1200 y=0.4000
  # gmz   size: x=0.5400 y=0.5400   enclosure: x=0.2100 y=0.0700
  # gm0   size: x=1.2010 y=0.6400   enclosure: x=0.5405 y=0.1200
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -0.2700 0.2700 0.2700 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER gm0  ; RECT -0.6005 -0.3200 0.6005 0.3200 ;
END VMZ_120X400_540V_1201V
VIA VMZ_120x400_540V_2130H_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -1.0650 0.2700 1.0650 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -0.2700 -1.0650 0.2700 1.0650 ;
END VMZ_120x400_540V_2130H_ARRAY_1x3
VIA VMZ_120x400_540V_2401H_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -1.2010 0.2700 1.2010 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -0.2700 -1.2010 0.2700 1.2010 ;
END VMZ_120x400_540V_2401H_ARRAY_1x3
VIA VMZ_120x400_540V_3980H_ARRAY_1x6
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.2700 -1.9900 0.2700 1.9900 ;
  LAYER vmz  ; RECT -0.0600 -1.8000 0.0600 -1.4000 ;
  LAYER vmz  ; RECT -0.0600 -1.1600 0.0600 -0.7600 ;
  LAYER vmz  ; RECT -0.0600 -0.5200 0.0600 -0.1200 ;
  LAYER vmz  ; RECT -0.0600 0.1200 0.0600 0.5200 ;
  LAYER vmz  ; RECT -0.0600 0.7600 0.0600 1.1600 ;
  LAYER vmz  ; RECT -0.0600 1.4000 0.0600 1.8000 ;
  LAYER gm0  ; RECT -0.2700 -1.9900 0.2700 1.9900 ;
END VMZ_120x400_540V_3980H_ARRAY_1x6
VIA VMZ_120x400_721V_2130H_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.3610 -1.0650 0.3610 1.0650 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -0.3610 -1.0650 0.3610 1.0650 ;
END VMZ_120x400_721V_2130H_ARRAY_1x3
VIA VMZ_120x400_721V_2401H_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.3610 -1.2010 0.3610 1.2010 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -0.3610 -1.2010 0.3610 1.2010 ;
END VMZ_120x400_721V_2401H_ARRAY_1x3
VIA VMZ_120x400_721V_3980H_ARRAY_1x6
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.3610 -1.9900 0.3610 1.9900 ;
  LAYER vmz  ; RECT -0.0600 -1.8000 0.0600 -1.4000 ;
  LAYER vmz  ; RECT -0.0600 -1.1600 0.0600 -0.7600 ;
  LAYER vmz  ; RECT -0.0600 -0.5200 0.0600 -0.1200 ;
  LAYER vmz  ; RECT -0.0600 0.1200 0.0600 0.5200 ;
  LAYER vmz  ; RECT -0.0600 0.7600 0.0600 1.1600 ;
  LAYER vmz  ; RECT -0.0600 1.4000 0.0600 1.8000 ;
  LAYER gm0  ; RECT -0.3610 -1.9900 0.3610 1.9900 ;
END VMZ_120x400_721V_3980H_ARRAY_1x6
VIA VMZ_120x400_1201V_2130H_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -1.0650 0.6010 1.0650 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -0.6010 -1.0650 0.6010 1.0650 ;
END VMZ_120x400_1201V_2130H_ARRAY_1x3
VIA VMZ_120x400_1201V_2401H_ARRAY_2x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -1.2010 0.6010 1.2010 ;
  LAYER vmz  ; RECT -0.2400 -0.8400 -0.1200 -0.4400 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT -0.2400 0.4400 -0.1200 0.8400 ;
  LAYER vmz  ; RECT 0.1200 -0.8400 0.2400 -0.4400 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.1200 0.4400 0.2400 0.8400 ;
  LAYER gm0  ; RECT -0.6010 -1.2010 0.6010 1.2010 ;
END VMZ_120x400_1201V_2401H_ARRAY_2x3
VIA VMZ_120x400_1201V_3980H_ARRAY_2x6
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.6010 -1.9900 0.6010 1.9900 ;
  LAYER vmz  ; RECT -0.2400 -1.8000 -0.1200 -1.4000 ;
  LAYER vmz  ; RECT -0.2400 -1.1600 -0.1200 -0.7600 ;
  LAYER vmz  ; RECT -0.2400 -0.5200 -0.1200 -0.1200 ;
  LAYER vmz  ; RECT -0.2400 0.1200 -0.1200 0.5200 ;
  LAYER vmz  ; RECT -0.2400 0.7600 -0.1200 1.1600 ;
  LAYER vmz  ; RECT -0.2400 1.4000 -0.1200 1.8000 ;
  LAYER vmz  ; RECT 0.1200 -1.8000 0.2400 -1.4000 ;
  LAYER vmz  ; RECT 0.1200 -1.1600 0.2400 -0.7600 ;
  LAYER vmz  ; RECT 0.1200 -0.5200 0.2400 -0.1200 ;
  LAYER vmz  ; RECT 0.1200 0.1200 0.2400 0.5200 ;
  LAYER vmz  ; RECT 0.1200 0.7600 0.2400 1.1600 ;
  LAYER vmz  ; RECT 0.1200 1.4000 0.2400 1.8000 ;
  LAYER gm0  ; RECT -0.6010 -1.9900 0.6010 1.9900 ;
END VMZ_120x400_1201V_3980H_ARRAY_2x6
VIA VMZ_120x400_2401V_721H_ARRAY_5x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -0.3610 1.2010 0.3610 ;
  LAYER vmz  ; RECT -0.7800 -0.2000 -0.6600 0.2000 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER vmz  ; RECT 0.6600 -0.2000 0.7800 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -0.3610 1.2010 0.3610 ;
END VMZ_120x400_2401V_721H_ARRAY_5x1
VIA VMZ_120x400_2401V_1080H_ARRAY_5x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -0.5400 1.2010 0.5400 ;
  LAYER vmz  ; RECT -0.7800 -0.2000 -0.6600 0.2000 ;
  LAYER vmz  ; RECT -0.4200 -0.2000 -0.3000 0.2000 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT 0.3000 -0.2000 0.4200 0.2000 ;
  LAYER vmz  ; RECT 0.6600 -0.2000 0.7800 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -0.5400 1.2010 0.5400 ;
END VMZ_120x400_2401V_1080H_ARRAY_5x1
VIA VMZ_120x400_2401V_1201H_ARRAY_4x1
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -0.6010 1.2010 0.6010 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER gm0  ; RECT -1.2010 -0.6010 1.2010 0.6010 ;
END VMZ_120x400_2401V_1201H_ARRAY_4x1
VIA VMZ_120x400_2401V_2130H_ARRAY_4x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -1.0650 1.2010 1.0650 ;
  LAYER vmz  ; RECT -0.6000 -0.8400 -0.4800 -0.4400 ;
  LAYER vmz  ; RECT -0.6000 -0.2000 -0.4800 0.2000 ;
  LAYER vmz  ; RECT -0.6000 0.4400 -0.4800 0.8400 ;
  LAYER vmz  ; RECT -0.2400 -0.8400 -0.1200 -0.4400 ;
  LAYER vmz  ; RECT -0.2400 -0.2000 -0.1200 0.2000 ;
  LAYER vmz  ; RECT -0.2400 0.4400 -0.1200 0.8400 ;
  LAYER vmz  ; RECT 0.1200 -0.8400 0.2400 -0.4400 ;
  LAYER vmz  ; RECT 0.1200 -0.2000 0.2400 0.2000 ;
  LAYER vmz  ; RECT 0.1200 0.4400 0.2400 0.8400 ;
  LAYER vmz  ; RECT 0.4800 -0.8400 0.6000 -0.4400 ;
  LAYER vmz  ; RECT 0.4800 -0.2000 0.6000 0.2000 ;
  LAYER vmz  ; RECT 0.4800 0.4400 0.6000 0.8400 ;
  LAYER gm0  ; RECT -1.2010 -1.0650 1.2010 1.0650 ;
END VMZ_120x400_2401V_2130H_ARRAY_4x3
VIA VMZ_120x400_2401V_2401H_ARRAY_1x3
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -1.2010 1.2010 1.2010 ;
  LAYER vmz  ; RECT -0.0600 -0.8400 0.0600 -0.4400 ;
  LAYER vmz  ; RECT -0.0600 -0.2000 0.0600 0.2000 ;
  LAYER vmz  ; RECT -0.0600 0.4400 0.0600 0.8400 ;
  LAYER gm0  ; RECT -1.2010 -1.2010 1.2010 1.2010 ;
END VMZ_120x400_2401V_2401H_ARRAY_1x3
VIA VMZ_120x400_2401V_3980H_ARRAY_1x6
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -1.2010 -1.9900 1.2010 1.9900 ;
  LAYER vmz  ; RECT -0.0600 -1.8000 0.0600 -1.4000 ;
  LAYER vmz  ; RECT -0.0600 -1.1600 0.0600 -0.7600 ;
  LAYER vmz  ; RECT -0.0600 -0.5200 0.0600 -0.1200 ;
  LAYER vmz  ; RECT -0.0600 0.1200 0.0600 0.5200 ;
  LAYER vmz  ; RECT -0.0600 0.7600 0.0600 1.1600 ;
  LAYER vmz  ; RECT -0.0600 1.4000 0.0600 1.8000 ;
  LAYER gm0  ; RECT -1.2010 -1.9900 1.2010 1.9900 ;
END VMZ_120x400_2401V_3980H_ARRAY_1x6
VIA GV0_800X7400_1080V_2000V
  # gv0   size: x=0.8000 y=7.4000
  # gm0   size: x=1.0800 y=7.6800   enclosure: x=0.1400 y=0.1400
  # gmb   size: x=2.0000 y=8.6000   enclosure: x=0.6000 y=0.6000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5400 -3.8400 0.5400 3.8400 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -1.0000 -4.3000 1.0000 4.3000 ;
END GV0_800X7400_1080V_2000V
VIA GV1_6000X18000_12000V_20000V
  # gv1   size: x=6.0000 y=18.0000
  # gmb   size: x=12.0000 y=24.0000   enclosure: x=3.0000 y=3.0000
  # c4emib   size: x=20.0000 y=20.0000   enclosure: x=7.0000 y=1.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -6.0000 -12.0000 6.0000 12.0000 ;
  LAYER gv1  ; RECT -3.0000 -9.0000 3.0000 9.0000 ;
  LAYER c4emib ; RECT -10.0000 -10.0000 10.0000 10.0000 ;
END GV1_6000X18000_12000V_20000V
VIA GV1_6000X10000_12000V_28000V
  # gv1   size: x=6.0000 y=10.0000
  # gmb   size: x=12.0000 y=16.0000   enclosure: x=3.0000 y=3.0000
  # c4emib   size: x=28.0000 y=28.0000   enclosure: x=11.0000 y=9.0000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -6.0000 -8.0000 6.0000 8.0000 ;
  LAYER gv1  ; RECT -3.0000 -5.0000 3.0000 5.0000 ;
  LAYER c4emib ; RECT -14.0000 -14.0000 14.0000 14.0000 ;
END GV1_6000X10000_12000V_28000V
VIA GV1_6000X30000_12000V_51000V
  # gv1   size: x=6.0000 y=30.0000
  # gmb   size: x=12.0000 y=36.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=51.0000 y=51.0000   enclosure: x=22.5000 y=10.5000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -6.0000 -18.0000 6.0000 18.0000 ;
  LAYER gv1  ; RECT -3.0000 -15.0000 3.0000 15.0000 ;
  LAYER c4   ; RECT -25.5000 -25.5000 25.5000 25.5000 ;
END GV1_6000X30000_12000V_51000V
VIA GV1_6000X30000_12000V_54000V
  # gv1   size: x=6.0000 y=30.0000
  # gmb   size: x=12.0000 y=36.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=54.0000 y=51.0000   enclosure: x=24.0000 y=10.5000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -6.0000 -18.0000 6.0000 18.0000 ;
  LAYER gv1  ; RECT -3.0000 -15.0000 3.0000 15.0000 ;
  LAYER c4   ; RECT -27.0000 -25.5000 27.0000 25.5000 ;
END GV1_6000X30000_12000V_54000V
VIA GV1_6000X30000_12000V_85000V
  # gv1   size: x=6.0000 y=30.0000
  # gmb   size: x=12.0000 y=36.0000   enclosure: x=3.0000 y=3.0000
  # c4   size: x=85.0000 y=51.0000   enclosure: x=39.5000 y=10.5000
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gmb  ; RECT -6.0000 -18.0000 6.0000 18.0000 ;
  LAYER gv1  ; RECT -3.0000 -15.0000 3.0000 15.0000 ;
  LAYER c4   ; RECT -42.5000 -25.5000 42.5000 25.5000 ;
END GV1_6000X30000_12000V_85000V
VIA GV0_800X7400_540V_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.2700 -0.5000 0.2700 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -0.2700 0.5000 0.2700 ;
END GV0_800X7400_540V_1000V_illegal
VIA GV0_800X7400_721V_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.3610 -0.5000 0.3610 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -0.3610 0.5000 0.3610 ;
END GV0_800X7400_721V_1000V_illegal
VIA GV0_800X7400_1080V_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.5400 -0.5000 0.5400 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -0.5400 0.5000 0.5400 ;
END GV0_800X7400_1080V_1000V_illegal
VIA GV0_800X7400_1201V_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.6010 -0.5000 0.6010 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -0.6010 0.5000 0.6010 ;
END GV0_800X7400_1201V_1000V_illegal
VIA GV0_800X7400_2130V_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.0650 -0.5000 1.0650 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -1.0650 0.5000 1.0650 ;
END GV0_800X7400_2130V_1000V_illegal
VIA GV0_800X7400_2401V_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.2010 -0.5000 1.2010 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -1.2010 0.5000 1.2010 ;
END GV0_800X7400_2401V_1000V_illegal
VIA GV0_800X7400_3980V_1000V_illegal
  DEFAULT
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.9900 -0.5000 1.9900 0.5000 ;
  LAYER gv0  ; RECT -0.4000 -3.7000 0.4000 3.7000 ;
  LAYER gmb  ; RECT -0.5000 -1.9900 0.5000 1.9900 ;
END GV0_800X7400_3980V_1000V_illegal


##################################################

VIA via1_108x52S_44H_108V
  # v1   size: x=0.108 y=0.052
  # m1   size: x=0.128 y=0.044   enclosure: x=0.010 y=-0.004
  # m2   size: x=0.108 y=0.096   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.064 -0.022 0.064 0.022 ;
  LAYER v1   ; RECT -0.054 -0.026 0.054 0.026 ;
  LAYER m2   ; RECT -0.054 -0.048 0.054 0.048 ;
END via1_108x52S_44H_108V

VIA via1_108x52S_100H_108V
  # v1   size: x=0.108 y=0.052
  # m1   size: x=0.128 y=0.100   enclosure: x=0.010 y=0.024
  # m2   size: x=0.108 y=0.096   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.064 -0.050 0.064 0.050 ;
  LAYER v1   ; RECT -0.054 -0.026 0.054 0.026 ;
  LAYER m2   ; RECT -0.054 -0.048 0.054 0.048 ;
END via1_108x52S_100H_108V

VIA via1_108x60S_100H_108V
  # v1   size: x=0.108 y=0.060
  # m1   size: x=0.128 y=0.100   enclosure: x=0.010 y=0.020
  # m2   size: x=0.108 y=0.104   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.064 -0.050 0.064 0.050 ;
  LAYER v1   ; RECT -0.054 -0.030 0.054 0.030 ;
  LAYER m2   ; RECT -0.054 -0.052 0.054 0.052 ;
END via1_108x60S_100H_108V

VIA via1_60Sx44_44H_44H
  # v1   size: x=0.060 y=0.044
  # m1   size: x=0.068 y=0.044   enclosure: x=0.004 y=0.000
  # m2   size: x=0.104 y=0.044   enclosure: x=0.022 y=0.000
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.034 -0.022 0.034 0.022 ;
  LAYER v1   ; RECT -0.030 -0.022 0.030 0.022 ;
  LAYER m2   ; RECT -0.052 -0.022 0.052 0.022 ;
END via1_60Sx44_44H_44H

VIA via1_60Sx44_100H_44H
  # v1   size: x=0.060 y=0.044
  # m1   size: x=0.080 y=0.100   enclosure: x=0.010 y=0.028
  # m2   size: x=0.104 y=0.044   enclosure: x=0.022 y=0.000
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.040 -0.050 0.040 0.050 ;
  LAYER v1   ; RECT -0.030 -0.022 0.030 0.022 ;
  LAYER m2   ; RECT -0.052 -0.022 0.052 0.022 ;
END via1_60Sx44_100H_44H

VIA via1_60Sx56_100H_56H
  # v1   size: x=0.060 y=0.056
  # m1   size: x=0.080 y=0.100   enclosure: x=0.010 y=0.022
  # m2   size: x=0.104 y=0.056   enclosure: x=0.022 y=0.000
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.040 -0.050 0.040 0.050 ;
  LAYER v1   ; RECT -0.030 -0.028 0.030 0.028 ;
  LAYER m2   ; RECT -0.052 -0.028 0.052 0.028 ;
END via1_60Sx56_100H_56H

VIA via1_60Sx76_100H_76H
  # v1   size: x=0.060 y=0.076
  # m1   size: x=0.080 y=0.100   enclosure: x=0.010 y=0.012
  # m2   size: x=0.104 y=0.076   enclosure: x=0.022 y=0.000
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.040 -0.050 0.040 0.050 ;
  LAYER v1   ; RECT -0.030 -0.038 0.030 0.038 ;
  LAYER m2   ; RECT -0.052 -0.038 0.052 0.038 ;
END via1_60Sx76_100H_76H

VIA via1_60Sx90_100H_90H
  # v1   size: x=0.060 y=0.090
  # m1   size: x=0.080 y=0.100   enclosure: x=0.010 y=0.005
  # m2   size: x=0.104 y=0.090   enclosure: x=0.022 y=0.000
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.040 -0.050 0.040 0.050 ;
  LAYER v1   ; RECT -0.030 -0.045 0.030 0.045 ;
  LAYER m2   ; RECT -0.052 -0.045 0.052 0.045 ;
END via1_60Sx90_100H_90H

VIA via1_70x70_100V_90H
  # v1   size: x=0.070 y=0.070
  # m1   size: x=0.100 y=0.090   enclosure: x=0.015 y=0.010
  # m2   size: x=0.114 y=0.090   enclosure: x=0.022 y=0.010
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.050 -0.045 0.050 0.045 ;
  LAYER v1   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m2   ; RECT -0.057 -0.045 0.057 0.045 ;
END via1_70x70_100V_90H

VIA via1_70x70_100V_108H
  # v1   size: x=0.070 y=0.070
  # m1   size: x=0.100 y=0.090   enclosure: x=0.015 y=0.010
  # m2   size: x=0.114 y=0.108   enclosure: x=0.022 y=0.019
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.050 -0.045 0.050 0.045 ;
  LAYER v1   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m2   ; RECT -0.057 -0.054 0.057 0.054 ;
END via1_70x70_100V_108H

VIA via1_70x70_100V_90V
  # v1   size: x=0.070 y=0.070
  # m1   size: x=0.100 y=0.090   enclosure: x=0.015 y=0.010
  # m2   size: x=0.090 y=0.114   enclosure: x=0.010 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.050 -0.045 0.050 0.045 ;
  LAYER v1   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m2   ; RECT -0.045 -0.057 0.045 0.057 ;
END via1_70x70_100V_90V

VIA via1_70x70_100V_108V
  # v1   size: x=0.070 y=0.070
  # m1   size: x=0.100 y=0.090   enclosure: x=0.015 y=0.010
  # m2   size: x=0.108 y=0.114   enclosure: x=0.019 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.050 -0.045 0.050 0.045 ;
  LAYER v1   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m2   ; RECT -0.054 -0.057 0.054 0.057 ;
END via1_70x70_100V_108V

VIA via1_70x70_100H_90H
  # v1   size: x=0.070 y=0.070
  # m1   size: x=0.090 y=0.100   enclosure: x=0.010 y=0.015
  # m2   size: x=0.114 y=0.090   enclosure: x=0.022 y=0.010
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.045 -0.050 0.045 0.050 ;
  LAYER v1   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m2   ; RECT -0.057 -0.045 0.057 0.045 ;
END via1_70x70_100H_90H

VIA via1_70x70_100H_108H
  # v1   size: x=0.070 y=0.070
  # m1   size: x=0.090 y=0.100   enclosure: x=0.010 y=0.015
  # m2   size: x=0.114 y=0.108   enclosure: x=0.022 y=0.019
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.045 -0.050 0.045 0.050 ;
  LAYER v1   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m2   ; RECT -0.057 -0.054 0.057 0.054 ;
END via1_70x70_100H_108H

VIA via1_70x70_100H_90V
  # v1   size: x=0.070 y=0.070
  # m1   size: x=0.090 y=0.100   enclosure: x=0.010 y=0.015
  # m2   size: x=0.090 y=0.114   enclosure: x=0.010 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.045 -0.050 0.045 0.050 ;
  LAYER v1   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m2   ; RECT -0.045 -0.057 0.045 0.057 ;
END via1_70x70_100H_90V

VIA via1_70x70_100H_108V
  # v1   size: x=0.070 y=0.070
  # m1   size: x=0.090 y=0.100   enclosure: x=0.010 y=0.015
  # m2   size: x=0.108 y=0.114   enclosure: x=0.019 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.045 -0.050 0.045 0.050 ;
  LAYER v1   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m2   ; RECT -0.054 -0.057 0.054 0.057 ;
END via1_70x70_100H_108V

VIA via1_76x52S_44H_76V
  # v1   size: x=0.076 y=0.052
  # m1   size: x=0.096 y=0.044   enclosure: x=0.010 y=-0.004
  # m2   size: x=0.076 y=0.096   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.048 -0.022 0.048 0.022 ;
  LAYER v1   ; RECT -0.038 -0.026 0.038 0.026 ;
  LAYER m2   ; RECT -0.038 -0.048 0.038 0.048 ;
END via1_76x52S_44H_76V

VIA via1_76x52S_100H_76V
  # v1   size: x=0.076 y=0.052
  # m1   size: x=0.096 y=0.100   enclosure: x=0.010 y=0.024
  # m2   size: x=0.076 y=0.096   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.048 -0.050 0.048 0.050 ;
  LAYER v1   ; RECT -0.038 -0.026 0.038 0.026 ;
  LAYER m2   ; RECT -0.038 -0.048 0.038 0.048 ;
END via1_76x52S_100H_76V

VIA via1_76x52S_100V_76V
  # v1   size: x=0.076 y=0.052
  # m1   size: x=0.100 y=0.072   enclosure: x=0.012 y=0.010
  # m2   size: x=0.076 y=0.096   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.050 -0.036 0.050 0.036 ;
  LAYER v1   ; RECT -0.038 -0.026 0.038 0.026 ;
  LAYER m2   ; RECT -0.038 -0.048 0.038 0.048 ;
END via1_76x52S_100V_76V

VIA via1_76x60S_100V_76V
  # v1   size: x=0.076 y=0.060
  # m1   size: x=0.100 y=0.080   enclosure: x=0.012 y=0.010
  # m2   size: x=0.076 y=0.104   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.050 -0.040 0.050 0.040 ;
  LAYER v1   ; RECT -0.038 -0.030 0.038 0.030 ;
  LAYER m2   ; RECT -0.038 -0.052 0.038 0.052 ;
END via1_76x60S_100V_76V

VIA via1_76x60S_100H_76V
  # v1   size: x=0.076 y=0.060
  # m1   size: x=0.096 y=0.100   enclosure: x=0.010 y=0.020
  # m2   size: x=0.076 y=0.104   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.048 -0.050 0.048 0.050 ;
  LAYER v1   ; RECT -0.038 -0.030 0.038 0.030 ;
  LAYER m2   ; RECT -0.038 -0.052 0.038 0.052 ;
END via1_76x60S_100H_76V

VIA via1_90x52S_44H_90V
  # v1   size: x=0.090 y=0.052
  # m1   size: x=0.110 y=0.044   enclosure: x=0.010 y=-0.004
  # m2   size: x=0.090 y=0.096   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.055 -0.022 0.055 0.022 ;
  LAYER v1   ; RECT -0.045 -0.026 0.045 0.026 ;
  LAYER m2   ; RECT -0.045 -0.048 0.045 0.048 ;
END via1_90x52S_44H_90V

VIA via1_90x52S_100H_90V
  # v1   size: x=0.090 y=0.052
  # m1   size: x=0.110 y=0.100   enclosure: x=0.010 y=0.024
  # m2   size: x=0.090 y=0.096   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.055 -0.050 0.055 0.050 ;
  LAYER v1   ; RECT -0.045 -0.026 0.045 0.026 ;
  LAYER m2   ; RECT -0.045 -0.048 0.045 0.048 ;
END via1_90x52S_100H_90V

VIA via1_90x52S_100V_90V
  # v1   size: x=0.090 y=0.052
  # m1   size: x=0.100 y=0.072   enclosure: x=0.005 y=0.010
  # m2   size: x=0.090 y=0.096   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.050 -0.036 0.050 0.036 ;
  LAYER v1   ; RECT -0.045 -0.026 0.045 0.026 ;
  LAYER m2   ; RECT -0.045 -0.048 0.045 0.048 ;
END via1_90x52S_100V_90V

VIA via1_90x60S_44H_90V
  # v1   size: x=0.090 y=0.060
  # m1   size: x=0.110 y=0.044   enclosure: x=0.010 y=-0.008
  # m2   size: x=0.090 y=0.104   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.055 -0.022 0.055 0.022 ;
  LAYER v1   ; RECT -0.045 -0.030 0.045 0.030 ;
  LAYER m2   ; RECT -0.045 -0.052 0.045 0.052 ;
END via1_90x60S_44H_90V

VIA via1_90x60S_100H_90V
  # v1   size: x=0.090 y=0.060
  # m1   size: x=0.110 y=0.100   enclosure: x=0.010 y=0.020
  # m2   size: x=0.090 y=0.104   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.055 -0.050 0.055 0.050 ;
  LAYER v1   ; RECT -0.045 -0.030 0.045 0.030 ;
  LAYER m2   ; RECT -0.045 -0.052 0.045 0.052 ;
END via1_90x60S_100H_90V

VIA via1_90x60S_100V_90V
  # v1   size: x=0.090 y=0.060
  # m1   size: x=0.100 y=0.080   enclosure: x=0.005 y=0.010
  # m2   size: x=0.090 y=0.104   enclosure: x=0.000 y=0.022
  RESISTANCE 1.000 ;
  LAYER m1   ; RECT -0.050 -0.040 0.050 0.040 ;
  LAYER v1   ; RECT -0.045 -0.030 0.045 0.030 ;
  LAYER m2   ; RECT -0.045 -0.052 0.045 0.052 ;
END via1_90x60S_100V_90V

VIA via2_44x58S_76V_44V
  # v2   size: x=0.044 y=0.058
  # m2   size: x=0.076 y=0.082   enclosure: x=0.016 y=0.012
  # m3   size: x=0.044 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.038 -0.041 0.038 0.041 ;
  LAYER v2   ; RECT -0.022 -0.029 0.022 0.029 ;
  LAYER m3   ; RECT -0.022 -0.050 0.022 0.050 ;
END via2_44x58S_76V_44V

VIA via2_44x58S_90V_44V
  # v2   size: x=0.044 y=0.058
  # m2   size: x=0.090 y=0.082   enclosure: x=0.023 y=0.012
  # m3   size: x=0.044 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.045 -0.041 0.045 0.041 ;
  LAYER v2   ; RECT -0.022 -0.029 0.022 0.029 ;
  LAYER m3   ; RECT -0.022 -0.050 0.022 0.050 ;
END via2_44x58S_90V_44V

VIA via2_44x58S_108V_44V
  # v2   size: x=0.044 y=0.058
  # m2   size: x=0.108 y=0.082   enclosure: x=0.032 y=0.012
  # m3   size: x=0.044 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v2   ; RECT -0.022 -0.029 0.022 0.029 ;
  LAYER m3   ; RECT -0.022 -0.050 0.022 0.050 ;
END via2_44x58S_108V_44V

VIA via2_56x58S_76V_56V
  # v2   size: x=0.056 y=0.058
  # m2   size: x=0.076 y=0.082   enclosure: x=0.010 y=0.012
  # m3   size: x=0.056 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.038 -0.041 0.038 0.041 ;
  LAYER v2   ; RECT -0.028 -0.029 0.028 0.029 ;
  LAYER m3   ; RECT -0.028 -0.050 0.028 0.050 ;
END via2_56x58S_76V_56V

VIA via2_56x58S_90V_56V
  # v2   size: x=0.056 y=0.058
  # m2   size: x=0.090 y=0.082   enclosure: x=0.017 y=0.012
  # m3   size: x=0.056 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.045 -0.041 0.045 0.041 ;
  LAYER v2   ; RECT -0.028 -0.029 0.028 0.029 ;
  LAYER m3   ; RECT -0.028 -0.050 0.028 0.050 ;
END via2_56x58S_90V_56V

VIA via2_56x58S_108V_56V
  # v2   size: x=0.056 y=0.058
  # m2   size: x=0.108 y=0.082   enclosure: x=0.026 y=0.012
  # m3   size: x=0.056 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v2   ; RECT -0.028 -0.029 0.028 0.029 ;
  LAYER m3   ; RECT -0.028 -0.050 0.028 0.050 ;
END via2_56x58S_108V_56V

VIA via2_58Sx108_76V_108H
  # v2   size: x=0.058 y=0.108
  # m2   size: x=0.076 y=0.132   enclosure: x=0.009 y=0.012
  # m3   size: x=0.100 y=0.108   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.038 -0.066 0.038 0.066 ;
  LAYER v2   ; RECT -0.029 -0.054 0.029 0.054 ;
  LAYER m3   ; RECT -0.050 -0.054 0.050 0.054 ;
END via2_58Sx108_76V_108H

VIA via2_58Sx108_90V_108H
  # v2   size: x=0.058 y=0.108
  # m2   size: x=0.090 y=0.132   enclosure: x=0.016 y=0.012
  # m3   size: x=0.100 y=0.108   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.045 -0.066 0.045 0.066 ;
  LAYER v2   ; RECT -0.029 -0.054 0.029 0.054 ;
  LAYER m3   ; RECT -0.050 -0.054 0.050 0.054 ;
END via2_58Sx108_90V_108H

VIA via2_58Sx108_108V_108H
  # v2   size: x=0.058 y=0.108
  # m2   size: x=0.108 y=0.132   enclosure: x=0.025 y=0.012
  # m3   size: x=0.100 y=0.108   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.054 -0.066 0.054 0.066 ;
  LAYER v2   ; RECT -0.029 -0.054 0.029 0.054 ;
  LAYER m3   ; RECT -0.050 -0.054 0.050 0.054 ;
END via2_58Sx108_108V_108H

VIA via2_58Sx76_76H_76H
  # v2   size: x=0.058 y=0.076
  # m2   size: x=0.082 y=0.076   enclosure: x=0.012 y=0.000
  # m3   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.041 -0.038 0.041 0.038 ;
  LAYER v2   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m3   ; RECT -0.050 -0.038 0.050 0.038 ;
END via2_58Sx76_76H_76H

VIA via2_58Sx76_90H_76H
  # v2   size: x=0.058 y=0.076
  # m2   size: x=0.082 y=0.090   enclosure: x=0.012 y=0.007
  # m3   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.041 -0.045 0.041 0.045 ;
  LAYER v2   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m3   ; RECT -0.050 -0.038 0.050 0.038 ;
END via2_58Sx76_90H_76H

VIA via2_58Sx76_108H_76H
  # v2   size: x=0.058 y=0.076
  # m2   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.016
  # m3   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v2   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m3   ; RECT -0.050 -0.038 0.050 0.038 ;
END via2_58Sx76_108H_76H

VIA via2_58Sx76_76V_76H
  # v2   size: x=0.058 y=0.076
  # m2   size: x=0.076 y=0.100   enclosure: x=0.009 y=0.012
  # m3   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.038 -0.050 0.038 0.050 ;
  LAYER v2   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m3   ; RECT -0.050 -0.038 0.050 0.038 ;
END via2_58Sx76_76V_76H

VIA via2_58Sx76_90V_76H
  # v2   size: x=0.058 y=0.076
  # m2   size: x=0.090 y=0.100   enclosure: x=0.016 y=0.012
  # m3   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.045 -0.050 0.045 0.050 ;
  LAYER v2   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m3   ; RECT -0.050 -0.038 0.050 0.038 ;
END via2_58Sx76_90V_76H

VIA via2_58Sx76_108V_76H
  # v2   size: x=0.058 y=0.076
  # m2   size: x=0.108 y=0.100   enclosure: x=0.025 y=0.012
  # m3   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.054 -0.050 0.054 0.050 ;
  LAYER v2   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m3   ; RECT -0.050 -0.038 0.050 0.038 ;
END via2_58Sx76_108V_76H

VIA via2_58Sx90_76V_90H
  # v2   size: x=0.058 y=0.090
  # m2   size: x=0.076 y=0.114   enclosure: x=0.009 y=0.012
  # m3   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.038 -0.057 0.038 0.057 ;
  LAYER v2   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m3   ; RECT -0.050 -0.045 0.050 0.045 ;
END via2_58Sx90_76V_90H

VIA via2_58Sx90_90V_90H
  # v2   size: x=0.058 y=0.090
  # m2   size: x=0.090 y=0.114   enclosure: x=0.016 y=0.012
  # m3   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.045 -0.057 0.045 0.057 ;
  LAYER v2   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m3   ; RECT -0.050 -0.045 0.050 0.045 ;
END via2_58Sx90_90V_90H

VIA via2_58Sx90_108V_90H
  # v2   size: x=0.058 y=0.090
  # m2   size: x=0.108 y=0.114   enclosure: x=0.025 y=0.012
  # m3   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.054 -0.057 0.054 0.057 ;
  LAYER v2   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m3   ; RECT -0.050 -0.045 0.050 0.045 ;
END via2_58Sx90_108V_90H

VIA via2_58Sx90_108H_90H
  # v2   size: x=0.058 y=0.090
  # m2   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.009
  # m3   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v2   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m3   ; RECT -0.050 -0.045 0.050 0.045 ;
END via2_58Sx90_108H_90H

VIA via2_70x70_56H_90V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.056   enclosure: x=0.012 y=-0.007
  # m3   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.028 0.047 0.028 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.045 -0.056 0.045 0.056 ;
END via2_70x70_56H_90V

VIA via2_70x70_56H_108V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.056   enclosure: x=0.012 y=-0.007
  # m3   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.028 0.047 0.028 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.054 -0.056 0.054 0.056 ;
END via2_70x70_56H_108V

VIA via2_70x70_76H_90V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m3   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.045 -0.056 0.045 0.056 ;
END via2_70x70_76H_90V

VIA via2_70x70_76H_108V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m3   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.054 -0.056 0.054 0.056 ;
END via2_70x70_76H_108V

VIA via2_70x70_90H_90V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m3   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.045 -0.056 0.045 0.056 ;
END via2_70x70_90H_90V

VIA via2_70x70_90H_108V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m3   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.054 -0.056 0.054 0.056 ;
END via2_70x70_90H_108V

VIA via2_70x70_108H_90V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m3   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.045 -0.056 0.045 0.056 ;
END via2_70x70_108H_90V

VIA via2_70x70_108H_108V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m3   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.054 -0.056 0.054 0.056 ;
END via2_70x70_108H_108V

VIA via2_70x70_76V_90V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m3   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.045 -0.056 0.045 0.056 ;
END via2_70x70_76V_90V

VIA via2_70x70_76V_108V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m3   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.054 -0.056 0.054 0.056 ;
END via2_70x70_76V_108V

VIA via2_70x70_76V_90H
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m3   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.056 -0.045 0.056 0.045 ;
END via2_70x70_76V_90H

VIA via2_70x70_76V_108H
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m3   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.056 -0.054 0.056 0.054 ;
END via2_70x70_76V_108H

VIA via2_70x70_90V_90V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m3   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.045 -0.056 0.045 0.056 ;
END via2_70x70_90V_90V

VIA via2_70x70_90V_108V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m3   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.054 -0.056 0.054 0.056 ;
END via2_70x70_90V_108V

VIA via2_70x70_90V_90H
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m3   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.056 -0.045 0.056 0.045 ;
END via2_70x70_90V_90H

VIA via2_70x70_90V_108H
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m3   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.056 -0.054 0.056 0.054 ;
END via2_70x70_90V_108H

VIA via2_70x70_108V_90V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m3   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.045 -0.056 0.045 0.056 ;
END via2_70x70_108V_90V

VIA via2_70x70_108V_108V
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m3   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.054 -0.056 0.054 0.056 ;
END via2_70x70_108V_108V

VIA via2_70x70_108V_90H
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m3   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.056 -0.045 0.056 0.045 ;
END via2_70x70_108V_90H

VIA via2_70x70_108V_108H
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m3   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.056 -0.054 0.056 0.054 ;
END via2_70x70_108V_108H

VIA via2_70x70_90H_90H
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m3   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.056 -0.045 0.056 0.045 ;
END via2_70x70_90H_90H

VIA via2_70x70_90H_108H
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m3   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.056 -0.054 0.056 0.054 ;
END via2_70x70_90H_108H

VIA via2_70x70_108H_90H
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m3   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.056 -0.045 0.056 0.045 ;
END via2_70x70_108H_90H

VIA via2_70x70_108H_108H
  # v2   size: x=0.070 y=0.070
  # m2   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m3   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v2   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m3   ; RECT -0.056 -0.054 0.056 0.054 ;
END via2_70x70_108H_108H

VIA via2_76x58S_76V_76V
  # v2   size: x=0.076 y=0.058
  # m2   size: x=0.076 y=0.082   enclosure: x=0.000 y=0.012
  # m3   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.038 -0.041 0.038 0.041 ;
  LAYER v2   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m3   ; RECT -0.038 -0.050 0.038 0.050 ;
END via2_76x58S_76V_76V

VIA via2_76x58S_90V_76V
  # v2   size: x=0.076 y=0.058
  # m2   size: x=0.090 y=0.082   enclosure: x=0.007 y=0.012
  # m3   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.045 -0.041 0.045 0.041 ;
  LAYER v2   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m3   ; RECT -0.038 -0.050 0.038 0.050 ;
END via2_76x58S_90V_76V

VIA via2_76x58S_108V_76V
  # v2   size: x=0.076 y=0.058
  # m2   size: x=0.108 y=0.082   enclosure: x=0.016 y=0.012
  # m3   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v2   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m3   ; RECT -0.038 -0.050 0.038 0.050 ;
END via2_76x58S_108V_76V

VIA via2_90x58S_108V_90V
  # v2   size: x=0.090 y=0.058
  # m2   size: x=0.108 y=0.082   enclosure: x=0.009 y=0.012
  # m3   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m2   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v2   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m3   ; RECT -0.045 -0.050 0.045 0.050 ;
END via2_90x58S_108V_90V

VIA via3_108x58S_76H_108V
  # v3   size: x=0.108 y=0.058
  # m3   size: x=0.132 y=0.076   enclosure: x=0.012 y=0.009
  # m4   size: x=0.108 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.066 -0.038 0.066 0.038 ;
  LAYER v3   ; RECT -0.054 -0.029 0.054 0.029 ;
  LAYER m4   ; RECT -0.054 -0.050 0.054 0.050 ;
END via3_108x58S_76H_108V

VIA via3_108x58S_90H_108V
  # v3   size: x=0.108 y=0.058
  # m3   size: x=0.132 y=0.090   enclosure: x=0.012 y=0.016
  # m4   size: x=0.108 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.066 -0.045 0.066 0.045 ;
  LAYER v3   ; RECT -0.054 -0.029 0.054 0.029 ;
  LAYER m4   ; RECT -0.054 -0.050 0.054 0.050 ;
END via3_108x58S_90H_108V

VIA via3_108x58S_108H_108V
  # v3   size: x=0.108 y=0.058
  # m3   size: x=0.132 y=0.108   enclosure: x=0.012 y=0.025
  # m4   size: x=0.108 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.066 -0.054 0.066 0.054 ;
  LAYER v3   ; RECT -0.054 -0.029 0.054 0.029 ;
  LAYER m4   ; RECT -0.054 -0.050 0.054 0.050 ;
END via3_108x58S_108H_108V

VIA via3_58Sx44_76H_44H
  # v3   size: x=0.058 y=0.044
  # m3   size: x=0.082 y=0.076   enclosure: x=0.012 y=0.016
  # m4   size: x=0.100 y=0.044   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.041 -0.038 0.041 0.038 ;
  LAYER v3   ; RECT -0.029 -0.022 0.029 0.022 ;
  LAYER m4   ; RECT -0.050 -0.022 0.050 0.022 ;
END via3_58Sx44_76H_44H

VIA via3_58Sx44_90H_44H
  # v3   size: x=0.058 y=0.044
  # m3   size: x=0.082 y=0.090   enclosure: x=0.012 y=0.023
  # m4   size: x=0.100 y=0.044   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.041 -0.045 0.041 0.045 ;
  LAYER v3   ; RECT -0.029 -0.022 0.029 0.022 ;
  LAYER m4   ; RECT -0.050 -0.022 0.050 0.022 ;
END via3_58Sx44_90H_44H

VIA via3_58Sx44_108H_44H
  # v3   size: x=0.058 y=0.044
  # m3   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.032
  # m4   size: x=0.100 y=0.044   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v3   ; RECT -0.029 -0.022 0.029 0.022 ;
  LAYER m4   ; RECT -0.050 -0.022 0.050 0.022 ;
END via3_58Sx44_108H_44H

VIA via3_58Sx56_76H_56H
  # v3   size: x=0.058 y=0.056
  # m3   size: x=0.082 y=0.076   enclosure: x=0.012 y=0.010
  # m4   size: x=0.100 y=0.056   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.041 -0.038 0.041 0.038 ;
  LAYER v3   ; RECT -0.029 -0.028 0.029 0.028 ;
  LAYER m4   ; RECT -0.050 -0.028 0.050 0.028 ;
END via3_58Sx56_76H_56H

VIA via3_58Sx56_90H_56H
  # v3   size: x=0.058 y=0.056
  # m3   size: x=0.082 y=0.090   enclosure: x=0.012 y=0.017
  # m4   size: x=0.100 y=0.056   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.041 -0.045 0.041 0.045 ;
  LAYER v3   ; RECT -0.029 -0.028 0.029 0.028 ;
  LAYER m4   ; RECT -0.050 -0.028 0.050 0.028 ;
END via3_58Sx56_90H_56H

VIA via3_58Sx56_108H_56H
  # v3   size: x=0.058 y=0.056
  # m3   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.026
  # m4   size: x=0.100 y=0.056   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v3   ; RECT -0.029 -0.028 0.029 0.028 ;
  LAYER m4   ; RECT -0.050 -0.028 0.050 0.028 ;
END via3_58Sx56_108H_56H

VIA via3_58Sx76_76H_76H
  # v3   size: x=0.058 y=0.076
  # m3   size: x=0.082 y=0.076   enclosure: x=0.012 y=0.000
  # m4   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.041 -0.038 0.041 0.038 ;
  LAYER v3   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m4   ; RECT -0.050 -0.038 0.050 0.038 ;
END via3_58Sx76_76H_76H

VIA via3_58Sx76_90H_76H
  # v3   size: x=0.058 y=0.076
  # m3   size: x=0.082 y=0.090   enclosure: x=0.012 y=0.007
  # m4   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.041 -0.045 0.041 0.045 ;
  LAYER v3   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m4   ; RECT -0.050 -0.038 0.050 0.038 ;
END via3_58Sx76_90H_76H

VIA via3_58Sx76_108H_76H
  # v3   size: x=0.058 y=0.076
  # m3   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.016
  # m4   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v3   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m4   ; RECT -0.050 -0.038 0.050 0.038 ;
END via3_58Sx76_108H_76H

VIA via3_58Sx90_108H_90H
  # v3   size: x=0.058 y=0.090
  # m3   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.009
  # m4   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v3   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m4   ; RECT -0.050 -0.045 0.050 0.045 ;
END via3_58Sx90_108H_90H

VIA via3_70x70_56V_90H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.056 y=0.094   enclosure: x=-0.007 y=0.012
  # m4   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.028 -0.047 0.028 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.045 0.056 0.045 ;
END via3_70x70_56V_90H

VIA via3_70x70_56V_108H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.056 y=0.094   enclosure: x=-0.007 y=0.012
  # m4   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.028 -0.047 0.028 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.054 0.056 0.054 ;
END via3_70x70_56V_108H

VIA via3_70x70_76V_90H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m4   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.045 0.056 0.045 ;
END via3_70x70_76V_90H

VIA via3_70x70_76V_108H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m4   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.054 0.056 0.054 ;
END via3_70x70_76V_108H

VIA via3_70x70_90V_90H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m4   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.045 0.056 0.045 ;
END via3_70x70_90V_90H

VIA via3_70x70_90V_108H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m4   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.054 0.056 0.054 ;
END via3_70x70_90V_108H

VIA via3_70x70_108V_90H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m4   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.045 0.056 0.045 ;
END via3_70x70_108V_90H

VIA via3_70x70_108V_108H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m4   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.054 0.056 0.054 ;
END via3_70x70_108V_108H

VIA via3_70x70_76H_90H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m4   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.045 0.056 0.045 ;
END via3_70x70_76H_90H

VIA via3_70x70_76H_108H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m4   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.054 0.056 0.054 ;
END via3_70x70_76H_108H

VIA via3_70x70_76H_90V
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m4   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.045 -0.056 0.045 0.056 ;
END via3_70x70_76H_90V

VIA via3_70x70_76H_108V
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m4   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.054 -0.056 0.054 0.056 ;
END via3_70x70_76H_108V

VIA via3_70x70_90H_90H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m4   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.045 0.056 0.045 ;
END via3_70x70_90H_90H

VIA via3_70x70_90H_108H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m4   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.054 0.056 0.054 ;
END via3_70x70_90H_108H

VIA via3_70x70_90H_90V
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m4   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.045 -0.056 0.045 0.056 ;
END via3_70x70_90H_90V

VIA via3_70x70_90H_108V
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m4   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.054 -0.056 0.054 0.056 ;
END via3_70x70_90H_108V

VIA via3_70x70_108H_90H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m4   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.045 0.056 0.045 ;
END via3_70x70_108H_90H

VIA via3_70x70_108H_108H
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m4   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.056 -0.054 0.056 0.054 ;
END via3_70x70_108H_108H

VIA via3_70x70_108H_90V
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m4   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.045 -0.056 0.045 0.056 ;
END via3_70x70_108H_90V

VIA via3_70x70_108H_108V
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m4   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.054 -0.056 0.054 0.056 ;
END via3_70x70_108H_108V

VIA via3_70x70_90V_90V
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m4   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.045 -0.056 0.045 0.056 ;
END via3_70x70_90V_90V

VIA via3_70x70_90V_108V
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m4   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.054 -0.056 0.054 0.056 ;
END via3_70x70_90V_108V

VIA via3_70x70_108V_90V
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m4   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.045 -0.056 0.045 0.056 ;
END via3_70x70_108V_90V

VIA via3_70x70_108V_108V
  # v3   size: x=0.070 y=0.070
  # m3   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m4   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v3   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m4   ; RECT -0.054 -0.056 0.054 0.056 ;
END via3_70x70_108V_108V

VIA via3_76x58S_76V_76V
  # v3   size: x=0.076 y=0.058
  # m3   size: x=0.076 y=0.082   enclosure: x=0.000 y=0.012
  # m4   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.038 -0.041 0.038 0.041 ;
  LAYER v3   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m4   ; RECT -0.038 -0.050 0.038 0.050 ;
END via3_76x58S_76V_76V

VIA via3_76x58S_90V_76V
  # v3   size: x=0.076 y=0.058
  # m3   size: x=0.090 y=0.082   enclosure: x=0.007 y=0.012
  # m4   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.045 -0.041 0.045 0.041 ;
  LAYER v3   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m4   ; RECT -0.038 -0.050 0.038 0.050 ;
END via3_76x58S_90V_76V

VIA via3_76x58S_108V_76V
  # v3   size: x=0.076 y=0.058
  # m3   size: x=0.108 y=0.082   enclosure: x=0.016 y=0.012
  # m4   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v3   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m4   ; RECT -0.038 -0.050 0.038 0.050 ;
END via3_76x58S_108V_76V

VIA via3_76x58S_76H_76V
  # v3   size: x=0.076 y=0.058
  # m3   size: x=0.100 y=0.076   enclosure: x=0.012 y=0.009
  # m4   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.050 -0.038 0.050 0.038 ;
  LAYER v3   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m4   ; RECT -0.038 -0.050 0.038 0.050 ;
END via3_76x58S_76H_76V

VIA via3_76x58S_90H_76V
  # v3   size: x=0.076 y=0.058
  # m3   size: x=0.100 y=0.090   enclosure: x=0.012 y=0.016
  # m4   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.050 -0.045 0.050 0.045 ;
  LAYER v3   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m4   ; RECT -0.038 -0.050 0.038 0.050 ;
END via3_76x58S_90H_76V

VIA via3_76x58S_108H_76V
  # v3   size: x=0.076 y=0.058
  # m3   size: x=0.100 y=0.108   enclosure: x=0.012 y=0.025
  # m4   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.050 -0.054 0.050 0.054 ;
  LAYER v3   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m4   ; RECT -0.038 -0.050 0.038 0.050 ;
END via3_76x58S_108H_76V

VIA via3_90x58S_76H_90V
  # v3   size: x=0.090 y=0.058
  # m3   size: x=0.114 y=0.076   enclosure: x=0.012 y=0.009
  # m4   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.057 -0.038 0.057 0.038 ;
  LAYER v3   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m4   ; RECT -0.045 -0.050 0.045 0.050 ;
END via3_90x58S_76H_90V

VIA via3_90x58S_90H_90V
  # v3   size: x=0.090 y=0.058
  # m3   size: x=0.114 y=0.090   enclosure: x=0.012 y=0.016
  # m4   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.057 -0.045 0.057 0.045 ;
  LAYER v3   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m4   ; RECT -0.045 -0.050 0.045 0.050 ;
END via3_90x58S_90H_90V

VIA via3_90x58S_108H_90V
  # v3   size: x=0.090 y=0.058
  # m3   size: x=0.114 y=0.108   enclosure: x=0.012 y=0.025
  # m4   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.057 -0.054 0.057 0.054 ;
  LAYER v3   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m4   ; RECT -0.045 -0.050 0.045 0.050 ;
END via3_90x58S_108H_90V

VIA via3_90x58S_108V_90V
  # v3   size: x=0.090 y=0.058
  # m3   size: x=0.108 y=0.082   enclosure: x=0.009 y=0.012
  # m4   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m3   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v3   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m4   ; RECT -0.045 -0.050 0.045 0.050 ;
END via3_90x58S_108V_90V

VIA via4_44x58S_76V_44V
  # v4   size: x=0.044 y=0.058
  # m4   size: x=0.076 y=0.082   enclosure: x=0.016 y=0.012
  # m5   size: x=0.044 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.041 0.038 0.041 ;
  LAYER v4   ; RECT -0.022 -0.029 0.022 0.029 ;
  LAYER m5   ; RECT -0.022 -0.050 0.022 0.050 ;
END via4_44x58S_76V_44V

VIA via4_44x58S_90V_44V
  # v4   size: x=0.044 y=0.058
  # m4   size: x=0.090 y=0.082   enclosure: x=0.023 y=0.012
  # m5   size: x=0.044 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.041 0.045 0.041 ;
  LAYER v4   ; RECT -0.022 -0.029 0.022 0.029 ;
  LAYER m5   ; RECT -0.022 -0.050 0.022 0.050 ;
END via4_44x58S_90V_44V

VIA via4_44x58S_108V_44V
  # v4   size: x=0.044 y=0.058
  # m4   size: x=0.108 y=0.082   enclosure: x=0.032 y=0.012
  # m5   size: x=0.044 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v4   ; RECT -0.022 -0.029 0.022 0.029 ;
  LAYER m5   ; RECT -0.022 -0.050 0.022 0.050 ;
END via4_44x58S_108V_44V

VIA via4_56x58S_76V_56V
  # v4   size: x=0.056 y=0.058
  # m4   size: x=0.076 y=0.082   enclosure: x=0.010 y=0.012
  # m5   size: x=0.056 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.041 0.038 0.041 ;
  LAYER v4   ; RECT -0.028 -0.029 0.028 0.029 ;
  LAYER m5   ; RECT -0.028 -0.050 0.028 0.050 ;
END via4_56x58S_76V_56V

VIA via4_56x58S_90V_56V
  # v4   size: x=0.056 y=0.058
  # m4   size: x=0.090 y=0.082   enclosure: x=0.017 y=0.012
  # m5   size: x=0.056 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.041 0.045 0.041 ;
  LAYER v4   ; RECT -0.028 -0.029 0.028 0.029 ;
  LAYER m5   ; RECT -0.028 -0.050 0.028 0.050 ;
END via4_56x58S_90V_56V

VIA via4_56x58S_108V_56V
  # v4   size: x=0.056 y=0.058
  # m4   size: x=0.108 y=0.082   enclosure: x=0.026 y=0.012
  # m5   size: x=0.056 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v4   ; RECT -0.028 -0.029 0.028 0.029 ;
  LAYER m5   ; RECT -0.028 -0.050 0.028 0.050 ;
END via4_56x58S_108V_56V

VIA via4_58Sx108_76V_108H
  # v4   size: x=0.058 y=0.108
  # m4   size: x=0.076 y=0.132   enclosure: x=0.009 y=0.012
  # m5   size: x=0.100 y=0.108   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.066 0.038 0.066 ;
  LAYER v4   ; RECT -0.029 -0.054 0.029 0.054 ;
  LAYER m5   ; RECT -0.050 -0.054 0.050 0.054 ;
END via4_58Sx108_76V_108H

VIA via4_58Sx108_90V_108H
  # v4   size: x=0.058 y=0.108
  # m4   size: x=0.090 y=0.132   enclosure: x=0.016 y=0.012
  # m5   size: x=0.100 y=0.108   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.066 0.045 0.066 ;
  LAYER v4   ; RECT -0.029 -0.054 0.029 0.054 ;
  LAYER m5   ; RECT -0.050 -0.054 0.050 0.054 ;
END via4_58Sx108_90V_108H

VIA via4_58Sx108_108V_108H
  # v4   size: x=0.058 y=0.108
  # m4   size: x=0.108 y=0.132   enclosure: x=0.025 y=0.012
  # m5   size: x=0.100 y=0.108   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.066 0.054 0.066 ;
  LAYER v4   ; RECT -0.029 -0.054 0.029 0.054 ;
  LAYER m5   ; RECT -0.050 -0.054 0.050 0.054 ;
END via4_58Sx108_108V_108H

VIA via4_58Sx160_76V_160H
  # v4   size: x=0.058 y=0.160
  # m4   size: x=0.076 y=0.184   enclosure: x=0.009 y=0.012
  # m5   size: x=0.100 y=0.160   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.092 0.038 0.092 ;
  LAYER v4   ; RECT -0.029 -0.080 0.029 0.080 ;
  LAYER m5   ; RECT -0.050 -0.080 0.050 0.080 ;
END via4_58Sx160_76V_160H

VIA via4_58Sx160_90V_160H
  # v4   size: x=0.058 y=0.160
  # m4   size: x=0.090 y=0.184   enclosure: x=0.016 y=0.012
  # m5   size: x=0.100 y=0.160   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.092 0.045 0.092 ;
  LAYER v4   ; RECT -0.029 -0.080 0.029 0.080 ;
  LAYER m5   ; RECT -0.050 -0.080 0.050 0.080 ;
END via4_58Sx160_90V_160H

VIA via4_58Sx160_108V_160H
  # v4   size: x=0.058 y=0.160
  # m4   size: x=0.108 y=0.184   enclosure: x=0.025 y=0.012
  # m5   size: x=0.100 y=0.160   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.092 0.054 0.092 ;
  LAYER v4   ; RECT -0.029 -0.080 0.029 0.080 ;
  LAYER m5   ; RECT -0.050 -0.080 0.050 0.080 ;
END via4_58Sx160_108V_160H

VIA via4_58Sx76_76H_76H
  # v4   size: x=0.058 y=0.076
  # m4   size: x=0.082 y=0.076   enclosure: x=0.012 y=0.000
  # m5   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.041 -0.038 0.041 0.038 ;
  LAYER v4   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m5   ; RECT -0.050 -0.038 0.050 0.038 ;
END via4_58Sx76_76H_76H

VIA via4_58Sx76_90H_76H
  # v4   size: x=0.058 y=0.076
  # m4   size: x=0.082 y=0.090   enclosure: x=0.012 y=0.007
  # m5   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.041 -0.045 0.041 0.045 ;
  LAYER v4   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m5   ; RECT -0.050 -0.038 0.050 0.038 ;
END via4_58Sx76_90H_76H

VIA via4_58Sx76_108H_76H
  # v4   size: x=0.058 y=0.076
  # m4   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.016
  # m5   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v4   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m5   ; RECT -0.050 -0.038 0.050 0.038 ;
END via4_58Sx76_108H_76H

VIA via4_58Sx76_76V_76H
  # v4   size: x=0.058 y=0.076
  # m4   size: x=0.076 y=0.100   enclosure: x=0.009 y=0.012
  # m5   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.050 0.038 0.050 ;
  LAYER v4   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m5   ; RECT -0.050 -0.038 0.050 0.038 ;
END via4_58Sx76_76V_76H

VIA via4_58Sx76_90V_76H
  # v4   size: x=0.058 y=0.076
  # m4   size: x=0.090 y=0.100   enclosure: x=0.016 y=0.012
  # m5   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.050 0.045 0.050 ;
  LAYER v4   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m5   ; RECT -0.050 -0.038 0.050 0.038 ;
END via4_58Sx76_90V_76H

VIA via4_58Sx76_108V_76H
  # v4   size: x=0.058 y=0.076
  # m4   size: x=0.108 y=0.100   enclosure: x=0.025 y=0.012
  # m5   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.050 0.054 0.050 ;
  LAYER v4   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m5   ; RECT -0.050 -0.038 0.050 0.038 ;
END via4_58Sx76_108V_76H

VIA via4_58Sx90_76V_90H
  # v4   size: x=0.058 y=0.090
  # m4   size: x=0.076 y=0.114   enclosure: x=0.009 y=0.012
  # m5   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.057 0.038 0.057 ;
  LAYER v4   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m5   ; RECT -0.050 -0.045 0.050 0.045 ;
END via4_58Sx90_76V_90H

VIA via4_58Sx90_90V_90H
  # v4   size: x=0.058 y=0.090
  # m4   size: x=0.090 y=0.114   enclosure: x=0.016 y=0.012
  # m5   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.057 0.045 0.057 ;
  LAYER v4   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m5   ; RECT -0.050 -0.045 0.050 0.045 ;
END via4_58Sx90_90V_90H

VIA via4_58Sx90_108V_90H
  # v4   size: x=0.058 y=0.090
  # m4   size: x=0.108 y=0.114   enclosure: x=0.025 y=0.012
  # m5   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.057 0.054 0.057 ;
  LAYER v4   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m5   ; RECT -0.050 -0.045 0.050 0.045 ;
END via4_58Sx90_108V_90H

VIA via4_58Sx90_108H_90H
  # v4   size: x=0.058 y=0.090
  # m4   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.009
  # m5   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v4   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m5   ; RECT -0.050 -0.045 0.050 0.045 ;
END via4_58Sx90_108H_90H

VIA via4_70x70_56H_90V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.056   enclosure: x=0.012 y=-0.007
  # m5   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.028 0.047 0.028 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.045 -0.056 0.045 0.056 ;
END via4_70x70_56H_90V

VIA via4_70x70_56H_108V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.056   enclosure: x=0.012 y=-0.007
  # m5   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.028 0.047 0.028 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.054 -0.056 0.054 0.056 ;
END via4_70x70_56H_108V

VIA via4_70x70_56H_160V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.056   enclosure: x=0.012 y=-0.007
  # m5   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.028 0.047 0.028 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.080 -0.056 0.080 0.056 ;
END via4_70x70_56H_160V

VIA via4_70x70_76H_90V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m5   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.045 -0.056 0.045 0.056 ;
END via4_70x70_76H_90V

VIA via4_70x70_76H_108V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m5   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.054 -0.056 0.054 0.056 ;
END via4_70x70_76H_108V

VIA via4_70x70_76H_160V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m5   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.080 -0.056 0.080 0.056 ;
END via4_70x70_76H_160V

VIA via4_70x70_90H_90V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m5   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.045 -0.056 0.045 0.056 ;
END via4_70x70_90H_90V

VIA via4_70x70_90H_108V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m5   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.054 -0.056 0.054 0.056 ;
END via4_70x70_90H_108V

VIA via4_70x70_90H_160V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m5   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.080 -0.056 0.080 0.056 ;
END via4_70x70_90H_160V

VIA via4_70x70_108H_90V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m5   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.045 -0.056 0.045 0.056 ;
END via4_70x70_108H_90V

VIA via4_70x70_108H_108V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m5   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.054 -0.056 0.054 0.056 ;
END via4_70x70_108H_108V

VIA via4_70x70_108H_160V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m5   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.080 -0.056 0.080 0.056 ;
END via4_70x70_108H_160V

VIA via4_70x70_108H_200V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m5   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.100 -0.056 0.100 0.056 ;
END via4_70x70_108H_200V

VIA via4_70x70_76V_90V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m5   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.045 -0.056 0.045 0.056 ;
END via4_70x70_76V_90V

VIA via4_70x70_76V_108V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m5   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.054 -0.056 0.054 0.056 ;
END via4_70x70_76V_108V

VIA via4_70x70_76V_160V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m5   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.080 -0.056 0.080 0.056 ;
END via4_70x70_76V_160V

VIA via4_70x70_76V_200V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m5   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.100 -0.056 0.100 0.056 ;
END via4_70x70_76V_200V

VIA via4_70x70_76V_90H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m5   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.045 0.056 0.045 ;
END via4_70x70_76V_90H

VIA via4_70x70_76V_108H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m5   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.054 0.056 0.054 ;
END via4_70x70_76V_108H

VIA via4_70x70_76V_160H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m5   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.080 0.056 0.080 ;
END via4_70x70_76V_160H

VIA via4_70x70_76V_200H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m5   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.100 0.056 0.100 ;
END via4_70x70_76V_200H

VIA via4_70x70_90V_90V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m5   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.045 -0.056 0.045 0.056 ;
END via4_70x70_90V_90V

VIA via4_70x70_90V_108V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m5   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.054 -0.056 0.054 0.056 ;
END via4_70x70_90V_108V

VIA via4_70x70_90V_160V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m5   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.080 -0.056 0.080 0.056 ;
END via4_70x70_90V_160V

VIA via4_70x70_90V_200V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m5   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.100 -0.056 0.100 0.056 ;
END via4_70x70_90V_200V

VIA via4_70x70_90V_90H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m5   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.045 0.056 0.045 ;
END via4_70x70_90V_90H

VIA via4_70x70_90V_108H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m5   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.054 0.056 0.054 ;
END via4_70x70_90V_108H

VIA via4_70x70_90V_160H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m5   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.080 0.056 0.080 ;
END via4_70x70_90V_160H

VIA via4_70x70_90V_200H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m5   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.100 0.056 0.100 ;
END via4_70x70_90V_200H

VIA via4_70x70_108V_90V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m5   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.045 -0.056 0.045 0.056 ;
END via4_70x70_108V_90V

VIA via4_70x70_108V_108V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m5   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.054 -0.056 0.054 0.056 ;
END via4_70x70_108V_108V

VIA via4_70x70_108V_160V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m5   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.080 -0.056 0.080 0.056 ;
END via4_70x70_108V_160V

VIA via4_70x70_108V_200V
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m5   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.100 -0.056 0.100 0.056 ;
END via4_70x70_108V_200V

VIA via4_70x70_108V_90H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m5   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.045 0.056 0.045 ;
END via4_70x70_108V_90H

VIA via4_70x70_108V_108H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m5   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.054 0.056 0.054 ;
END via4_70x70_108V_108H

VIA via4_70x70_108V_160H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m5   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.080 0.056 0.080 ;
END via4_70x70_108V_160H

VIA via4_70x70_108V_200H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m5   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.100 0.056 0.100 ;
END via4_70x70_108V_200H

VIA via4_70x70_90H_90H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m5   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.045 0.056 0.045 ;
END via4_70x70_90H_90H

VIA via4_70x70_90H_108H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m5   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.054 0.056 0.054 ;
END via4_70x70_90H_108H

VIA via4_70x70_90H_160H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m5   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.080 0.056 0.080 ;
END via4_70x70_90H_160H

VIA via4_70x70_90H_200H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m5   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.100 0.056 0.100 ;
END via4_70x70_90H_200H

VIA via4_70x70_108H_90H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m5   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.045 0.056 0.045 ;
END via4_70x70_108H_90H

VIA via4_70x70_108H_108H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m5   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.054 0.056 0.054 ;
END via4_70x70_108H_108H

VIA via4_70x70_108H_160H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m5   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.080 0.056 0.080 ;
END via4_70x70_108H_160H

VIA via4_70x70_108H_200H
  # v4   size: x=0.070 y=0.070
  # m4   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m5   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v4   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m5   ; RECT -0.056 -0.100 0.056 0.100 ;
END via4_70x70_108H_200H

VIA via4_76x58S_76V_76V
  # v4   size: x=0.076 y=0.058
  # m4   size: x=0.076 y=0.082   enclosure: x=0.000 y=0.012
  # m5   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.038 -0.041 0.038 0.041 ;
  LAYER v4   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m5   ; RECT -0.038 -0.050 0.038 0.050 ;
END via4_76x58S_76V_76V

VIA via4_76x58S_90V_76V
  # v4   size: x=0.076 y=0.058
  # m4   size: x=0.090 y=0.082   enclosure: x=0.007 y=0.012
  # m5   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.045 -0.041 0.045 0.041 ;
  LAYER v4   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m5   ; RECT -0.038 -0.050 0.038 0.050 ;
END via4_76x58S_90V_76V

VIA via4_76x58S_108V_76V
  # v4   size: x=0.076 y=0.058
  # m4   size: x=0.108 y=0.082   enclosure: x=0.016 y=0.012
  # m5   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v4   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m5   ; RECT -0.038 -0.050 0.038 0.050 ;
END via4_76x58S_108V_76V

VIA via4_90x58S_108V_90V
  # v4   size: x=0.090 y=0.058
  # m4   size: x=0.108 y=0.082   enclosure: x=0.009 y=0.012
  # m5   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v4   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m5   ; RECT -0.045 -0.050 0.045 0.050 ;
END via4_90x58S_108V_90V

VIA via4_90x90_108H_160V
  # v4   size: x=0.090 y=0.090
  # m4   size: x=0.114 y=0.108   enclosure: x=0.012 y=0.009
  # m5   size: x=0.160 y=0.170   enclosure: x=0.035 y=0.040
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.057 -0.054 0.057 0.054 ;
  LAYER v4   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m5   ; RECT -0.080 -0.085 0.080 0.085 ;
END via4_90x90_108H_160V

VIA via4_90x90_108H_160H
  # v4   size: x=0.090 y=0.090
  # m4   size: x=0.114 y=0.108   enclosure: x=0.012 y=0.009
  # m5   size: x=0.170 y=0.160   enclosure: x=0.040 y=0.035
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.057 -0.054 0.057 0.054 ;
  LAYER v4   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m5   ; RECT -0.085 -0.080 0.085 0.080 ;
END via4_90x90_108H_160H

VIA via4_90x90_108H_200H
  # v4   size: x=0.090 y=0.090
  # m4   size: x=0.114 y=0.108   enclosure: x=0.012 y=0.009
  # m5   size: x=0.170 y=0.200   enclosure: x=0.040 y=0.055
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.057 -0.054 0.057 0.054 ;
  LAYER v4   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m5   ; RECT -0.085 -0.100 0.085 0.100 ;
END via4_90x90_108H_200H

VIA via4_90x90_108V_160V
  # v4   size: x=0.090 y=0.090
  # m4   size: x=0.108 y=0.114   enclosure: x=0.009 y=0.012
  # m5   size: x=0.160 y=0.170   enclosure: x=0.035 y=0.040
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.057 0.054 0.057 ;
  LAYER v4   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m5   ; RECT -0.080 -0.085 0.080 0.085 ;
END via4_90x90_108V_160V

VIA via4_90x90_108V_200V
  # v4   size: x=0.090 y=0.090
  # m4   size: x=0.108 y=0.114   enclosure: x=0.009 y=0.012
  # m5   size: x=0.200 y=0.170   enclosure: x=0.055 y=0.040
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.057 0.054 0.057 ;
  LAYER v4   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m5   ; RECT -0.100 -0.085 0.100 0.085 ;
END via4_90x90_108V_200V

VIA via4_90x90_108V_160H
  # v4   size: x=0.090 y=0.090
  # m4   size: x=0.108 y=0.114   enclosure: x=0.009 y=0.012
  # m5   size: x=0.170 y=0.160   enclosure: x=0.040 y=0.035
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.057 0.054 0.057 ;
  LAYER v4   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m5   ; RECT -0.085 -0.080 0.085 0.080 ;
END via4_90x90_108V_160H

VIA via4_90x90_108V_200H
  # v4   size: x=0.090 y=0.090
  # m4   size: x=0.108 y=0.114   enclosure: x=0.009 y=0.012
  # m5   size: x=0.170 y=0.200   enclosure: x=0.040 y=0.055
  RESISTANCE 1.000 ;
  LAYER m4   ; RECT -0.054 -0.057 0.054 0.057 ;
  LAYER v4   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m5   ; RECT -0.085 -0.100 0.085 0.100 ;
END via4_90x90_108V_200H

VIA via5_108x58S_76H_108V
  # v5   size: x=0.108 y=0.058
  # m5   size: x=0.132 y=0.076   enclosure: x=0.012 y=0.009
  # m6   size: x=0.108 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.066 -0.038 0.066 0.038 ;
  LAYER v5   ; RECT -0.054 -0.029 0.054 0.029 ;
  LAYER m6   ; RECT -0.054 -0.050 0.054 0.050 ;
END via5_108x58S_76H_108V

VIA via5_108x58S_90H_108V
  # v5   size: x=0.108 y=0.058
  # m5   size: x=0.132 y=0.090   enclosure: x=0.012 y=0.016
  # m6   size: x=0.108 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.066 -0.045 0.066 0.045 ;
  LAYER v5   ; RECT -0.054 -0.029 0.054 0.029 ;
  LAYER m6   ; RECT -0.054 -0.050 0.054 0.050 ;
END via5_108x58S_90H_108V

VIA via5_108x58S_108H_108V
  # v5   size: x=0.108 y=0.058
  # m5   size: x=0.132 y=0.108   enclosure: x=0.012 y=0.025
  # m6   size: x=0.108 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.066 -0.054 0.066 0.054 ;
  LAYER v5   ; RECT -0.054 -0.029 0.054 0.029 ;
  LAYER m6   ; RECT -0.054 -0.050 0.054 0.050 ;
END via5_108x58S_108H_108V

VIA via5_108x58S_160H_108V
  # v5   size: x=0.108 y=0.058
  # m5   size: x=0.132 y=0.160   enclosure: x=0.012 y=0.051
  # m6   size: x=0.108 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.066 -0.080 0.066 0.080 ;
  LAYER v5   ; RECT -0.054 -0.029 0.054 0.029 ;
  LAYER m6   ; RECT -0.054 -0.050 0.054 0.050 ;
END via5_108x58S_160H_108V

VIA via5_108x58S_200H_108V
  # v5   size: x=0.108 y=0.058
  # m5   size: x=0.132 y=0.200   enclosure: x=0.012 y=0.071
  # m6   size: x=0.108 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.066 -0.100 0.066 0.100 ;
  LAYER v5   ; RECT -0.054 -0.029 0.054 0.029 ;
  LAYER m6   ; RECT -0.054 -0.050 0.054 0.050 ;
END via5_108x58S_200H_108V

VIA via5_108x58S_160V_108V
  # v5   size: x=0.108 y=0.058
  # m5   size: x=0.160 y=0.082   enclosure: x=0.026 y=0.012
  # m6   size: x=0.108 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.041 0.080 0.041 ;
  LAYER v5   ; RECT -0.054 -0.029 0.054 0.029 ;
  LAYER m6   ; RECT -0.054 -0.050 0.054 0.050 ;
END via5_108x58S_160V_108V

VIA via5_108x58S_200V_108V
  # v5   size: x=0.108 y=0.058
  # m5   size: x=0.200 y=0.082   enclosure: x=0.046 y=0.012
  # m6   size: x=0.108 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.041 0.100 0.041 ;
  LAYER v5   ; RECT -0.054 -0.029 0.054 0.029 ;
  LAYER m6   ; RECT -0.054 -0.050 0.054 0.050 ;
END via5_108x58S_200V_108V

VIA via5_160x58S_76H_160V
  # v5   size: x=0.160 y=0.058
  # m5   size: x=0.184 y=0.076   enclosure: x=0.012 y=0.009
  # m6   size: x=0.160 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.092 -0.038 0.092 0.038 ;
  LAYER v5   ; RECT -0.080 -0.029 0.080 0.029 ;
  LAYER m6   ; RECT -0.080 -0.050 0.080 0.050 ;
END via5_160x58S_76H_160V

VIA via5_160x58S_90H_160V
  # v5   size: x=0.160 y=0.058
  # m5   size: x=0.184 y=0.090   enclosure: x=0.012 y=0.016
  # m6   size: x=0.160 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.092 -0.045 0.092 0.045 ;
  LAYER v5   ; RECT -0.080 -0.029 0.080 0.029 ;
  LAYER m6   ; RECT -0.080 -0.050 0.080 0.050 ;
END via5_160x58S_90H_160V

VIA via5_160x58S_108H_160V
  # v5   size: x=0.160 y=0.058
  # m5   size: x=0.184 y=0.108   enclosure: x=0.012 y=0.025
  # m6   size: x=0.160 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.092 -0.054 0.092 0.054 ;
  LAYER v5   ; RECT -0.080 -0.029 0.080 0.029 ;
  LAYER m6   ; RECT -0.080 -0.050 0.080 0.050 ;
END via5_160x58S_108H_160V

VIA via5_160x58S_160H_160V
  # v5   size: x=0.160 y=0.058
  # m5   size: x=0.184 y=0.160   enclosure: x=0.012 y=0.051
  # m6   size: x=0.160 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.092 -0.080 0.092 0.080 ;
  LAYER v5   ; RECT -0.080 -0.029 0.080 0.029 ;
  LAYER m6   ; RECT -0.080 -0.050 0.080 0.050 ;
END via5_160x58S_160H_160V

VIA via5_160x58S_200H_160V
  # v5   size: x=0.160 y=0.058
  # m5   size: x=0.184 y=0.200   enclosure: x=0.012 y=0.071
  # m6   size: x=0.160 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.092 -0.100 0.092 0.100 ;
  LAYER v5   ; RECT -0.080 -0.029 0.080 0.029 ;
  LAYER m6   ; RECT -0.080 -0.050 0.080 0.050 ;
END via5_160x58S_200H_160V

VIA via5_160x58S_200V_160V
  # v5   size: x=0.160 y=0.058
  # m5   size: x=0.200 y=0.082   enclosure: x=0.020 y=0.012
  # m6   size: x=0.160 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.041 0.100 0.041 ;
  LAYER v5   ; RECT -0.080 -0.029 0.080 0.029 ;
  LAYER m6   ; RECT -0.080 -0.050 0.080 0.050 ;
END via5_160x58S_200V_160V

VIA via5_58Sx108_160H_108H
  # v5   size: x=0.058 y=0.108
  # m5   size: x=0.082 y=0.160   enclosure: x=0.012 y=0.026
  # m6   size: x=0.100 y=0.108   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.080 0.041 0.080 ;
  LAYER v5   ; RECT -0.029 -0.054 0.029 0.054 ;
  LAYER m6   ; RECT -0.050 -0.054 0.050 0.054 ;
END via5_58Sx108_160H_108H

VIA via5_58Sx108_200H_108H
  # v5   size: x=0.058 y=0.108
  # m5   size: x=0.082 y=0.200   enclosure: x=0.012 y=0.046
  # m6   size: x=0.100 y=0.108   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.100 0.041 0.100 ;
  LAYER v5   ; RECT -0.029 -0.054 0.029 0.054 ;
  LAYER m6   ; RECT -0.050 -0.054 0.050 0.054 ;
END via5_58Sx108_200H_108H

VIA via5_58Sx160_200H_160H
  # v5   size: x=0.058 y=0.160
  # m5   size: x=0.082 y=0.200   enclosure: x=0.012 y=0.020
  # m6   size: x=0.100 y=0.160   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.100 0.041 0.100 ;
  LAYER v5   ; RECT -0.029 -0.080 0.029 0.080 ;
  LAYER m6   ; RECT -0.050 -0.080 0.050 0.080 ;
END via5_58Sx160_200H_160H

VIA via5_58Sx44_76H_44H
  # v5   size: x=0.058 y=0.044
  # m5   size: x=0.082 y=0.076   enclosure: x=0.012 y=0.016
  # m6   size: x=0.100 y=0.044   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.038 0.041 0.038 ;
  LAYER v5   ; RECT -0.029 -0.022 0.029 0.022 ;
  LAYER m6   ; RECT -0.050 -0.022 0.050 0.022 ;
END via5_58Sx44_76H_44H

VIA via5_58Sx44_90H_44H
  # v5   size: x=0.058 y=0.044
  # m5   size: x=0.082 y=0.090   enclosure: x=0.012 y=0.023
  # m6   size: x=0.100 y=0.044   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.045 0.041 0.045 ;
  LAYER v5   ; RECT -0.029 -0.022 0.029 0.022 ;
  LAYER m6   ; RECT -0.050 -0.022 0.050 0.022 ;
END via5_58Sx44_90H_44H

VIA via5_58Sx44_108H_44H
  # v5   size: x=0.058 y=0.044
  # m5   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.032
  # m6   size: x=0.100 y=0.044   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v5   ; RECT -0.029 -0.022 0.029 0.022 ;
  LAYER m6   ; RECT -0.050 -0.022 0.050 0.022 ;
END via5_58Sx44_108H_44H

VIA via5_58Sx44_160H_44H
  # v5   size: x=0.058 y=0.044
  # m5   size: x=0.082 y=0.160   enclosure: x=0.012 y=0.058
  # m6   size: x=0.100 y=0.044   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.080 0.041 0.080 ;
  LAYER v5   ; RECT -0.029 -0.022 0.029 0.022 ;
  LAYER m6   ; RECT -0.050 -0.022 0.050 0.022 ;
END via5_58Sx44_160H_44H

VIA via5_58Sx44_200H_44H
  # v5   size: x=0.058 y=0.044
  # m5   size: x=0.082 y=0.200   enclosure: x=0.012 y=0.078
  # m6   size: x=0.100 y=0.044   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.100 0.041 0.100 ;
  LAYER v5   ; RECT -0.029 -0.022 0.029 0.022 ;
  LAYER m6   ; RECT -0.050 -0.022 0.050 0.022 ;
END via5_58Sx44_200H_44H

VIA via5_58Sx56_76H_56H
  # v5   size: x=0.058 y=0.056
  # m5   size: x=0.082 y=0.076   enclosure: x=0.012 y=0.010
  # m6   size: x=0.100 y=0.056   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.038 0.041 0.038 ;
  LAYER v5   ; RECT -0.029 -0.028 0.029 0.028 ;
  LAYER m6   ; RECT -0.050 -0.028 0.050 0.028 ;
END via5_58Sx56_76H_56H

VIA via5_58Sx56_90H_56H
  # v5   size: x=0.058 y=0.056
  # m5   size: x=0.082 y=0.090   enclosure: x=0.012 y=0.017
  # m6   size: x=0.100 y=0.056   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.045 0.041 0.045 ;
  LAYER v5   ; RECT -0.029 -0.028 0.029 0.028 ;
  LAYER m6   ; RECT -0.050 -0.028 0.050 0.028 ;
END via5_58Sx56_90H_56H

VIA via5_58Sx56_108H_56H
  # v5   size: x=0.058 y=0.056
  # m5   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.026
  # m6   size: x=0.100 y=0.056   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v5   ; RECT -0.029 -0.028 0.029 0.028 ;
  LAYER m6   ; RECT -0.050 -0.028 0.050 0.028 ;
END via5_58Sx56_108H_56H

VIA via5_58Sx56_160H_56H
  # v5   size: x=0.058 y=0.056
  # m5   size: x=0.082 y=0.160   enclosure: x=0.012 y=0.052
  # m6   size: x=0.100 y=0.056   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.080 0.041 0.080 ;
  LAYER v5   ; RECT -0.029 -0.028 0.029 0.028 ;
  LAYER m6   ; RECT -0.050 -0.028 0.050 0.028 ;
END via5_58Sx56_160H_56H

VIA via5_58Sx56_200H_56H
  # v5   size: x=0.058 y=0.056
  # m5   size: x=0.082 y=0.200   enclosure: x=0.012 y=0.072
  # m6   size: x=0.100 y=0.056   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.100 0.041 0.100 ;
  LAYER v5   ; RECT -0.029 -0.028 0.029 0.028 ;
  LAYER m6   ; RECT -0.050 -0.028 0.050 0.028 ;
END via5_58Sx56_200H_56H

VIA via5_58Sx76_76H_76H
  # v5   size: x=0.058 y=0.076
  # m5   size: x=0.082 y=0.076   enclosure: x=0.012 y=0.000
  # m6   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.038 0.041 0.038 ;
  LAYER v5   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m6   ; RECT -0.050 -0.038 0.050 0.038 ;
END via5_58Sx76_76H_76H

VIA via5_58Sx76_90H_76H
  # v5   size: x=0.058 y=0.076
  # m5   size: x=0.082 y=0.090   enclosure: x=0.012 y=0.007
  # m6   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.045 0.041 0.045 ;
  LAYER v5   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m6   ; RECT -0.050 -0.038 0.050 0.038 ;
END via5_58Sx76_90H_76H

VIA via5_58Sx76_108H_76H
  # v5   size: x=0.058 y=0.076
  # m5   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.016
  # m6   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v5   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m6   ; RECT -0.050 -0.038 0.050 0.038 ;
END via5_58Sx76_108H_76H

VIA via5_58Sx76_160H_76H
  # v5   size: x=0.058 y=0.076
  # m5   size: x=0.082 y=0.160   enclosure: x=0.012 y=0.042
  # m6   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.080 0.041 0.080 ;
  LAYER v5   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m6   ; RECT -0.050 -0.038 0.050 0.038 ;
END via5_58Sx76_160H_76H

VIA via5_58Sx76_200H_76H
  # v5   size: x=0.058 y=0.076
  # m5   size: x=0.082 y=0.200   enclosure: x=0.012 y=0.062
  # m6   size: x=0.100 y=0.076   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.100 0.041 0.100 ;
  LAYER v5   ; RECT -0.029 -0.038 0.029 0.038 ;
  LAYER m6   ; RECT -0.050 -0.038 0.050 0.038 ;
END via5_58Sx76_200H_76H

VIA via5_58Sx90_108H_90H
  # v5   size: x=0.058 y=0.090
  # m5   size: x=0.082 y=0.108   enclosure: x=0.012 y=0.009
  # m6   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.054 0.041 0.054 ;
  LAYER v5   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m6   ; RECT -0.050 -0.045 0.050 0.045 ;
END via5_58Sx90_108H_90H

VIA via5_58Sx90_160H_90H
  # v5   size: x=0.058 y=0.090
  # m5   size: x=0.082 y=0.160   enclosure: x=0.012 y=0.035
  # m6   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.080 0.041 0.080 ;
  LAYER v5   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m6   ; RECT -0.050 -0.045 0.050 0.045 ;
END via5_58Sx90_160H_90H

VIA via5_58Sx90_200H_90H
  # v5   size: x=0.058 y=0.090
  # m5   size: x=0.082 y=0.200   enclosure: x=0.012 y=0.055
  # m6   size: x=0.100 y=0.090   enclosure: x=0.021 y=0.000
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.041 -0.100 0.041 0.100 ;
  LAYER v5   ; RECT -0.029 -0.045 0.029 0.045 ;
  LAYER m6   ; RECT -0.050 -0.045 0.050 0.045 ;
END via5_58Sx90_200H_90H

VIA via5_70x70_56V_90H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.056 y=0.094   enclosure: x=-0.007 y=0.012
  # m6   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.028 -0.047 0.028 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.045 0.056 0.045 ;
END via5_70x70_56V_90H

VIA via5_70x70_56V_108H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.056 y=0.094   enclosure: x=-0.007 y=0.012
  # m6   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.028 -0.047 0.028 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.054 0.056 0.054 ;
END via5_70x70_56V_108H

VIA via5_70x70_56V_160H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.056 y=0.094   enclosure: x=-0.007 y=0.012
  # m6   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.028 -0.047 0.028 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.080 0.056 0.080 ;
END via5_70x70_56V_160H

VIA via5_70x70_76V_90H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m6   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.045 0.056 0.045 ;
END via5_70x70_76V_90H

VIA via5_70x70_76V_108H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m6   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.054 0.056 0.054 ;
END via5_70x70_76V_108H

VIA via5_70x70_76V_160H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.076 y=0.094   enclosure: x=0.003 y=0.012
  # m6   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.038 -0.047 0.038 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.080 0.056 0.080 ;
END via5_70x70_76V_160H

VIA via5_70x70_90V_90H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m6   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.045 0.056 0.045 ;
END via5_70x70_90V_90H

VIA via5_70x70_90V_108H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m6   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.054 0.056 0.054 ;
END via5_70x70_90V_108H

VIA via5_70x70_90V_160H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m6   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.080 0.056 0.080 ;
END via5_70x70_90V_160H

VIA via5_70x70_108V_90H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m6   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.045 0.056 0.045 ;
END via5_70x70_108V_90H

VIA via5_70x70_108V_108H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m6   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.054 0.056 0.054 ;
END via5_70x70_108V_108H

VIA via5_70x70_108V_160H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m6   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.080 0.056 0.080 ;
END via5_70x70_108V_160H

VIA via5_70x70_108V_200H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m6   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.100 0.056 0.100 ;
END via5_70x70_108V_200H

VIA via5_70x70_108V_400H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m6   size: x=0.112 y=0.400   enclosure: x=0.021 y=0.165
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.200 0.056 0.200 ;
END via5_70x70_108V_400H

VIA via5_70x70_160V_90H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.160 y=0.094   enclosure: x=0.045 y=0.012
  # m6   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.047 0.080 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.045 0.056 0.045 ;
END via5_70x70_160V_90H

VIA via5_70x70_160V_108H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.160 y=0.094   enclosure: x=0.045 y=0.012
  # m6   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.047 0.080 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.054 0.056 0.054 ;
END via5_70x70_160V_108H

VIA via5_70x70_160V_160H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.160 y=0.094   enclosure: x=0.045 y=0.012
  # m6   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.047 0.080 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.080 0.056 0.080 ;
END via5_70x70_160V_160H

VIA via5_70x70_160V_200H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.160 y=0.094   enclosure: x=0.045 y=0.012
  # m6   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.047 0.080 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.100 0.056 0.100 ;
END via5_70x70_160V_200H

VIA via5_70x70_160V_400H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.160 y=0.094   enclosure: x=0.045 y=0.012
  # m6   size: x=0.112 y=0.400   enclosure: x=0.021 y=0.165
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.047 0.080 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.200 0.056 0.200 ;
END via5_70x70_160V_400H

VIA via5_70x70_200V_90H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.200 y=0.094   enclosure: x=0.065 y=0.012
  # m6   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.047 0.100 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.045 0.056 0.045 ;
END via5_70x70_200V_90H

VIA via5_70x70_200V_108H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.200 y=0.094   enclosure: x=0.065 y=0.012
  # m6   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.047 0.100 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.054 0.056 0.054 ;
END via5_70x70_200V_108H

VIA via5_70x70_200V_160H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.200 y=0.094   enclosure: x=0.065 y=0.012
  # m6   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.047 0.100 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.080 0.056 0.080 ;
END via5_70x70_200V_160H

VIA via5_70x70_200V_200H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.200 y=0.094   enclosure: x=0.065 y=0.012
  # m6   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.047 0.100 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.100 0.056 0.100 ;
END via5_70x70_200V_200H

VIA via5_70x70_200V_400H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.200 y=0.094   enclosure: x=0.065 y=0.012
  # m6   size: x=0.112 y=0.400   enclosure: x=0.021 y=0.165
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.047 0.100 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.200 0.056 0.200 ;
END via5_70x70_200V_400H

VIA via5_70x70_76H_90H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m6   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.045 0.056 0.045 ;
END via5_70x70_76H_90H

VIA via5_70x70_76H_108H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m6   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.054 0.056 0.054 ;
END via5_70x70_76H_108H

VIA via5_70x70_76H_160H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m6   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.080 0.056 0.080 ;
END via5_70x70_76H_160H

VIA via5_70x70_76H_200H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m6   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.100 0.056 0.100 ;
END via5_70x70_76H_200H

VIA via5_70x70_76H_400H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m6   size: x=0.112 y=0.400   enclosure: x=0.021 y=0.165
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.200 0.056 0.200 ;
END via5_70x70_76H_400H

VIA via5_70x70_76H_90V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m6   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.045 -0.056 0.045 0.056 ;
END via5_70x70_76H_90V

VIA via5_70x70_76H_108V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m6   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.054 -0.056 0.054 0.056 ;
END via5_70x70_76H_108V

VIA via5_70x70_76H_160V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m6   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.080 -0.056 0.080 0.056 ;
END via5_70x70_76H_160V

VIA via5_70x70_76H_200V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m6   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.100 -0.056 0.100 0.056 ;
END via5_70x70_76H_200V

VIA via5_70x70_76H_400V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.076   enclosure: x=0.012 y=0.003
  # m6   size: x=0.400 y=0.112   enclosure: x=0.165 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.038 0.047 0.038 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.200 -0.056 0.200 0.056 ;
END via5_70x70_76H_400V

VIA via5_70x70_90H_90H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m6   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.045 0.056 0.045 ;
END via5_70x70_90H_90H

VIA via5_70x70_90H_108H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m6   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.054 0.056 0.054 ;
END via5_70x70_90H_108H

VIA via5_70x70_90H_160H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m6   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.080 0.056 0.080 ;
END via5_70x70_90H_160H

VIA via5_70x70_90H_200H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m6   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.100 0.056 0.100 ;
END via5_70x70_90H_200H

VIA via5_70x70_90H_400H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m6   size: x=0.112 y=0.400   enclosure: x=0.021 y=0.165
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.200 0.056 0.200 ;
END via5_70x70_90H_400H

VIA via5_70x70_90H_90V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m6   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.045 -0.056 0.045 0.056 ;
END via5_70x70_90H_90V

VIA via5_70x70_90H_108V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m6   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.054 -0.056 0.054 0.056 ;
END via5_70x70_90H_108V

VIA via5_70x70_90H_160V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m6   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.080 -0.056 0.080 0.056 ;
END via5_70x70_90H_160V

VIA via5_70x70_90H_200V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m6   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.100 -0.056 0.100 0.056 ;
END via5_70x70_90H_200V

VIA via5_70x70_90H_400V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.090   enclosure: x=0.012 y=0.010
  # m6   size: x=0.400 y=0.112   enclosure: x=0.165 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.045 0.047 0.045 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.200 -0.056 0.200 0.056 ;
END via5_70x70_90H_400V

VIA via5_70x70_108H_90H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m6   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.045 0.056 0.045 ;
END via5_70x70_108H_90H

VIA via5_70x70_108H_108H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m6   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.054 0.056 0.054 ;
END via5_70x70_108H_108H

VIA via5_70x70_108H_160H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m6   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.080 0.056 0.080 ;
END via5_70x70_108H_160H

VIA via5_70x70_108H_200H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m6   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.100 0.056 0.100 ;
END via5_70x70_108H_200H

VIA via5_70x70_108H_400H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m6   size: x=0.112 y=0.400   enclosure: x=0.021 y=0.165
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.200 0.056 0.200 ;
END via5_70x70_108H_400H

VIA via5_70x70_108H_90V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m6   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.045 -0.056 0.045 0.056 ;
END via5_70x70_108H_90V

VIA via5_70x70_108H_108V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m6   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.054 -0.056 0.054 0.056 ;
END via5_70x70_108H_108V

VIA via5_70x70_108H_160V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m6   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.080 -0.056 0.080 0.056 ;
END via5_70x70_108H_160V

VIA via5_70x70_108H_200V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m6   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.100 -0.056 0.100 0.056 ;
END via5_70x70_108H_200V

VIA via5_70x70_108H_400V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.108   enclosure: x=0.012 y=0.019
  # m6   size: x=0.400 y=0.112   enclosure: x=0.165 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.054 0.047 0.054 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.200 -0.056 0.200 0.056 ;
END via5_70x70_108H_400V

VIA via5_70x70_160H_90H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.160   enclosure: x=0.012 y=0.045
  # m6   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.080 0.047 0.080 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.045 0.056 0.045 ;
END via5_70x70_160H_90H

VIA via5_70x70_160H_108H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.160   enclosure: x=0.012 y=0.045
  # m6   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.080 0.047 0.080 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.054 0.056 0.054 ;
END via5_70x70_160H_108H

VIA via5_70x70_160H_160H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.160   enclosure: x=0.012 y=0.045
  # m6   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.080 0.047 0.080 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.080 0.056 0.080 ;
END via5_70x70_160H_160H

VIA via5_70x70_160H_200H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.160   enclosure: x=0.012 y=0.045
  # m6   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.080 0.047 0.080 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.100 0.056 0.100 ;
END via5_70x70_160H_200H

VIA via5_70x70_160H_400H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.160   enclosure: x=0.012 y=0.045
  # m6   size: x=0.112 y=0.400   enclosure: x=0.021 y=0.165
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.080 0.047 0.080 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.200 0.056 0.200 ;
END via5_70x70_160H_400H

VIA via5_70x70_160H_90V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.160   enclosure: x=0.012 y=0.045
  # m6   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.080 0.047 0.080 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.045 -0.056 0.045 0.056 ;
END via5_70x70_160H_90V

VIA via5_70x70_160H_108V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.160   enclosure: x=0.012 y=0.045
  # m6   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.080 0.047 0.080 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.054 -0.056 0.054 0.056 ;
END via5_70x70_160H_108V

VIA via5_70x70_160H_160V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.160   enclosure: x=0.012 y=0.045
  # m6   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.080 0.047 0.080 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.080 -0.056 0.080 0.056 ;
END via5_70x70_160H_160V

VIA via5_70x70_160H_200V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.160   enclosure: x=0.012 y=0.045
  # m6   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.080 0.047 0.080 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.100 -0.056 0.100 0.056 ;
END via5_70x70_160H_200V

VIA via5_70x70_160H_400V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.160   enclosure: x=0.012 y=0.045
  # m6   size: x=0.400 y=0.112   enclosure: x=0.165 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.080 0.047 0.080 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.200 -0.056 0.200 0.056 ;
END via5_70x70_160H_400V

VIA via5_70x70_200H_90H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.200   enclosure: x=0.012 y=0.065
  # m6   size: x=0.112 y=0.090   enclosure: x=0.021 y=0.010
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.100 0.047 0.100 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.045 0.056 0.045 ;
END via5_70x70_200H_90H

VIA via5_70x70_200H_108H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.200   enclosure: x=0.012 y=0.065
  # m6   size: x=0.112 y=0.108   enclosure: x=0.021 y=0.019
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.100 0.047 0.100 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.054 0.056 0.054 ;
END via5_70x70_200H_108H

VIA via5_70x70_200H_160H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.200   enclosure: x=0.012 y=0.065
  # m6   size: x=0.112 y=0.160   enclosure: x=0.021 y=0.045
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.100 0.047 0.100 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.080 0.056 0.080 ;
END via5_70x70_200H_160H

VIA via5_70x70_200H_200H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.200   enclosure: x=0.012 y=0.065
  # m6   size: x=0.112 y=0.200   enclosure: x=0.021 y=0.065
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.100 0.047 0.100 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.100 0.056 0.100 ;
END via5_70x70_200H_200H

VIA via5_70x70_200H_400H
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.200   enclosure: x=0.012 y=0.065
  # m6   size: x=0.112 y=0.400   enclosure: x=0.021 y=0.165
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.100 0.047 0.100 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.056 -0.200 0.056 0.200 ;
END via5_70x70_200H_400H

VIA via5_70x70_200H_90V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.200   enclosure: x=0.012 y=0.065
  # m6   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.100 0.047 0.100 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.045 -0.056 0.045 0.056 ;
END via5_70x70_200H_90V

VIA via5_70x70_200H_108V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.200   enclosure: x=0.012 y=0.065
  # m6   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.100 0.047 0.100 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.054 -0.056 0.054 0.056 ;
END via5_70x70_200H_108V

VIA via5_70x70_200H_160V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.200   enclosure: x=0.012 y=0.065
  # m6   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.100 0.047 0.100 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.080 -0.056 0.080 0.056 ;
END via5_70x70_200H_160V

VIA via5_70x70_200H_200V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.200   enclosure: x=0.012 y=0.065
  # m6   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.100 0.047 0.100 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.100 -0.056 0.100 0.056 ;
END via5_70x70_200H_200V

VIA via5_70x70_200H_400V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.094 y=0.200   enclosure: x=0.012 y=0.065
  # m6   size: x=0.400 y=0.112   enclosure: x=0.165 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.047 -0.100 0.047 0.100 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.200 -0.056 0.200 0.056 ;
END via5_70x70_200H_400V

VIA via5_70x70_90V_90V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m6   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.045 -0.056 0.045 0.056 ;
END via5_70x70_90V_90V

VIA via5_70x70_90V_108V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m6   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.054 -0.056 0.054 0.056 ;
END via5_70x70_90V_108V

VIA via5_70x70_90V_160V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m6   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.080 -0.056 0.080 0.056 ;
END via5_70x70_90V_160V

VIA via5_70x70_90V_200V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m6   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.100 -0.056 0.100 0.056 ;
END via5_70x70_90V_200V

VIA via5_70x70_90V_400V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.090 y=0.094   enclosure: x=0.010 y=0.012
  # m6   size: x=0.400 y=0.112   enclosure: x=0.165 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.045 -0.047 0.045 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.200 -0.056 0.200 0.056 ;
END via5_70x70_90V_400V

VIA via5_70x70_108V_90V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m6   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.045 -0.056 0.045 0.056 ;
END via5_70x70_108V_90V

VIA via5_70x70_108V_108V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m6   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.054 -0.056 0.054 0.056 ;
END via5_70x70_108V_108V

VIA via5_70x70_108V_160V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m6   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.080 -0.056 0.080 0.056 ;
END via5_70x70_108V_160V

VIA via5_70x70_108V_200V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m6   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.100 -0.056 0.100 0.056 ;
END via5_70x70_108V_200V

VIA via5_70x70_108V_400V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.108 y=0.094   enclosure: x=0.019 y=0.012
  # m6   size: x=0.400 y=0.112   enclosure: x=0.165 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.047 0.054 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.200 -0.056 0.200 0.056 ;
END via5_70x70_108V_400V

VIA via5_70x70_160V_90V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.160 y=0.094   enclosure: x=0.045 y=0.012
  # m6   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.047 0.080 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.045 -0.056 0.045 0.056 ;
END via5_70x70_160V_90V

VIA via5_70x70_160V_108V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.160 y=0.094   enclosure: x=0.045 y=0.012
  # m6   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.047 0.080 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.054 -0.056 0.054 0.056 ;
END via5_70x70_160V_108V

VIA via5_70x70_160V_160V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.160 y=0.094   enclosure: x=0.045 y=0.012
  # m6   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.047 0.080 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.080 -0.056 0.080 0.056 ;
END via5_70x70_160V_160V

VIA via5_70x70_160V_200V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.160 y=0.094   enclosure: x=0.045 y=0.012
  # m6   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.047 0.080 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.100 -0.056 0.100 0.056 ;
END via5_70x70_160V_200V

VIA via5_70x70_160V_400V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.160 y=0.094   enclosure: x=0.045 y=0.012
  # m6   size: x=0.400 y=0.112   enclosure: x=0.165 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.047 0.080 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.200 -0.056 0.200 0.056 ;
END via5_70x70_160V_400V

VIA via5_70x70_200V_90V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.200 y=0.094   enclosure: x=0.065 y=0.012
  # m6   size: x=0.090 y=0.112   enclosure: x=0.010 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.047 0.100 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.045 -0.056 0.045 0.056 ;
END via5_70x70_200V_90V

VIA via5_70x70_200V_108V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.200 y=0.094   enclosure: x=0.065 y=0.012
  # m6   size: x=0.108 y=0.112   enclosure: x=0.019 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.047 0.100 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.054 -0.056 0.054 0.056 ;
END via5_70x70_200V_108V

VIA via5_70x70_200V_160V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.200 y=0.094   enclosure: x=0.065 y=0.012
  # m6   size: x=0.160 y=0.112   enclosure: x=0.045 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.047 0.100 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.080 -0.056 0.080 0.056 ;
END via5_70x70_200V_160V

VIA via5_70x70_200V_200V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.200 y=0.094   enclosure: x=0.065 y=0.012
  # m6   size: x=0.200 y=0.112   enclosure: x=0.065 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.047 0.100 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.100 -0.056 0.100 0.056 ;
END via5_70x70_200V_200V

VIA via5_70x70_200V_400V
  # v5   size: x=0.070 y=0.070
  # m5   size: x=0.200 y=0.094   enclosure: x=0.065 y=0.012
  # m6   size: x=0.400 y=0.112   enclosure: x=0.165 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.047 0.100 0.047 ;
  LAYER v5   ; RECT -0.035 -0.035 0.035 0.035 ;
  LAYER m6   ; RECT -0.200 -0.056 0.200 0.056 ;
END via5_70x70_200V_400V

VIA via5_76x58S_76V_76V
  # v5   size: x=0.076 y=0.058
  # m5   size: x=0.076 y=0.082   enclosure: x=0.000 y=0.012
  # m6   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.038 -0.041 0.038 0.041 ;
  LAYER v5   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m6   ; RECT -0.038 -0.050 0.038 0.050 ;
END via5_76x58S_76V_76V

VIA via5_76x58S_90V_76V
  # v5   size: x=0.076 y=0.058
  # m5   size: x=0.090 y=0.082   enclosure: x=0.007 y=0.012
  # m6   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.045 -0.041 0.045 0.041 ;
  LAYER v5   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m6   ; RECT -0.038 -0.050 0.038 0.050 ;
END via5_76x58S_90V_76V

VIA via5_76x58S_108V_76V
  # v5   size: x=0.076 y=0.058
  # m5   size: x=0.108 y=0.082   enclosure: x=0.016 y=0.012
  # m6   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v5   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m6   ; RECT -0.038 -0.050 0.038 0.050 ;
END via5_76x58S_108V_76V

VIA via5_76x58S_160V_76V
  # v5   size: x=0.076 y=0.058
  # m5   size: x=0.160 y=0.082   enclosure: x=0.042 y=0.012
  # m6   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.041 0.080 0.041 ;
  LAYER v5   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m6   ; RECT -0.038 -0.050 0.038 0.050 ;
END via5_76x58S_160V_76V

VIA via5_76x58S_200V_76V
  # v5   size: x=0.076 y=0.058
  # m5   size: x=0.200 y=0.082   enclosure: x=0.062 y=0.012
  # m6   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.041 0.100 0.041 ;
  LAYER v5   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m6   ; RECT -0.038 -0.050 0.038 0.050 ;
END via5_76x58S_200V_76V

VIA via5_76x58S_76H_76V
  # v5   size: x=0.076 y=0.058
  # m5   size: x=0.100 y=0.076   enclosure: x=0.012 y=0.009
  # m6   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.050 -0.038 0.050 0.038 ;
  LAYER v5   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m6   ; RECT -0.038 -0.050 0.038 0.050 ;
END via5_76x58S_76H_76V

VIA via5_76x58S_90H_76V
  # v5   size: x=0.076 y=0.058
  # m5   size: x=0.100 y=0.090   enclosure: x=0.012 y=0.016
  # m6   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.050 -0.045 0.050 0.045 ;
  LAYER v5   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m6   ; RECT -0.038 -0.050 0.038 0.050 ;
END via5_76x58S_90H_76V

VIA via5_76x58S_108H_76V
  # v5   size: x=0.076 y=0.058
  # m5   size: x=0.100 y=0.108   enclosure: x=0.012 y=0.025
  # m6   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.050 -0.054 0.050 0.054 ;
  LAYER v5   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m6   ; RECT -0.038 -0.050 0.038 0.050 ;
END via5_76x58S_108H_76V

VIA via5_76x58S_160H_76V
  # v5   size: x=0.076 y=0.058
  # m5   size: x=0.100 y=0.160   enclosure: x=0.012 y=0.051
  # m6   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.050 -0.080 0.050 0.080 ;
  LAYER v5   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m6   ; RECT -0.038 -0.050 0.038 0.050 ;
END via5_76x58S_160H_76V

VIA via5_76x58S_200H_76V
  # v5   size: x=0.076 y=0.058
  # m5   size: x=0.100 y=0.200   enclosure: x=0.012 y=0.071
  # m6   size: x=0.076 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.050 -0.100 0.050 0.100 ;
  LAYER v5   ; RECT -0.038 -0.029 0.038 0.029 ;
  LAYER m6   ; RECT -0.038 -0.050 0.038 0.050 ;
END via5_76x58S_200H_76V

VIA via5_90x58S_76H_90V
  # v5   size: x=0.090 y=0.058
  # m5   size: x=0.114 y=0.076   enclosure: x=0.012 y=0.009
  # m6   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.038 0.057 0.038 ;
  LAYER v5   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m6   ; RECT -0.045 -0.050 0.045 0.050 ;
END via5_90x58S_76H_90V

VIA via5_90x58S_90H_90V
  # v5   size: x=0.090 y=0.058
  # m5   size: x=0.114 y=0.090   enclosure: x=0.012 y=0.016
  # m6   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.045 0.057 0.045 ;
  LAYER v5   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m6   ; RECT -0.045 -0.050 0.045 0.050 ;
END via5_90x58S_90H_90V

VIA via5_90x58S_108H_90V
  # v5   size: x=0.090 y=0.058
  # m5   size: x=0.114 y=0.108   enclosure: x=0.012 y=0.025
  # m6   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.054 0.057 0.054 ;
  LAYER v5   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m6   ; RECT -0.045 -0.050 0.045 0.050 ;
END via5_90x58S_108H_90V

VIA via5_90x58S_160H_90V
  # v5   size: x=0.090 y=0.058
  # m5   size: x=0.114 y=0.160   enclosure: x=0.012 y=0.051
  # m6   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.080 0.057 0.080 ;
  LAYER v5   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m6   ; RECT -0.045 -0.050 0.045 0.050 ;
END via5_90x58S_160H_90V

VIA via5_90x58S_200H_90V
  # v5   size: x=0.090 y=0.058
  # m5   size: x=0.114 y=0.200   enclosure: x=0.012 y=0.071
  # m6   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.100 0.057 0.100 ;
  LAYER v5   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m6   ; RECT -0.045 -0.050 0.045 0.050 ;
END via5_90x58S_200H_90V

VIA via5_90x58S_108V_90V
  # v5   size: x=0.090 y=0.058
  # m5   size: x=0.108 y=0.082   enclosure: x=0.009 y=0.012
  # m6   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.041 0.054 0.041 ;
  LAYER v5   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m6   ; RECT -0.045 -0.050 0.045 0.050 ;
END via5_90x58S_108V_90V

VIA via5_90x58S_160V_90V
  # v5   size: x=0.090 y=0.058
  # m5   size: x=0.160 y=0.082   enclosure: x=0.035 y=0.012
  # m6   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.041 0.080 0.041 ;
  LAYER v5   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m6   ; RECT -0.045 -0.050 0.045 0.050 ;
END via5_90x58S_160V_90V

VIA via5_90x58S_200V_90V
  # v5   size: x=0.090 y=0.058
  # m5   size: x=0.200 y=0.082   enclosure: x=0.055 y=0.012
  # m6   size: x=0.090 y=0.100   enclosure: x=0.000 y=0.021
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.041 0.100 0.041 ;
  LAYER v5   ; RECT -0.045 -0.029 0.045 0.029 ;
  LAYER m6   ; RECT -0.045 -0.050 0.045 0.050 ;
END via5_90x58S_200V_90V

VIA via5_90x90_108V_160H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.108 y=0.114   enclosure: x=0.009 y=0.012
  # m6   size: x=0.170 y=0.160   enclosure: x=0.040 y=0.035
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.057 0.054 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.080 0.085 0.080 ;
END via5_90x90_108V_160H

VIA via5_90x90_108V_160V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.108 y=0.114   enclosure: x=0.009 y=0.012
  # m6   size: x=0.160 y=0.170   enclosure: x=0.035 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.057 0.054 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.080 -0.085 0.080 0.085 ;
END via5_90x90_108V_160V

VIA via5_90x90_108V_200V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.108 y=0.114   enclosure: x=0.009 y=0.012
  # m6   size: x=0.200 y=0.170   enclosure: x=0.055 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.057 0.054 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.100 -0.085 0.100 0.085 ;
END via5_90x90_108V_200V

VIA via5_90x90_108V_400V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.108 y=0.114   enclosure: x=0.009 y=0.012
  # m6   size: x=0.400 y=0.170   enclosure: x=0.155 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.054 -0.057 0.054 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.200 -0.085 0.200 0.085 ;
END via5_90x90_108V_400V

VIA via5_90x90_160V_160H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.160 y=0.114   enclosure: x=0.035 y=0.012
  # m6   size: x=0.170 y=0.160   enclosure: x=0.040 y=0.035
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.057 0.080 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.080 0.085 0.080 ;
END via5_90x90_160V_160H

VIA via5_90x90_160V_160V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.160 y=0.114   enclosure: x=0.035 y=0.012
  # m6   size: x=0.160 y=0.170   enclosure: x=0.035 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.057 0.080 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.080 -0.085 0.080 0.085 ;
END via5_90x90_160V_160V

VIA via5_90x90_160V_200V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.160 y=0.114   enclosure: x=0.035 y=0.012
  # m6   size: x=0.200 y=0.170   enclosure: x=0.055 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.057 0.080 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.100 -0.085 0.100 0.085 ;
END via5_90x90_160V_200V

VIA via5_90x90_160V_400V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.160 y=0.114   enclosure: x=0.035 y=0.012
  # m6   size: x=0.400 y=0.170   enclosure: x=0.155 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.080 -0.057 0.080 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.200 -0.085 0.200 0.085 ;
END via5_90x90_160V_400V

VIA via5_90x90_200V_160H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.200 y=0.114   enclosure: x=0.055 y=0.012
  # m6   size: x=0.170 y=0.160   enclosure: x=0.040 y=0.035
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.057 0.100 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.080 0.085 0.080 ;
END via5_90x90_200V_160H

VIA via5_90x90_200V_160V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.200 y=0.114   enclosure: x=0.055 y=0.012
  # m6   size: x=0.160 y=0.170   enclosure: x=0.035 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.057 0.100 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.080 -0.085 0.080 0.085 ;
END via5_90x90_200V_160V

VIA via5_90x90_200V_200V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.200 y=0.114   enclosure: x=0.055 y=0.012
  # m6   size: x=0.200 y=0.170   enclosure: x=0.055 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.057 0.100 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.100 -0.085 0.100 0.085 ;
END via5_90x90_200V_200V

VIA via5_90x90_200V_400V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.200 y=0.114   enclosure: x=0.055 y=0.012
  # m6   size: x=0.400 y=0.170   enclosure: x=0.155 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.100 -0.057 0.100 0.057 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.200 -0.085 0.200 0.085 ;
END via5_90x90_200V_400V

VIA via5_90x90_108H_160H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.108   enclosure: x=0.012 y=0.009
  # m6   size: x=0.170 y=0.160   enclosure: x=0.040 y=0.035
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.054 0.057 0.054 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.080 0.085 0.080 ;
END via5_90x90_108H_160H

VIA via5_90x90_108H_200H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.108   enclosure: x=0.012 y=0.009
  # m6   size: x=0.170 y=0.200   enclosure: x=0.040 y=0.055
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.054 0.057 0.054 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.100 0.085 0.100 ;
END via5_90x90_108H_200H

VIA via5_90x90_108H_400H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.108   enclosure: x=0.012 y=0.009
  # m6   size: x=0.170 y=0.400   enclosure: x=0.040 y=0.155
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.054 0.057 0.054 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.200 0.085 0.200 ;
END via5_90x90_108H_400H

VIA via5_90x90_108H_160V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.108   enclosure: x=0.012 y=0.009
  # m6   size: x=0.160 y=0.170   enclosure: x=0.035 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.054 0.057 0.054 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.080 -0.085 0.080 0.085 ;
END via5_90x90_108H_160V

VIA via5_90x90_108H_200V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.108   enclosure: x=0.012 y=0.009
  # m6   size: x=0.200 y=0.170   enclosure: x=0.055 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.054 0.057 0.054 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.100 -0.085 0.100 0.085 ;
END via5_90x90_108H_200V

VIA via5_90x90_108H_400V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.108   enclosure: x=0.012 y=0.009
  # m6   size: x=0.400 y=0.170   enclosure: x=0.155 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.054 0.057 0.054 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.200 -0.085 0.200 0.085 ;
END via5_90x90_108H_400V

VIA via5_90x90_160H_160H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.160   enclosure: x=0.012 y=0.035
  # m6   size: x=0.170 y=0.160   enclosure: x=0.040 y=0.035
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.080 0.057 0.080 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.080 0.085 0.080 ;
END via5_90x90_160H_160H

VIA via5_90x90_160H_200H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.160   enclosure: x=0.012 y=0.035
  # m6   size: x=0.170 y=0.200   enclosure: x=0.040 y=0.055
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.080 0.057 0.080 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.100 0.085 0.100 ;
END via5_90x90_160H_200H

VIA via5_90x90_160H_400H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.160   enclosure: x=0.012 y=0.035
  # m6   size: x=0.170 y=0.400   enclosure: x=0.040 y=0.155
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.080 0.057 0.080 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.200 0.085 0.200 ;
END via5_90x90_160H_400H

VIA via5_90x90_160H_160V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.160   enclosure: x=0.012 y=0.035
  # m6   size: x=0.160 y=0.170   enclosure: x=0.035 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.080 0.057 0.080 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.080 -0.085 0.080 0.085 ;
END via5_90x90_160H_160V

VIA via5_90x90_160H_200V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.160   enclosure: x=0.012 y=0.035
  # m6   size: x=0.200 y=0.170   enclosure: x=0.055 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.080 0.057 0.080 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.100 -0.085 0.100 0.085 ;
END via5_90x90_160H_200V

VIA via5_90x90_160H_400V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.160   enclosure: x=0.012 y=0.035
  # m6   size: x=0.400 y=0.170   enclosure: x=0.155 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.080 0.057 0.080 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.200 -0.085 0.200 0.085 ;
END via5_90x90_160H_400V

VIA via5_90x90_200H_160H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.200   enclosure: x=0.012 y=0.055
  # m6   size: x=0.170 y=0.160   enclosure: x=0.040 y=0.035
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.100 0.057 0.100 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.080 0.085 0.080 ;
END via5_90x90_200H_160H

VIA via5_90x90_200H_200H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.200   enclosure: x=0.012 y=0.055
  # m6   size: x=0.170 y=0.200   enclosure: x=0.040 y=0.055
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.100 0.057 0.100 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.100 0.085 0.100 ;
END via5_90x90_200H_200H

VIA via5_90x90_200H_400H
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.200   enclosure: x=0.012 y=0.055
  # m6   size: x=0.170 y=0.400   enclosure: x=0.040 y=0.155
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.100 0.057 0.100 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.085 -0.200 0.085 0.200 ;
END via5_90x90_200H_400H

VIA via5_90x90_200H_160V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.200   enclosure: x=0.012 y=0.055
  # m6   size: x=0.160 y=0.170   enclosure: x=0.035 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.100 0.057 0.100 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.080 -0.085 0.080 0.085 ;
END via5_90x90_200H_160V

VIA via5_90x90_200H_200V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.200   enclosure: x=0.012 y=0.055
  # m6   size: x=0.200 y=0.170   enclosure: x=0.055 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.100 0.057 0.100 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.100 -0.085 0.100 0.085 ;
END via5_90x90_200H_200V

VIA via5_90x90_200H_400V
  # v5   size: x=0.090 y=0.090
  # m5   size: x=0.114 y=0.200   enclosure: x=0.012 y=0.055
  # m6   size: x=0.400 y=0.170   enclosure: x=0.155 y=0.040
  RESISTANCE 1.000 ;
  LAYER m5   ; RECT -0.057 -0.100 0.057 0.100 ;
  LAYER v5   ; RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m6   ; RECT -0.200 -0.085 0.200 0.085 ;
END via5_90x90_200H_400V

VIA via6_120Ux200_160V_180H
  # v6   size: x=0.120 y=0.200
  # m6   size: x=0.160 y=0.320   enclosure: x=0.020 y=0.060
  # m7   size: x=0.240 y=0.180   enclosure: x=0.060 y=-0.010
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.080 -0.160 0.080 0.160 ;
  LAYER v6   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m7   ; RECT -0.120 -0.090 0.120 0.090 ;
END via6_120Ux200_160V_180H

VIA via6_120Ux200_200V_180H
  # v6   size: x=0.120 y=0.200
  # m6   size: x=0.200 y=0.320   enclosure: x=0.040 y=0.060
  # m7   size: x=0.240 y=0.180   enclosure: x=0.060 y=-0.010
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.100 -0.160 0.100 0.160 ;
  LAYER v6   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m7   ; RECT -0.120 -0.090 0.120 0.090 ;
END via6_120Ux200_200V_180H

VIA via6_120Ux200_400V_180H
  # v6   size: x=0.120 y=0.200
  # m6   size: x=0.400 y=0.320   enclosure: x=0.140 y=0.060
  # m7   size: x=0.240 y=0.180   enclosure: x=0.060 y=-0.010
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.200 -0.160 0.200 0.160 ;
  LAYER v6   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m7   ; RECT -0.120 -0.090 0.120 0.090 ;
END via6_120Ux200_400V_180H

VIA via6_120Ux200_400H_180H
  # v6   size: x=0.120 y=0.200
  # m6   size: x=0.240 y=0.400   enclosure: x=0.060 y=0.100
  # m7   size: x=0.240 y=0.180   enclosure: x=0.060 y=-0.010
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.120 -0.200 0.120 0.200 ;
  LAYER v6   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m7   ; RECT -0.120 -0.090 0.120 0.090 ;
END via6_120Ux200_400H_180H

VIA via6_120x200_160V_180V
  # v6   size: x=0.120 y=0.200
  # m6   size: x=0.160 y=0.320   enclosure: x=0.020 y=0.060
  # m7   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.080 -0.160 0.080 0.160 ;
  LAYER v6   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m7   ; RECT -0.090 -0.160 0.090 0.160 ;
END via6_120x200_160V_180V

VIA via6_120x200_200V_180V
  # v6   size: x=0.120 y=0.200
  # m6   size: x=0.200 y=0.320   enclosure: x=0.040 y=0.060
  # m7   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.100 -0.160 0.100 0.160 ;
  LAYER v6   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m7   ; RECT -0.090 -0.160 0.090 0.160 ;
END via6_120x200_200V_180V

VIA via6_120x200_400V_180V
  # v6   size: x=0.120 y=0.200
  # m6   size: x=0.400 y=0.320   enclosure: x=0.140 y=0.060
  # m7   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.200 -0.160 0.200 0.160 ;
  LAYER v6   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m7   ; RECT -0.090 -0.160 0.090 0.160 ;
END via6_120x200_400V_180V

VIA via6_120x200_160V_260H
  # v6   size: x=0.120 y=0.200
  # m6   size: x=0.160 y=0.320   enclosure: x=0.020 y=0.060
  # m7   size: x=0.240 y=0.260   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.080 -0.160 0.080 0.160 ;
  LAYER v6   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m7   ; RECT -0.120 -0.130 0.120 0.130 ;
END via6_120x200_160V_260H

VIA via6_120x200_200V_260H
  # v6   size: x=0.120 y=0.200
  # m6   size: x=0.200 y=0.320   enclosure: x=0.040 y=0.060
  # m7   size: x=0.240 y=0.260   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.100 -0.160 0.100 0.160 ;
  LAYER v6   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m7   ; RECT -0.120 -0.130 0.120 0.130 ;
END via6_120x200_200V_260H

VIA via6_120x200_400V_260H
  # v6   size: x=0.120 y=0.200
  # m6   size: x=0.400 y=0.320   enclosure: x=0.140 y=0.060
  # m7   size: x=0.240 y=0.260   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.200 -0.160 0.200 0.160 ;
  LAYER v6   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m7   ; RECT -0.120 -0.130 0.120 0.130 ;
END via6_120x200_400V_260H

VIA via6_120x200_400H_260H
  # v6   size: x=0.120 y=0.200
  # m6   size: x=0.240 y=0.400   enclosure: x=0.060 y=0.100
  # m7   size: x=0.240 y=0.260   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.120 -0.200 0.120 0.200 ;
  LAYER v6   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m7   ; RECT -0.120 -0.130 0.120 0.130 ;
END via6_120x200_400H_260H

VIA via6_120x400_160V_180V
  # v6   size: x=0.120 y=0.400
  # m6   size: x=0.160 y=0.520   enclosure: x=0.020 y=0.060
  # m7   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.080 -0.260 0.080 0.260 ;
  LAYER v6   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER m7   ; RECT -0.090 -0.260 0.090 0.260 ;
END via6_120x400_160V_180V

VIA via6_120x400_200V_180V
  # v6   size: x=0.120 y=0.400
  # m6   size: x=0.200 y=0.520   enclosure: x=0.040 y=0.060
  # m7   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.100 -0.260 0.100 0.260 ;
  LAYER v6   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER m7   ; RECT -0.090 -0.260 0.090 0.260 ;
END via6_120x400_200V_180V

VIA via6_120x400_400V_180V
  # v6   size: x=0.120 y=0.400
  # m6   size: x=0.400 y=0.520   enclosure: x=0.140 y=0.060
  # m7   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.200 -0.260 0.200 0.260 ;
  LAYER v6   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER m7   ; RECT -0.090 -0.260 0.090 0.260 ;
END via6_120x400_400V_180V

VIA via6_120x400_160V_460H
  # v6   size: x=0.120 y=0.400
  # m6   size: x=0.160 y=0.520   enclosure: x=0.020 y=0.060
  # m7   size: x=0.240 y=0.460   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.080 -0.260 0.080 0.260 ;
  LAYER v6   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER m7   ; RECT -0.120 -0.230 0.120 0.230 ;
END via6_120x400_160V_460H

VIA via6_120x400_200V_460H
  # v6   size: x=0.120 y=0.400
  # m6   size: x=0.200 y=0.520   enclosure: x=0.040 y=0.060
  # m7   size: x=0.240 y=0.460   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.100 -0.260 0.100 0.260 ;
  LAYER v6   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER m7   ; RECT -0.120 -0.230 0.120 0.230 ;
END via6_120x400_200V_460H

VIA via6_120x400_400V_460H
  # v6   size: x=0.120 y=0.400
  # m6   size: x=0.400 y=0.520   enclosure: x=0.140 y=0.060
  # m7   size: x=0.240 y=0.460   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.200 -0.260 0.200 0.260 ;
  LAYER v6   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER m7   ; RECT -0.120 -0.230 0.120 0.230 ;
END via6_120x400_400V_460H

VIA via6_200x120_400H_260V
  # v6   size: x=0.200 y=0.120
  # m6   size: x=0.320 y=0.400   enclosure: x=0.060 y=0.140
  # m7   size: x=0.260 y=0.240   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.160 -0.200 0.160 0.200 ;
  LAYER v6   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m7   ; RECT -0.130 -0.120 0.130 0.120 ;
END via6_200x120_400H_260V

VIA via6_200x120_400V_260V
  # v6   size: x=0.200 y=0.120
  # m6   size: x=0.400 y=0.240   enclosure: x=0.100 y=0.060
  # m7   size: x=0.260 y=0.240   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.200 -0.120 0.200 0.120 ;
  LAYER v6   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m7   ; RECT -0.130 -0.120 0.130 0.120 ;
END via6_200x120_400V_260V

VIA via6_200x120_160H_180H
  # v6   size: x=0.200 y=0.120
  # m6   size: x=0.320 y=0.160   enclosure: x=0.060 y=0.020
  # m7   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.160 -0.080 0.160 0.080 ;
  LAYER v6   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m7   ; RECT -0.160 -0.090 0.160 0.090 ;
END via6_200x120_160H_180H

VIA via6_200x120_200H_180H
  # v6   size: x=0.200 y=0.120
  # m6   size: x=0.320 y=0.200   enclosure: x=0.060 y=0.040
  # m7   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.160 -0.100 0.160 0.100 ;
  LAYER v6   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m7   ; RECT -0.160 -0.090 0.160 0.090 ;
END via6_200x120_200H_180H

VIA via6_200x120_400H_180H
  # v6   size: x=0.200 y=0.120
  # m6   size: x=0.320 y=0.400   enclosure: x=0.060 y=0.140
  # m7   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.160 -0.200 0.160 0.200 ;
  LAYER v6   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m7   ; RECT -0.160 -0.090 0.160 0.090 ;
END via6_200x120_400H_180H

VIA via6_200x120_400V_180H
  # v6   size: x=0.200 y=0.120
  # m6   size: x=0.400 y=0.240   enclosure: x=0.100 y=0.060
  # m7   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.200 -0.120 0.200 0.120 ;
  LAYER v6   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m7   ; RECT -0.160 -0.090 0.160 0.090 ;
END via6_200x120_400V_180H

VIA via6_200x120U_400H_180V
  # v6   size: x=0.200 y=0.120
  # m6   size: x=0.320 y=0.400   enclosure: x=0.060 y=0.140
  # m7   size: x=0.180 y=0.240   enclosure: x=-0.010 y=0.060
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.160 -0.200 0.160 0.200 ;
  LAYER v6   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m7   ; RECT -0.090 -0.120 0.090 0.120 ;
END via6_200x120U_400H_180V

VIA via6_200x120U_400V_180V
  # v6   size: x=0.200 y=0.120
  # m6   size: x=0.400 y=0.240   enclosure: x=0.100 y=0.060
  # m7   size: x=0.180 y=0.240   enclosure: x=-0.010 y=0.060
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.200 -0.120 0.200 0.120 ;
  LAYER v6   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m7   ; RECT -0.090 -0.120 0.090 0.120 ;
END via6_200x120U_400V_180V

VIA via6_400x120_160H_180H
  # v6   size: x=0.400 y=0.120
  # m6   size: x=0.520 y=0.160   enclosure: x=0.060 y=0.020
  # m7   size: x=0.520 y=0.180   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.260 -0.080 0.260 0.080 ;
  LAYER v6   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER m7   ; RECT -0.260 -0.090 0.260 0.090 ;
END via6_400x120_160H_180H

VIA via6_400x120_200H_180H
  # v6   size: x=0.400 y=0.120
  # m6   size: x=0.520 y=0.200   enclosure: x=0.060 y=0.040
  # m7   size: x=0.520 y=0.180   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.260 -0.100 0.260 0.100 ;
  LAYER v6   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER m7   ; RECT -0.260 -0.090 0.260 0.090 ;
END via6_400x120_200H_180H

VIA via6_400x120_400H_180H
  # v6   size: x=0.400 y=0.120
  # m6   size: x=0.520 y=0.400   enclosure: x=0.060 y=0.140
  # m7   size: x=0.520 y=0.180   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m6   ; RECT -0.260 -0.200 0.260 0.200 ;
  LAYER v6   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER m7   ; RECT -0.260 -0.090 0.260 0.090 ;
END via6_400x120_400H_180H

VIA via7_120Ux200_240H_180H
  # v7   size: x=0.120 y=0.200
  # m7   size: x=0.240 y=0.240   enclosure: x=0.060 y=0.020
  # m8   size: x=0.240 y=0.180   enclosure: x=0.060 y=-0.010
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v7   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m8   ; RECT -0.120 -0.090 0.120 0.090 ;
END via7_120Ux200_240H_180H

VIA via7_120x200_180V_180V
  # v7   size: x=0.120 y=0.200
  # m7   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  # m8   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.090 -0.160 0.090 0.160 ;
  LAYER v7   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m8   ; RECT -0.090 -0.160 0.090 0.160 ;
END via7_120x200_180V_180V

VIA via7_120x200_240H_180V
  # v7   size: x=0.120 y=0.200
  # m7   size: x=0.240 y=0.240   enclosure: x=0.060 y=0.020
  # m8   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v7   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m8   ; RECT -0.090 -0.160 0.090 0.160 ;
END via7_120x200_240H_180V

VIA via7_120x200_240H_260H
  # v7   size: x=0.120 y=0.200
  # m7   size: x=0.240 y=0.240   enclosure: x=0.060 y=0.020
  # m8   size: x=0.240 y=0.260   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v7   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER m8   ; RECT -0.120 -0.130 0.120 0.130 ;
END via7_120x200_240H_260H

VIA via7_120x400_180V_180V
  # v7   size: x=0.120 y=0.400
  # m7   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  # m8   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.090 -0.260 0.090 0.260 ;
  LAYER v7   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER m8   ; RECT -0.090 -0.260 0.090 0.260 ;
END via7_120x400_180V_180V

VIA via7_120x400_440H_180V
  # v7   size: x=0.120 y=0.400
  # m7   size: x=0.240 y=0.440   enclosure: x=0.060 y=0.020
  # m8   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.120 -0.220 0.120 0.220 ;
  LAYER v7   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER m8   ; RECT -0.090 -0.260 0.090 0.260 ;
END via7_120x400_440H_180V

VIA via7_120x400_440H_460H
  # v7   size: x=0.120 y=0.400
  # m7   size: x=0.240 y=0.440   enclosure: x=0.060 y=0.020
  # m8   size: x=0.240 y=0.460   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.120 -0.220 0.120 0.220 ;
  LAYER v7   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER m8   ; RECT -0.120 -0.230 0.120 0.230 ;
END via7_120x400_440H_460H

VIA via7_200x120_240V_260V
  # v7   size: x=0.200 y=0.120
  # m7   size: x=0.240 y=0.240   enclosure: x=0.020 y=0.060
  # m8   size: x=0.260 y=0.240   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v7   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m8   ; RECT -0.130 -0.120 0.130 0.120 ;
END via7_200x120_240V_260V

VIA via7_200x120_180H_260V
  # v7   size: x=0.200 y=0.120
  # m7   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  # m8   size: x=0.260 y=0.240   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.160 -0.090 0.160 0.090 ;
  LAYER v7   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m8   ; RECT -0.130 -0.120 0.130 0.120 ;
END via7_200x120_180H_260V

VIA via7_200x120_180H_180H
  # v7   size: x=0.200 y=0.120
  # m7   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  # m8   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.160 -0.090 0.160 0.090 ;
  LAYER v7   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m8   ; RECT -0.160 -0.090 0.160 0.090 ;
END via7_200x120_180H_180H

VIA via7_200x120U_240V_180V
  # v7   size: x=0.200 y=0.120
  # m7   size: x=0.240 y=0.240   enclosure: x=0.020 y=0.060
  # m8   size: x=0.180 y=0.240   enclosure: x=-0.010 y=0.060
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v7   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m8   ; RECT -0.090 -0.120 0.090 0.120 ;
END via7_200x120U_240V_180V

VIA via7_200x120U_180H_180V
  # v7   size: x=0.200 y=0.120
  # m7   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  # m8   size: x=0.180 y=0.240   enclosure: x=-0.010 y=0.060
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.160 -0.090 0.160 0.090 ;
  LAYER v7   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER m8   ; RECT -0.090 -0.120 0.090 0.120 ;
END via7_200x120U_180H_180V

VIA via7_400x120_440V_460V
  # v7   size: x=0.400 y=0.120
  # m7   size: x=0.440 y=0.240   enclosure: x=0.020 y=0.060
  # m8   size: x=0.460 y=0.240   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.220 -0.120 0.220 0.120 ;
  LAYER v7   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER m8   ; RECT -0.230 -0.120 0.230 0.120 ;
END via7_400x120_440V_460V

VIA via7_400x120_180H_460V
  # v7   size: x=0.400 y=0.120
  # m7   size: x=0.520 y=0.180   enclosure: x=0.060 y=0.030
  # m8   size: x=0.460 y=0.240   enclosure: x=0.030 y=0.060
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.260 -0.090 0.260 0.090 ;
  LAYER v7   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER m8   ; RECT -0.230 -0.120 0.230 0.120 ;
END via7_400x120_180H_460V

VIA via7_400x120_180H_180H
  # v7   size: x=0.400 y=0.120
  # m7   size: x=0.520 y=0.180   enclosure: x=0.060 y=0.030
  # m8   size: x=0.520 y=0.180   enclosure: x=0.060 y=0.030
  RESISTANCE 1.000 ;
  LAYER m7   ; RECT -0.260 -0.090 0.260 0.090 ;
  LAYER v7   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER m8   ; RECT -0.260 -0.090 0.260 0.090 ;
END via7_400x120_180H_180H

VIA via8_120x200_180V_1201V
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  # gmz   size: x=1.200 y=0.440   enclosure: x=0.540 y=0.120
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.160 0.090 0.160 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.600 -0.220 0.600 0.220 ;
END via8_120x200_180V_1201V

VIA via8_120x200_180V_1201H
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.360 y=1.200   enclosure: x=0.120 y=0.500
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.160 0.090 0.160 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.180 -0.600 0.180 0.600 ;
END via8_120x200_180V_1201H

VIA via8_120x200_240H_1201V
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.240 y=0.240   enclosure: x=0.060 y=0.020
  # gmz   size: x=1.200 y=0.440   enclosure: x=0.540 y=0.120
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.600 -0.220 0.600 0.220 ;
END via8_120x200_240H_1201V

VIA via8_120x200_240H_1201H
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.240 y=0.240   enclosure: x=0.060 y=0.020
  # gmz   size: x=0.360 y=1.200   enclosure: x=0.120 y=0.500
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.180 -0.600 0.180 0.600 ;
END via8_120x200_240H_1201H

VIA via8_120x200_180V_2401V
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  # gmz   size: x=2.400 y=0.540   enclosure: x=1.140 y=0.170
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.160 0.090 0.160 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -1.200 -0.270 1.200 0.270 ;
END via8_120x200_180V_2401V

VIA via8_120x200_180V_2401H
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.460 y=2.400   enclosure: x=0.170 y=1.100
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.160 0.090 0.160 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.230 -1.200 0.230 1.200 ;
END via8_120x200_180V_2401H

VIA via8_120x200_240H_2401V
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.240 y=0.240   enclosure: x=0.060 y=0.020
  # gmz   size: x=2.400 y=0.540   enclosure: x=1.140 y=0.170
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -1.200 -0.270 1.200 0.270 ;
END via8_120x200_240H_2401V

VIA via8_120x200_240H_2401H
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.240 y=0.240   enclosure: x=0.060 y=0.020
  # gmz   size: x=0.460 y=2.400   enclosure: x=0.170 y=1.100
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.230 -1.200 0.230 1.200 ;
END via8_120x200_240H_2401H

VIA via8_120x200_180V_540V
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.210 y=0.060
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.160 0.090 0.160 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
END via8_120x200_180V_540V

VIA via8_120x200_180V_540H
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.240 y=0.540   enclosure: x=0.060 y=0.170
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.160 0.090 0.160 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.120 -0.270 0.120 0.270 ;
END via8_120x200_180V_540H

VIA via8_120x200_240H_540V
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.240 y=0.240   enclosure: x=0.060 y=0.020
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.210 y=0.060
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
END via8_120x200_240H_540V

VIA via8_120x200_240H_540H
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.240 y=0.240   enclosure: x=0.060 y=0.020
  # gmz   size: x=0.240 y=0.540   enclosure: x=0.060 y=0.170
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.120 -0.270 0.120 0.270 ;
END via8_120x200_240H_540H

VIA via8_120x200_180V_721V
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.720 y=0.370   enclosure: x=0.300 y=0.085
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.160 0.090 0.160 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.360 -0.185 0.360 0.185 ;
END via8_120x200_180V_721V

VIA via8_120x200_180V_721H
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.180 y=0.320   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.290 y=0.720   enclosure: x=0.085 y=0.260
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.160 0.090 0.160 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.145 -0.360 0.145 0.360 ;
END via8_120x200_180V_721H

VIA via8_120x200_240H_721V
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.240 y=0.240   enclosure: x=0.060 y=0.020
  # gmz   size: x=0.720 y=0.370   enclosure: x=0.300 y=0.085
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.360 -0.185 0.360 0.185 ;
END via8_120x200_240H_721V

VIA via8_120x200_240H_721H
  # v8   size: x=0.120 y=0.200
  # m8   size: x=0.240 y=0.240   enclosure: x=0.060 y=0.020
  # gmz   size: x=0.290 y=0.720   enclosure: x=0.085 y=0.260
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gmz  ; RECT -0.145 -0.360 0.145 0.360 ;
END via8_120x200_240H_721H

VIA via8_120x400_180V_1201V
  # v8   size: x=0.120 y=0.400
  # m8   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  # gmz   size: x=1.200 y=0.640   enclosure: x=0.540 y=0.120
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.260 0.090 0.260 ;
  LAYER v8   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gmz  ; RECT -0.600 -0.320 0.600 0.320 ;
END via8_120x400_180V_1201V

VIA via8_120x400_180V_1201H
  # v8   size: x=0.120 y=0.400
  # m8   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.360 y=1.200   enclosure: x=0.120 y=0.400
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.260 0.090 0.260 ;
  LAYER v8   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gmz  ; RECT -0.180 -0.600 0.180 0.600 ;
END via8_120x400_180V_1201H

VIA via8_120x400_440H_1201H
  # v8   size: x=0.120 y=0.400
  # m8   size: x=0.240 y=0.440   enclosure: x=0.060 y=0.020
  # gmz   size: x=0.360 y=1.200   enclosure: x=0.120 y=0.400
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.220 0.120 0.220 ;
  LAYER v8   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gmz  ; RECT -0.180 -0.600 0.180 0.600 ;
END via8_120x400_440H_1201H

VIA via8_120x400_180V_2401V
  # v8   size: x=0.120 y=0.400
  # m8   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  # gmz   size: x=2.400 y=0.740   enclosure: x=1.140 y=0.170
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.260 0.090 0.260 ;
  LAYER v8   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gmz  ; RECT -1.200 -0.370 1.200 0.370 ;
END via8_120x400_180V_2401V

VIA via8_120x400_180V_2401H
  # v8   size: x=0.120 y=0.400
  # m8   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.460 y=2.400   enclosure: x=0.170 y=1.000
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.260 0.090 0.260 ;
  LAYER v8   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gmz  ; RECT -0.230 -1.200 0.230 1.200 ;
END via8_120x400_180V_2401H

VIA via8_120x400_440H_2401H
  # v8   size: x=0.120 y=0.400
  # m8   size: x=0.240 y=0.440   enclosure: x=0.060 y=0.020
  # gmz   size: x=0.460 y=2.400   enclosure: x=0.170 y=1.000
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.220 0.120 0.220 ;
  LAYER v8   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gmz  ; RECT -0.230 -1.200 0.230 1.200 ;
END via8_120x400_440H_2401H

VIA via8_120x400_180V_540V
  # v8   size: x=0.120 y=0.400
  # m8   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.540 y=0.520   enclosure: x=0.210 y=0.060
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.260 0.090 0.260 ;
  LAYER v8   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gmz  ; RECT -0.270 -0.260 0.270 0.260 ;
END via8_120x400_180V_540V

VIA via8_120x400_180V_540H
  # v8   size: x=0.120 y=0.400
  # m8   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.240 y=0.540   enclosure: x=0.060 y=0.070
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.260 0.090 0.260 ;
  LAYER v8   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gmz  ; RECT -0.120 -0.270 0.120 0.270 ;
END via8_120x400_180V_540H

VIA via8_120x400_180V_721V
  # v8   size: x=0.120 y=0.400
  # m8   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.720 y=0.570   enclosure: x=0.300 y=0.085
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.260 0.090 0.260 ;
  LAYER v8   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gmz  ; RECT -0.360 -0.285 0.360 0.285 ;
END via8_120x400_180V_721V

VIA via8_120x400_180V_721H
  # v8   size: x=0.120 y=0.400
  # m8   size: x=0.180 y=0.520   enclosure: x=0.030 y=0.060
  # gmz   size: x=0.290 y=0.720   enclosure: x=0.085 y=0.160
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.090 -0.260 0.090 0.260 ;
  LAYER v8   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gmz  ; RECT -0.145 -0.360 0.145 0.360 ;
END via8_120x400_180V_721H

VIA via8_120x400_440H_721H
  # v8   size: x=0.120 y=0.400
  # m8   size: x=0.240 y=0.440   enclosure: x=0.060 y=0.020
  # gmz   size: x=0.290 y=0.720   enclosure: x=0.085 y=0.160
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.220 0.120 0.220 ;
  LAYER v8   ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gmz  ; RECT -0.145 -0.360 0.145 0.360 ;
END via8_120x400_440H_721H

VIA via8_200x120_240V_1201V
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.240 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=1.200 y=0.360   enclosure: x=0.500 y=0.120
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.600 -0.180 0.600 0.180 ;
END via8_200x120_240V_1201V

VIA via8_200x120_240V_1201H
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.240 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.440 y=1.200   enclosure: x=0.120 y=0.540
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.220 -0.600 0.220 0.600 ;
END via8_200x120_240V_1201H

VIA via8_200x120_180H_1201V
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  # gmz   size: x=1.200 y=0.360   enclosure: x=0.500 y=0.120
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.160 -0.090 0.160 0.090 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.600 -0.180 0.600 0.180 ;
END via8_200x120_180H_1201V

VIA via8_200x120_180H_1201H
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  # gmz   size: x=0.440 y=1.200   enclosure: x=0.120 y=0.540
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.160 -0.090 0.160 0.090 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.220 -0.600 0.220 0.600 ;
END via8_200x120_180H_1201H

VIA via8_200x120_240V_2401V
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.240 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=2.400 y=0.460   enclosure: x=1.100 y=0.170
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -1.200 -0.230 1.200 0.230 ;
END via8_200x120_240V_2401V

VIA via8_200x120_240V_2401H
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.240 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.540 y=2.400   enclosure: x=0.170 y=1.140
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.270 -1.200 0.270 1.200 ;
END via8_200x120_240V_2401H

VIA via8_200x120_180H_2401V
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  # gmz   size: x=2.400 y=0.460   enclosure: x=1.100 y=0.170
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.160 -0.090 0.160 0.090 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -1.200 -0.230 1.200 0.230 ;
END via8_200x120_180H_2401V

VIA via8_200x120_180H_2401H
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  # gmz   size: x=0.540 y=2.400   enclosure: x=0.170 y=1.140
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.160 -0.090 0.160 0.090 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.270 -1.200 0.270 1.200 ;
END via8_200x120_180H_2401H

VIA via8_200x120_240V_540V
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.240 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.540 y=0.240   enclosure: x=0.170 y=0.060
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.270 -0.120 0.270 0.120 ;
END via8_200x120_240V_540V

VIA via8_200x120_240V_540H
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.240 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.060 y=0.210
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
END via8_200x120_240V_540H

VIA via8_200x120_180H_540V
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  # gmz   size: x=0.540 y=0.240   enclosure: x=0.170 y=0.060
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.160 -0.090 0.160 0.090 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.270 -0.120 0.270 0.120 ;
END via8_200x120_180H_540V

VIA via8_200x120_180H_540H
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.060 y=0.210
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.160 -0.090 0.160 0.090 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
END via8_200x120_180H_540H

VIA via8_200x120_240V_721V
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.240 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.720 y=0.290   enclosure: x=0.260 y=0.085
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.360 -0.145 0.360 0.145 ;
END via8_200x120_240V_721V

VIA via8_200x120_240V_721H
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.240 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.370 y=0.720   enclosure: x=0.085 y=0.300
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.120 -0.120 0.120 0.120 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.185 -0.360 0.185 0.360 ;
END via8_200x120_240V_721H

VIA via8_200x120_180H_721V
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  # gmz   size: x=0.720 y=0.290   enclosure: x=0.260 y=0.085
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.160 -0.090 0.160 0.090 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.360 -0.145 0.360 0.145 ;
END via8_200x120_180H_721V

VIA via8_200x120_180H_721H
  # v8   size: x=0.200 y=0.120
  # m8   size: x=0.320 y=0.180   enclosure: x=0.060 y=0.030
  # gmz   size: x=0.370 y=0.720   enclosure: x=0.085 y=0.300
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.160 -0.090 0.160 0.090 ;
  LAYER v8   ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gmz  ; RECT -0.185 -0.360 0.185 0.360 ;
END via8_200x120_180H_721H

VIA via8_400x120_440V_1201V
  # v8   size: x=0.400 y=0.120
  # m8   size: x=0.440 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=1.200 y=0.360   enclosure: x=0.400 y=0.120
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.220 -0.120 0.220 0.120 ;
  LAYER v8   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gmz  ; RECT -0.600 -0.180 0.600 0.180 ;
END via8_400x120_440V_1201V

VIA via8_400x120_440V_1201H
  # v8   size: x=0.400 y=0.120
  # m8   size: x=0.440 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.640 y=1.200   enclosure: x=0.120 y=0.540
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.220 -0.120 0.220 0.120 ;
  LAYER v8   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gmz  ; RECT -0.320 -0.600 0.320 0.600 ;
END via8_400x120_440V_1201H

VIA via8_400x120_440V_2401V
  # v8   size: x=0.400 y=0.120
  # m8   size: x=0.440 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=2.400 y=0.460   enclosure: x=1.000 y=0.170
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.220 -0.120 0.220 0.120 ;
  LAYER v8   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gmz  ; RECT -1.200 -0.230 1.200 0.230 ;
END via8_400x120_440V_2401V

VIA via8_400x120_440V_2401H
  # v8   size: x=0.400 y=0.120
  # m8   size: x=0.440 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.740 y=2.400   enclosure: x=0.170 y=1.140
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.220 -0.120 0.220 0.120 ;
  LAYER v8   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gmz  ; RECT -0.370 -1.200 0.370 1.200 ;
END via8_400x120_440V_2401H

VIA via8_400x120_180H_2401H
  # v8   size: x=0.400 y=0.120
  # m8   size: x=0.520 y=0.180   enclosure: x=0.060 y=0.030
  # gmz   size: x=0.740 y=2.400   enclosure: x=0.170 y=1.140
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.260 -0.090 0.260 0.090 ;
  LAYER v8   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gmz  ; RECT -0.370 -1.200 0.370 1.200 ;
END via8_400x120_180H_2401H

VIA via8_400x120_440V_540V
  # v8   size: x=0.400 y=0.120
  # m8   size: x=0.440 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.540 y=0.240   enclosure: x=0.070 y=0.060
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.220 -0.120 0.220 0.120 ;
  LAYER v8   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gmz  ; RECT -0.270 -0.120 0.270 0.120 ;
END via8_400x120_440V_540V

VIA via8_400x120_440V_540H
  # v8   size: x=0.400 y=0.120
  # m8   size: x=0.440 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.520 y=0.540   enclosure: x=0.060 y=0.210
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.220 -0.120 0.220 0.120 ;
  LAYER v8   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gmz  ; RECT -0.260 -0.270 0.260 0.270 ;
END via8_400x120_440V_540H

VIA via8_400x120_440V_721V
  # v8   size: x=0.400 y=0.120
  # m8   size: x=0.440 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.720 y=0.290   enclosure: x=0.160 y=0.085
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.220 -0.120 0.220 0.120 ;
  LAYER v8   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gmz  ; RECT -0.360 -0.145 0.360 0.145 ;
END via8_400x120_440V_721V

VIA via8_400x120_440V_721H
  # v8   size: x=0.400 y=0.120
  # m8   size: x=0.440 y=0.240   enclosure: x=0.020 y=0.060
  # gmz   size: x=0.570 y=0.720   enclosure: x=0.085 y=0.300
  RESISTANCE 1.000 ;
  LAYER m8   ; RECT -0.220 -0.120 0.220 0.120 ;
  LAYER v8   ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gmz  ; RECT -0.285 -0.360 0.285 0.360 ;
END via8_400x120_440V_721H

VIA GV0_1850x800_2130V_3050V
  # gv0   size: x=1.850 y=0.800
  # gm0   size: x=2.130 y=1.080   enclosure: x=0.140 y=0.140
  # gmb   size: x=3.050 y=2.000   enclosure: x=0.600 y=0.600
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.065 -0.540 1.065 0.540 ;
  LAYER gv0  ; RECT -0.925 -0.400 0.925 0.400 ;
  LAYER gmb  ; RECT -1.525 -1.000 1.525 1.000 ;
END GV0_1850x800_2130V_3050V

VIA GV0_1850x800_1080H_2000H
  # gv0   size: x=1.850 y=0.800
  # gm0   size: x=2.130 y=1.080   enclosure: x=0.140 y=0.140
  # gmb   size: x=3.050 y=2.000   enclosure: x=0.600 y=0.600
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.065 -0.540 1.065 0.540 ;
  LAYER gv0  ; RECT -0.925 -0.400 0.925 0.400 ;
  LAYER gmb  ; RECT -1.525 -1.000 1.525 1.000 ;
END GV0_1850x800_1080H_2000H

VIA GV0_3700x800_3980V_4900V
  # gv0   size: x=3.700 y=0.800
  # gm0   size: x=3.980 y=1.080   enclosure: x=0.140 y=0.140
  # gmb   size: x=4.900 y=2.000   enclosure: x=0.600 y=0.600
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.990 -0.540 1.990 0.540 ;
  LAYER gv0  ; RECT -1.850 -0.400 1.850 0.400 ;
  LAYER gmb  ; RECT -2.450 -1.000 2.450 1.000 ;
END GV0_3700x800_3980V_4900V

VIA GV0_3700x800_1080H_2000H
  # gv0   size: x=3.700 y=0.800
  # gm0   size: x=3.980 y=1.080   enclosure: x=0.140 y=0.140
  # gmb   size: x=4.900 y=2.000   enclosure: x=0.600 y=0.600
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -1.990 -0.540 1.990 0.540 ;
  LAYER gv0  ; RECT -1.850 -0.400 1.850 0.400 ;
  LAYER gmb  ; RECT -2.450 -1.000 2.450 1.000 ;
END GV0_3700x800_1080H_2000H

VIA GV0_800x1850_1080V_2000V
  # gv0   size: x=0.800 y=1.850
  # gm0   size: x=1.080 y=2.130   enclosure: x=0.140 y=0.140
  # gmb   size: x=2.000 y=3.050   enclosure: x=0.600 y=0.600
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.540 -1.065 0.540 1.065 ;
  LAYER gv0  ; RECT -0.400 -0.925 0.400 0.925 ;
  LAYER gmb  ; RECT -1.000 -1.525 1.000 1.525 ;
END GV0_800x1850_1080V_2000V

VIA GV0_800x1850_2130H_3050H
  # gv0   size: x=0.800 y=1.850
  # gm0   size: x=1.080 y=2.130   enclosure: x=0.140 y=0.140
  # gmb   size: x=2.000 y=3.050   enclosure: x=0.600 y=0.600
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.540 -1.065 0.540 1.065 ;
  LAYER gv0  ; RECT -0.400 -0.925 0.400 0.925 ;
  LAYER gmb  ; RECT -1.000 -1.525 1.000 1.525 ;
END GV0_800x1850_2130H_3050H

VIA GV0_800x3700_1080V_2000V
  # gv0   size: x=0.800 y=3.700
  # gm0   size: x=1.080 y=3.980   enclosure: x=0.140 y=0.140
  # gmb   size: x=2.000 y=4.900   enclosure: x=0.600 y=0.600
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.540 -1.990 0.540 1.990 ;
  LAYER gv0  ; RECT -0.400 -1.850 0.400 1.850 ;
  LAYER gmb  ; RECT -1.000 -2.450 1.000 2.450 ;
END GV0_800x3700_1080V_2000V

VIA GV0_800x3700_3980H_4900H
  # gv0   size: x=0.800 y=3.700
  # gm0   size: x=1.080 y=3.980   enclosure: x=0.140 y=0.140
  # gmb   size: x=2.000 y=4.900   enclosure: x=0.600 y=0.600
  RESISTANCE 1.000 ;
  LAYER gm0  ; RECT -0.540 -1.990 0.540 1.990 ;
  LAYER gv0  ; RECT -0.400 -1.850 0.400 1.850 ;
  LAYER gmb  ; RECT -1.000 -2.450 1.000 2.450 ;
END GV0_800x3700_3980H_4900H

VIA VMZ_120x200_540V_1201H
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.540 y=0.340   enclosure: x=0.210 y=0.070
  # gm0   size: x=0.360 y=1.200   enclosure: x=0.120 y=0.500
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.170 0.270 0.170 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.180 -0.600 0.180 0.600 ;
END VMZ_120x200_540V_1201H

VIA VMZ_120x200_540V_1201V
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.540 y=0.340   enclosure: x=0.210 y=0.070
  # gm0   size: x=1.200 y=0.440   enclosure: x=0.540 y=0.120
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.170 0.270 0.170 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.600 -0.220 0.600 0.220 ;
END VMZ_120x200_540V_1201V

VIA VMZ_120x200_540V_2401H
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.540 y=0.340   enclosure: x=0.210 y=0.070
  # gm0   size: x=0.460 y=2.400   enclosure: x=0.170 y=1.100
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.170 0.270 0.170 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.230 -1.200 0.230 1.200 ;
END VMZ_120x200_540V_2401H

VIA VMZ_120x200_540V_2401V
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.540 y=0.340   enclosure: x=0.210 y=0.070
  # gm0   size: x=2.400 y=0.540   enclosure: x=1.140 y=0.170
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.170 0.270 0.170 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -1.200 -0.270 1.200 0.270 ;
END VMZ_120x200_540V_2401V

VIA VMZ_120x200_540V_540H
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.540 y=0.340   enclosure: x=0.210 y=0.070
  # gm0   size: x=0.240 y=0.540   enclosure: x=0.060 y=0.170
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.170 0.270 0.170 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.120 -0.270 0.120 0.270 ;
END VMZ_120x200_540V_540H

VIA VMZ_120x200_540V_540V
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.540 y=0.340   enclosure: x=0.210 y=0.070
  # gm0   size: x=0.540 y=0.320   enclosure: x=0.210 y=0.060
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.170 0.270 0.170 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.270 -0.160 0.270 0.160 ;
END VMZ_120x200_540V_540V

VIA VMZ_120x200_540V_721H
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.540 y=0.340   enclosure: x=0.210 y=0.070
  # gm0   size: x=0.290 y=0.720   enclosure: x=0.085 y=0.260
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.170 0.270 0.170 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.145 -0.360 0.145 0.360 ;
END VMZ_120x200_540V_721H

VIA VMZ_120x200_540V_721V
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.540 y=0.340   enclosure: x=0.210 y=0.070
  # gm0   size: x=0.720 y=0.370   enclosure: x=0.300 y=0.085
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.170 0.270 0.170 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.360 -0.185 0.360 0.185 ;
END VMZ_120x200_540V_721V

VIA VMZ_120x200_540H_1201H
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.100 y=0.170
  # gm0   size: x=0.360 y=1.200   enclosure: x=0.120 y=0.500
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.180 -0.600 0.180 0.600 ;
END VMZ_120x200_540H_1201H

VIA VMZ_120x200_540H_1201V
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.100 y=0.170
  # gm0   size: x=1.200 y=0.440   enclosure: x=0.540 y=0.120
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.600 -0.220 0.600 0.220 ;
END VMZ_120x200_540H_1201V

VIA VMZ_120x200_540H_2401H
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.100 y=0.170
  # gm0   size: x=0.460 y=2.400   enclosure: x=0.170 y=1.100
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.230 -1.200 0.230 1.200 ;
END VMZ_120x200_540H_2401H

VIA VMZ_120x200_540H_2401V
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.100 y=0.170
  # gm0   size: x=2.400 y=0.540   enclosure: x=1.140 y=0.170
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -1.200 -0.270 1.200 0.270 ;
END VMZ_120x200_540H_2401V

VIA VMZ_120x200_540H_540H
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.100 y=0.170
  # gm0   size: x=0.240 y=0.540   enclosure: x=0.060 y=0.170
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.120 -0.270 0.120 0.270 ;
END VMZ_120x200_540H_540H

VIA VMZ_120x200_540H_540V
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.100 y=0.170
  # gm0   size: x=0.540 y=0.320   enclosure: x=0.210 y=0.060
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.270 -0.160 0.270 0.160 ;
END VMZ_120x200_540H_540V

VIA VMZ_120x200_540H_721H
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.100 y=0.170
  # gm0   size: x=0.290 y=0.720   enclosure: x=0.085 y=0.260
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.145 -0.360 0.145 0.360 ;
END VMZ_120x200_540H_721H

VIA VMZ_120x200_540H_721V
  # vmz   size: x=0.120 y=0.200
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.100 y=0.170
  # gm0   size: x=0.720 y=0.370   enclosure: x=0.300 y=0.085
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.100 0.060 0.100 ;
  LAYER gm0  ; RECT -0.360 -0.185 0.360 0.185 ;
END VMZ_120x200_540H_721V

VIA VMZ_120x400_540V_2401V
  # vmz   size: x=0.120 y=0.400
  # gmz   size: x=0.540 y=0.540   enclosure: x=0.210 y=0.070
  # gm0   size: x=2.400 y=0.740   enclosure: x=1.140 y=0.170
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.270 0.270 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gm0  ; RECT -1.200 -0.370 1.200 0.370 ;
END VMZ_120x400_540V_2401V

VIA VMZ_120x400_540H_1201H
  # vmz   size: x=0.120 y=0.400
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.100 y=0.070
  # gm0   size: x=0.360 y=1.200   enclosure: x=0.120 y=0.400
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gm0  ; RECT -0.180 -0.600 0.180 0.600 ;
END VMZ_120x400_540H_1201H

VIA VMZ_120x400_540H_2401H
  # vmz   size: x=0.120 y=0.400
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.100 y=0.070
  # gm0   size: x=0.460 y=2.400   enclosure: x=0.170 y=1.000
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gm0  ; RECT -0.230 -1.200 0.230 1.200 ;
END VMZ_120x400_540H_2401H

VIA VMZ_120x400_540H_721H
  # vmz   size: x=0.120 y=0.400
  # gmz   size: x=0.320 y=0.540   enclosure: x=0.100 y=0.070
  # gm0   size: x=0.290 y=0.720   enclosure: x=0.085 y=0.160
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.160 -0.270 0.160 0.270 ;
  LAYER vmz  ; RECT -0.060 -0.200 0.060 0.200 ;
  LAYER gm0  ; RECT -0.145 -0.360 0.145 0.360 ;
END VMZ_120x400_540H_721H

VIA VMZ_200x120_540H_1201H
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.340 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.440 y=1.200   enclosure: x=0.120 y=0.540
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.170 -0.270 0.170 0.270 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.220 -0.600 0.220 0.600 ;
END VMZ_200x120_540H_1201H

VIA VMZ_200x120_540H_1201V
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.340 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=1.200 y=0.360   enclosure: x=0.500 y=0.120
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.170 -0.270 0.170 0.270 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.600 -0.180 0.600 0.180 ;
END VMZ_200x120_540H_1201V

VIA VMZ_200x120_540H_2401H
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.340 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.540 y=2.400   enclosure: x=0.170 y=1.140
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.170 -0.270 0.170 0.270 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.270 -1.200 0.270 1.200 ;
END VMZ_200x120_540H_2401H

VIA VMZ_200x120_540H_2401V
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.340 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=2.400 y=0.460   enclosure: x=1.100 y=0.170
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.170 -0.270 0.170 0.270 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -1.200 -0.230 1.200 0.230 ;
END VMZ_200x120_540H_2401V

VIA VMZ_200x120_540H_540H
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.340 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.320 y=0.540   enclosure: x=0.060 y=0.210
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.170 -0.270 0.170 0.270 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.160 -0.270 0.160 0.270 ;
END VMZ_200x120_540H_540H

VIA VMZ_200x120_540H_540V
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.340 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.540 y=0.240   enclosure: x=0.170 y=0.060
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.170 -0.270 0.170 0.270 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.270 -0.120 0.270 0.120 ;
END VMZ_200x120_540H_540V

VIA VMZ_200x120_540H_721H
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.340 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.370 y=0.720   enclosure: x=0.085 y=0.300
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.170 -0.270 0.170 0.270 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.185 -0.360 0.185 0.360 ;
END VMZ_200x120_540H_721H

VIA VMZ_200x120_540H_721V
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.340 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.720 y=0.290   enclosure: x=0.260 y=0.085
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.170 -0.270 0.170 0.270 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.360 -0.145 0.360 0.145 ;
END VMZ_200x120_540H_721V

VIA VMZ_200x120_540V_1201H
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.170 y=0.100
  # gm0   size: x=0.440 y=1.200   enclosure: x=0.120 y=0.540
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.220 -0.600 0.220 0.600 ;
END VMZ_200x120_540V_1201H

VIA VMZ_200x120_540V_1201V
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.170 y=0.100
  # gm0   size: x=1.200 y=0.360   enclosure: x=0.500 y=0.120
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.600 -0.180 0.600 0.180 ;
END VMZ_200x120_540V_1201V

VIA VMZ_200x120_540V_2401H
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.170 y=0.100
  # gm0   size: x=0.540 y=2.400   enclosure: x=0.170 y=1.140
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.270 -1.200 0.270 1.200 ;
END VMZ_200x120_540V_2401H

VIA VMZ_200x120_540V_2401V
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.170 y=0.100
  # gm0   size: x=2.400 y=0.460   enclosure: x=1.100 y=0.170
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -1.200 -0.230 1.200 0.230 ;
END VMZ_200x120_540V_2401V

VIA VMZ_200x120_540V_540H
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.170 y=0.100
  # gm0   size: x=0.320 y=0.540   enclosure: x=0.060 y=0.210
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.160 -0.270 0.160 0.270 ;
END VMZ_200x120_540V_540H

VIA VMZ_200x120_540V_540V
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.170 y=0.100
  # gm0   size: x=0.540 y=0.240   enclosure: x=0.170 y=0.060
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.270 -0.120 0.270 0.120 ;
END VMZ_200x120_540V_540V

VIA VMZ_200x120_540V_721H
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.170 y=0.100
  # gm0   size: x=0.370 y=0.720   enclosure: x=0.085 y=0.300
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.185 -0.360 0.185 0.360 ;
END VMZ_200x120_540V_721H

VIA VMZ_200x120_540V_721V
  # vmz   size: x=0.200 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.170 y=0.100
  # gm0   size: x=0.720 y=0.290   enclosure: x=0.260 y=0.085
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.100 -0.060 0.100 0.060 ;
  LAYER gm0  ; RECT -0.360 -0.145 0.360 0.145 ;
END VMZ_200x120_540V_721V

VIA VMZ_400x120_540H_1201H
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.640 y=1.200   enclosure: x=0.120 y=0.540
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.270 0.270 0.270 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.320 -0.600 0.320 0.600 ;
END VMZ_400x120_540H_1201H

VIA VMZ_400x120_540H_1201V
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=1.200 y=0.360   enclosure: x=0.400 y=0.120
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.270 0.270 0.270 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.600 -0.180 0.600 0.180 ;
END VMZ_400x120_540H_1201V

VIA VMZ_400x120_540H_2401H
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.740 y=2.400   enclosure: x=0.170 y=1.140
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.270 0.270 0.270 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.370 -1.200 0.370 1.200 ;
END VMZ_400x120_540H_2401H

VIA VMZ_400x120_540H_2401V
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=2.400 y=0.460   enclosure: x=1.000 y=0.170
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.270 0.270 0.270 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -1.200 -0.230 1.200 0.230 ;
END VMZ_400x120_540H_2401V

VIA VMZ_400x120_540H_540H
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.520 y=0.540   enclosure: x=0.060 y=0.210
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.270 0.270 0.270 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.260 -0.270 0.260 0.270 ;
END VMZ_400x120_540H_540H

VIA VMZ_400x120_540H_540V
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.540 y=0.240   enclosure: x=0.070 y=0.060
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.270 0.270 0.270 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.270 -0.120 0.270 0.120 ;
END VMZ_400x120_540H_540V

VIA VMZ_400x120_540H_721H
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.570 y=0.720   enclosure: x=0.085 y=0.300
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.270 0.270 0.270 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.285 -0.360 0.285 0.360 ;
END VMZ_400x120_540H_721H

VIA VMZ_400x120_540H_721V
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.540   enclosure: x=0.070 y=0.210
  # gm0   size: x=0.720 y=0.290   enclosure: x=0.160 y=0.085
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.270 0.270 0.270 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.360 -0.145 0.360 0.145 ;
END VMZ_400x120_540H_721V

VIA VMZ_400x120_540V_1201H
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.070 y=0.100
  # gm0   size: x=0.640 y=1.200   enclosure: x=0.120 y=0.540
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.320 -0.600 0.320 0.600 ;
END VMZ_400x120_540V_1201H

VIA VMZ_400x120_540V_1201V
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.070 y=0.100
  # gm0   size: x=1.200 y=0.360   enclosure: x=0.400 y=0.120
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.600 -0.180 0.600 0.180 ;
END VMZ_400x120_540V_1201V

VIA VMZ_400x120_540V_2401H
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.070 y=0.100
  # gm0   size: x=0.740 y=2.400   enclosure: x=0.170 y=1.140
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.370 -1.200 0.370 1.200 ;
END VMZ_400x120_540V_2401H

VIA VMZ_400x120_540V_2401V
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.070 y=0.100
  # gm0   size: x=2.400 y=0.460   enclosure: x=1.000 y=0.170
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -1.200 -0.230 1.200 0.230 ;
END VMZ_400x120_540V_2401V

VIA VMZ_400x120_540V_540H
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.070 y=0.100
  # gm0   size: x=0.520 y=0.540   enclosure: x=0.060 y=0.210
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.260 -0.270 0.260 0.270 ;
END VMZ_400x120_540V_540H

VIA VMZ_400x120_540V_540V
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.070 y=0.100
  # gm0   size: x=0.540 y=0.240   enclosure: x=0.070 y=0.060
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.270 -0.120 0.270 0.120 ;
END VMZ_400x120_540V_540V

VIA VMZ_400x120_540V_721H
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.070 y=0.100
  # gm0   size: x=0.570 y=0.720   enclosure: x=0.085 y=0.300
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.285 -0.360 0.285 0.360 ;
END VMZ_400x120_540V_721H

VIA VMZ_400x120_540V_721V
  # vmz   size: x=0.400 y=0.120
  # gmz   size: x=0.540 y=0.320   enclosure: x=0.070 y=0.100
  # gm0   size: x=0.720 y=0.290   enclosure: x=0.160 y=0.085
  RESISTANCE 1.000 ;
  LAYER gmz  ; RECT -0.270 -0.160 0.270 0.160 ;
  LAYER vmz  ; RECT -0.200 -0.060 0.200 0.060 ;
  LAYER gm0  ; RECT -0.360 -0.145 0.360 0.145 ;
END VMZ_400x120_540V_721V

##################################################
# Via Map Table 
##################################################
# |-------------------------------------------------------------------------------------------|
# | Via Map Table                                                                             |
# |-------------------------------------------------------------------------------------------|
# | This table specifies which specific via to use given a metal width below and above.       |
# | If a via is specified in this table, it should also include the "DEFAULT" keyword in      |
# | the previous Via Definitions section.                                                     |
# |-------------------------------------------------------------------------------------------|
# | The format of the via map table is:                                                       |
# |                                                                                           |
# | VIA  Cut_layer  Lower_metal_width  Upper_metal_width  Via_name                            |
# | ---  ---------  -----------------  -----------------  -------------------------           |
# | VIA     v1         0.020             0.068            via1_20Sx68_20V_68H                 |
# | VIA     v5         0.064             0.108            via5_52Sx108_64V_108H               |
# |-------------------------------------------------------------------------------------------|
# | NOTE                                                                                      |
# |-------------------------------------------------------------------------------------------|
# | Dummy vias are created to include all metal width transitions in the via map table. Dummy |
# | vias are not drc clean and not intended to be used, but exist to prevent routing errors   |
# | occurring for an incomplete via map table.                                                |
# |-------------------------------------------------------------------------------------------|

PROPERTYDEFINITIONS
 LIBRARY LEF58_METALWIDTHVIAMAP STRING "
  METALWIDTHVIAMAP
   VIA   v1    0.068              0.044               VIA1_60SX44_68V_44H
   VIA   v1    0.068              0.056               VIA1_60SX56_68V_56H
   VIA   v1    0.068              0.076               VIA1_60SX76_68V_76H
   VIA   v1    0.068              0.09                VIA1_60SX90_68V_90H
   VIA   v1    0.068              0.108               VIA1_60SX108_68V_108H
   VIA   v1    0.1                0.044               VIA1_60SX44_100V_44H
   VIA   v1    0.1                0.056               VIA1_60SX56_100V_56H
   VIA   v1    0.1                0.076               VIA1_60SX76_100V_76H
   VIA   v1    0.1                0.09                VIA1_60SX90_100V_90H
   VIA   v1    0.1                0.108               VIA1_60SX108_100V_108H
   VIA   v2    0.044              0.044               VIA2_44X58S_44H_44V
   VIA   v2    0.044              0.056               VIA2_56X58S_44H_56V
   VIA   v2    0.044              0.076               VIA2_76X58S_44H_76V
   VIA   v2    0.044              0.09                VIA2_90X58S_44H_90V
   VIA   v2    0.044              0.108               VIA2_108X58S_44H_108V
   VIA   v2    0.056              0.044               VIA2_44X58S_56H_44V
   VIA   v2    0.056              0.056               VIA2_56X58S_56H_56V
   VIA   v2    0.056              0.076               VIA2_76X58S_56H_76V
   VIA   v2    0.056              0.09                VIA2_90X58S_56H_90V
   VIA   v2    0.056              0.108               VIA2_108X58S_56H_108V
   VIA   v2    0.076              0.044               VIA2_44X58S_76H_44V
   VIA   v2    0.076              0.056               VIA2_56X58S_76H_56V
   VIA   v2    0.076              0.076               VIA2_76X58S_76H_76V
   VIA   v2    0.076              0.09                VIA2_90X58S_76H_90V
   VIA   v2    0.076              0.108               VIA2_108X58S_76H_108V
   VIA   v2    0.09               0.044               VIA2_44X58S_90H_44V
   VIA   v2    0.09               0.056               VIA2_56X58S_90H_56V
   VIA   v2    0.09               0.076               VIA2_76X58S_90H_76V
   VIA   v2    0.09               0.09                VIA2_90X58S_90H_90V
   VIA   v2    0.09               0.108               VIA2_108X58S_90H_108V
   VIA   v2    0.108              0.044               VIA2_44X58S_108H_44V
   VIA   v2    0.108              0.056               VIA2_56X58S_108H_56V
   VIA   v2    0.108              0.076               VIA2_76X58S_108H_76V
   VIA   v2    0.108              0.09                VIA2_90X58S_108H_90V
   VIA   v2    0.108              0.108               VIA2_108X58S_108H_108V
   VIA   v3    0.044              0.044               VIA3_58SX44_44V_44H
   VIA   v3    0.044              0.056               VIA3_58SX56_44V_56H
   VIA   v3    0.044              0.076               VIA3_58SX76_44V_76H
   VIA   v3    0.044              0.09                VIA3_58SX90_44V_90H
   VIA   v3    0.044              0.108               VIA3_58SX108_44V_108H
   VIA   v3    0.056              0.044               VIA3_58SX44_56V_44H
   VIA   v3    0.056              0.056               VIA3_58SX56_56V_56H
   VIA   v3    0.056              0.076               VIA3_58SX76_56V_76H
   VIA   v3    0.056              0.09                VIA3_58SX90_56V_90H
   VIA   v3    0.056              0.108               VIA3_58SX108_56V_108H
   VIA   v3    0.076              0.044               VIA3_58SX44_76V_44H
   VIA   v3    0.076              0.056               VIA3_58SX56_76V_56H
   VIA   v3    0.076              0.076               VIA3_58SX76_76V_76H
   VIA   v3    0.076              0.09                VIA3_58SX90_76V_90H
   VIA   v3    0.076              0.108               VIA3_58SX108_76V_108H
   VIA   v3    0.09               0.044               VIA3_58SX44_90V_44H
   VIA   v3    0.09               0.056               VIA3_58SX56_90V_56H
   VIA   v3    0.09               0.076               VIA3_58SX76_90V_76H
   VIA   v3    0.09               0.09                VIA3_58SX90_90V_90H
   VIA   v3    0.09               0.108               VIA3_58SX108_90V_108H
   VIA   v3    0.108              0.044               VIA3_58SX44_108V_44H
   VIA   v3    0.108              0.056               VIA3_58SX56_108V_56H
   VIA   v3    0.108              0.076               VIA3_58SX76_108V_76H
   VIA   v3    0.108              0.09                VIA3_58SX90_108V_90H
   VIA   v3    0.108              0.108               VIA3_58SX108_108V_108H
   VIA   v4    0.044              0.044               VIA4_44X58S_44H_44V
   VIA   v4    0.044              0.056               VIA4_56X58S_44H_56V
   VIA   v4    0.044              0.076               VIA4_76X58S_44H_76V
   VIA   v4    0.044              0.09                VIA4_90X58S_44H_90V
   VIA   v4    0.044              0.108               VIA4_108X58S_44H_108V
   VIA   v4    0.044              0.16                VIA4_160X58S_44H_160V
   VIA   v4    0.044              0.2                 VIA4_70X70_56H_200V
   VIA   v4    0.056              0.044               VIA4_44X58S_56H_44V
   VIA   v4    0.056              0.056               VIA4_56X58S_56H_56V
   VIA   v4    0.056              0.076               VIA4_76X58S_56H_76V
   VIA   v4    0.056              0.09                VIA4_90X58S_56H_90V
   VIA   v4    0.056              0.108               VIA4_108X58S_56H_108V
   VIA   v4    0.056              0.16                VIA4_160X58S_56H_160V
   VIA   v4    0.056              0.2                 VIA4_70X70_56H_200V
   VIA   v4    0.076              0.044               VIA4_44X58S_76H_44V
   VIA   v4    0.076              0.056               VIA4_56X58S_76H_56V
   VIA   v4    0.076              0.076               VIA4_76X58S_76H_76V
   VIA   v4    0.076              0.09                VIA4_90X58S_76H_90V
   VIA   v4    0.076              0.108               VIA4_108X58S_76H_108V
   VIA   v4    0.076              0.16                VIA4_160X58S_76H_160V
   VIA   v4    0.076              0.2                 VIA4_70X70_76H_200V
   VIA   v4    0.09               0.044               VIA4_44X58S_90H_44V
   VIA   v4    0.09               0.056               VIA4_56X58S_90H_56V
   VIA   v4    0.09               0.076               VIA4_76X58S_90H_76V
   VIA   v4    0.09               0.09                VIA4_90X58S_90H_90V
   VIA   v4    0.09               0.108               VIA4_108X58S_90H_108V
   VIA   v4    0.09               0.16                VIA4_160X58S_90H_160V
   VIA   v4    0.09               0.2                 VIA4_70X70_90H_200V
   VIA   v4    0.108              0.044               VIA4_44X58S_108H_44V
   VIA   v4    0.108              0.056               VIA4_56X58S_108H_56V
   VIA   v4    0.108              0.076               VIA4_76X58S_108H_76V
   VIA   v4    0.108              0.09                VIA4_90X58S_108H_90V
   VIA   v4    0.108              0.108               VIA4_108X58S_108H_108V
   VIA   v4    0.108              0.16                VIA4_160X58S_108H_160V
   VIA   v4    0.108              0.2                 VIA4_90X90_108H_200V
   VIA   v5    0.044              0.044               VIA5_58SX44_44V_44H
   VIA   v5    0.044              0.056               VIA5_58SX56_44V_56H
   VIA   v5    0.044              0.076               VIA5_58SX76_44V_76H
   VIA   v5    0.044              0.09                VIA5_58SX90_44V_90H
   VIA   v5    0.044              0.108               VIA5_58SX108_44V_108H
   VIA   v5    0.044              0.16                VIA5_58SX160_44V_160H
   VIA   v5    0.044              0.2                 VIA5_70X70_56V_200H
   VIA   v5    0.044              0.4                 VIA5_70X70_56V_400H
   VIA   v5    0.056              0.044               VIA5_58SX44_56V_44H
   VIA   v5    0.056              0.056               VIA5_58SX56_56V_56H
   VIA   v5    0.056              0.076               VIA5_58SX76_56V_76H
   VIA   v5    0.056              0.09                VIA5_58SX90_56V_90H
   VIA   v5    0.056              0.108               VIA5_58SX108_56V_108H
   VIA   v5    0.056              0.16                VIA5_58SX160_56V_160H
   VIA   v5    0.056              0.2                 VIA5_70X70_56V_200H
   VIA   v5    0.056              0.4                 VIA5_70X70_56V_400H
   VIA   v5    0.076              0.044               VIA5_58SX44_76V_44H
   VIA   v5    0.076              0.056               VIA5_58SX56_76V_56H
   VIA   v5    0.076              0.076               VIA5_58SX76_76V_76H
   VIA   v5    0.076              0.09                VIA5_58SX90_76V_90H
   VIA   v5    0.076              0.108               VIA5_58SX108_76V_108H
   VIA   v5    0.076              0.16                VIA5_58SX160_76V_160H
   VIA   v5    0.076              0.2                 VIA5_70X70_76V_200H
   VIA   v5    0.076              0.4                 VIA5_70X70_76V_400H
   VIA   v5    0.09               0.044               VIA5_58SX44_90V_44H
   VIA   v5    0.09               0.056               VIA5_58SX56_90V_56H
   VIA   v5    0.09               0.076               VIA5_58SX76_90V_76H
   VIA   v5    0.09               0.09                VIA5_58SX90_90V_90H
   VIA   v5    0.09               0.108               VIA5_58SX108_90V_108H
   VIA   v5    0.09               0.16                VIA5_58SX160_90V_160H
   VIA   v5    0.09               0.2                 VIA5_70X70_90V_200H
   VIA   v5    0.09               0.4                 VIA5_70X70_90V_400H
   VIA   v5    0.108              0.044               VIA5_58SX44_108V_44H
   VIA   v5    0.108              0.056               VIA5_58SX56_108V_56H
   VIA   v5    0.108              0.076               VIA5_58SX76_108V_76H
   VIA   v5    0.108              0.09                VIA5_58SX90_108V_90H
   VIA   v5    0.108              0.108               VIA5_58SX108_108V_108H
   VIA   v5    0.108              0.16                VIA5_58SX160_108V_160H
   VIA   v5    0.108              0.2                 VIA5_90X90_108V_200H
   VIA   v5    0.108              0.4                 VIA5_90X90_108V_400H
   VIA   v5    0.16               0.044               VIA5_58SX44_160V_44H
   VIA   v5    0.16               0.056               VIA5_58SX56_160V_56H
   VIA   v5    0.16               0.076               VIA5_58SX76_160V_76H
   VIA   v5    0.16               0.09                VIA5_58SX90_160V_90H
   VIA   v5    0.16               0.108               VIA5_58SX108_160V_108H
   VIA   v5    0.16               0.16                VIA5_58SX160_160V_160H
   VIA   v5    0.16               0.2                 VIA5_90X90_160V_200H
   VIA   v5    0.16               0.4                 VIA5_90X90_160V_400H
   VIA   v5    0.2                0.044               VIA5_58SX44_200V_44H
   VIA   v5    0.2                0.056               VIA5_58SX56_200V_56H
   VIA   v5    0.2                0.076               VIA5_58SX76_200V_76H
   VIA   v5    0.2                0.09                VIA5_58SX90_200V_90H
   VIA   v5    0.2                0.108               VIA5_58SX108_200V_108H
   VIA   v5    0.2                0.16                VIA5_58SX160_200V_160H
   VIA   v5    0.2                0.2                 VIA5_90X90_200V_200H
   VIA   v5    0.2                0.4                 VIA5_90X90_200V_400H
   VIA   v6    0.044 0.16         0.18 0.18           VIA6_200X120U_160H_180V
   VIA   v6    0.044 0.16         0.26 0.4            VIA6_200X120_160H_260V
   VIA   v6    0.044 0.16         0.46 0.9            VIA6_400X120_160H_460V
   VIA   v6    0.2 0.2            0.18 0.18           VIA6_200X120U_200H_180V
   VIA   v6    0.2 0.2            0.26 0.4            VIA6_200X120_200H_260V
   VIA   v6    0.2 0.2            0.46 0.9            VIA6_400X120_200H_460V
   VIA   v6    0.4 0.4            0.18 0.4            VIA6_120X200_400H_180V
   VIA   v6    0.4 0.4            0.46 0.9            VIA6_400X120_400H_460V
   VIA   v7    0.18 0.4           0.18 0.18           VIA7_120UX200_180V_180H
   VIA   v7    0.18 0.4           0.181 0.19          VIA7_200X120_240V_180H
   VIA   v7    0.18 0.4           0.26 0.4            VIA7_120X200_180V_260H
   VIA   v7    0.18 0.5           0.46 0.9            VIA7_120X400_180V_460H
   VIA   v7    0.46 0.9           0.18 0.4            VIA7_400X120_440V_180H
   VIA   v7    0.6 0.6            0.46 0.46           via7_120x400_600V_460H_ARRAY_2x1
   VIA   v7    0.6 0.6            0.5 0.5             via7_120x400_600V_500H_ARRAY_2x1
   VIA   v7    0.6 0.6            0.6 0.6             via7_120x400_600V_600H_ARRAY_2x1
   VIA   v7    0.6 0.6            0.7 0.7             via7_120x400_600V_700H_ARRAY_2x1
   VIA   v7    0.6 0.6            0.8 0.8             via7_120x400_600V_800H_ARRAY_2x1
   VIA   v7    0.6 0.6            0.9 0.9             via7_120x400_600V_900H_ARRAY_2x1
   VIA   v7    0.7 0.7            0.46 0.46           via7_120x400_700V_460H_ARRAY_2x1
   VIA   v7    0.7 0.7            0.5 0.5             via7_120x400_700V_500H_ARRAY_2x1
   VIA   v7    0.7 0.7            0.6 0.6             via7_120x400_700V_600H_ARRAY_2x1
   VIA   v7    0.7 0.7            0.7 0.7             via7_120x400_700V_700H_ARRAY_2x1
   VIA   v7    0.7 0.7            0.8 0.8             via7_120x400_700V_800H_ARRAY_2x1
   VIA   v7    0.7 0.7            0.9 0.9             via7_120x400_700V_900H_ARRAY_2x1
   VIA   v7    0.8 0.8            0.46 0.46           via7_120x400_800V_460H_ARRAY_2x1
   VIA   v7    0.8 0.8            0.5 0.5             via7_120x400_800V_500H_ARRAY_2x1
   VIA   v7    0.8 0.8            0.6 0.6             via7_120x400_800V_600H_ARRAY_2x1
   VIA   v7    0.8 0.8            0.7 0.7             via7_120x400_800V_700H_ARRAY_2x1
   VIA   v7    0.8 0.8            0.8 0.8             via7_120x400_800V_800H_ARRAY_2x1
   VIA   v7    0.8 0.8            0.9 0.9             via7_120x400_800V_900H_ARRAY_2x1
   VIA   v7    0.9 0.9            0.46 0.46           via7_120x400_900V_460H_ARRAY_2x1
   VIA   v7    0.9 0.9            0.5 0.5             via7_120x400_900V_500H_ARRAY_2x1
   VIA   v7    0.9 0.9            0.6 0.6             via7_120x400_900V_600H_ARRAY_2x1
   VIA   v7    0.9 0.9            0.7 0.7             via7_120x400_900V_700H_ARRAY_2x1
   VIA   v7    0.9 0.9            0.8 0.8             via7_120x400_900V_800H_ARRAY_2x1
   VIA   v7    0.9 0.9            0.9 0.9             via7_120x400_900V_900H_ARRAY_2x1
   VIA   v8    0.18 0.4           0.54 0.54           VIA8_400X120_180H_540V
   VIA   v8    0.18 0.4           0.721 0.721         VIA8_400X120_180H_721V
   VIA   v8    0.18 0.4           1.201 1.201         VIA8_400X120_180H_1201V
   VIA   v8    0.18 0.4           2.401 2.401         VIA8_400X120_180H_2401V
   VIA   v8    0.46 0.9           0.54 0.54           VIA8_120X400_440H_540V
   VIA   v8    0.46 0.9           0.721 0.721         VIA8_120X400_440H_721V
   VIA   v8    0.46 0.9           1.201 1.201         VIA8_120X400_440H_1201V
   VIA   v8    0.46 0.9           2.401 2.401         VIA8_120X400_440H_2401V
   VIA   v8    0.18 0.4           0.54 0.54           VIA8_400X120_180H_540H PGVIA
   VIA   v8    0.18 0.4           0.721 0.721         VIA8_400X120_180H_721H PGVIA
   VIA   v8    0.18 0.4           1.201 1.201         VIA8_400X120_180H_1201H PGVIA
   VIA   v8    0.18 0.18          2.401 2.401         via8_400x120_180H_2401V_ARRAY_3x1 PGVIA
   VIA   v8    0.181 0.181        2.401 2.401         via8_400x120_181H_2401V_ARRAY_3x1 PGVIA
   VIA   v8    0.19 0.19          2.401 2.401         via8_400x120_190H_2401V_ARRAY_3x1 PGVIA
   VIA   v8    0.26 0.26          2.401 2.401         via8_400x120_260H_2401V_ARRAY_3x1 PGVIA
   VIA   v8    0.3 0.3            2.401 2.401         via8_400x120_300H_2401V_ARRAY_3x1 PGVIA
   VIA   v8    0.4 0.4            2.401 2.401         via8_400x120_400H_2401V_ARRAY_3x1 PGVIA
   VIA   v8    0.46 0.9           0.54 0.54           VIA8_120X400_440H_540H PGVIA
   VIA   v8    0.46 0.46          0.721 0.721         via8_120x400_460H_721V_ARRAY_2x1 PGVIA
   VIA   v8    0.46 0.46          1.201 1.201         via8_120x400_460H_1201V_ARRAY_3x1 PGVIA
   VIA   v8    0.46 0.46          2.401 2.401         via8_120x400_460H_2401V_ARRAY_6x1 PGVIA
   VIA   v8    0.5 0.5            0.721 0.721         via8_120x400_500H_721V_ARRAY_2x1 PGVIA
   VIA   v8    0.5 0.5            1.201 1.201         via8_120x400_500H_1201V_ARRAY_3x1 PGVIA
   VIA   v8    0.5 0.5            2.401 2.401         via8_120x400_500H_2401V_ARRAY_6x1 PGVIA
   VIA   v8    0.6 0.6            0.721 0.721         via8_120x400_600H_721V_ARRAY_2x1 PGVIA
   VIA   v8    0.6 0.6            1.201 1.201         via8_120x400_600H_1201V_ARRAY_3x1 PGVIA
   VIA   v8    0.6 0.6            2.401 2.401         via8_120x400_600H_2401V_ARRAY_6x1 PGVIA
   VIA   v8    0.7 0.7            0.721 0.721         via8_120x400_700H_721V_ARRAY_2x1 PGVIA
   VIA   v8    0.7 0.7            1.201 1.201         via8_120x400_700H_1201V_ARRAY_3x1 PGVIA
   VIA   v8    0.7 0.7            2.401 2.401         via8_120x400_700H_2401V_ARRAY_6x1 PGVIA
   VIA   v8    0.8 0.8            0.721 0.721         via8_120x400_800H_721V_ARRAY_2x1 PGVIA
   VIA   v8    0.8 0.8            1.201 1.201         via8_120x400_800H_1201V_ARRAY_3x1 PGVIA
   VIA   v8    0.8 0.8            2.401 2.401         via8_120x400_800H_2401V_ARRAY_6x1 PGVIA
   VIA   v8    0.9 0.9            0.721 0.721         via8_120x400_900H_721V_ARRAY_2x1 PGVIA
   VIA   v8    0.9 0.9            1.201 1.201         via8_120x400_900H_1201V_ARRAY_3x1 PGVIA
   VIA   v8    0.9 0.9            2.401 2.401         via8_120x400_900H_2401V_ARRAY_6x1 PGVIA
   VIA   vmz   0.54 0.721         0.54 0.54           VMZ_120X400_540V_540H
   VIA   vmz   0.54 0.721         0.721 1.08          VMZ_120X400_540V_721H
   VIA   vmz   0.54 0.721         1.201 1.201         VMZ_120X400_540V_1201H
   VIA   vmz   0.54 0.54          2.13 2.13           VMZ_120x400_540V_2130H_ARRAY_1x2
   VIA   vmz   0.54 0.721         2.401 2.401         VMZ_120X400_540V_2401H
   VIA   vmz   0.54 0.54          3.98 3.98           VMZ_120x400_540V_3980H_ARRAY_1x3
   VIA   vmz   0.721 0.721        2.13 2.13           VMZ_120x400_721V_2130H_ARRAY_1x2
   VIA   vmz   0.721 0.721        3.98 3.98           VMZ_120x400_721V_3980H_ARRAY_1x3
   VIA   vmz   1.201 1.201        0.54 0.54           VMZ_120x400_1201V_540H_ARRAY_2x1
   VIA   vmz   1.201 1.201        0.721 0.721         VMZ_120x400_1201V_721H_ARRAY_2x1
   VIA   vmz   1.201 1.201        1.08 1.08           VMZ_120x400_1201V_1080H_ARRAY_2x1
   VIA   vmz   1.201 1.201        1.201 1.201         VMZ_120x400_1201V_1201H_ARRAY_2x1
   VIA   vmz   1.201 1.201        2.13 2.13           VMZ_120x400_1201V_2130H_ARRAY_2x2
   VIA   vmz   1.201 1.201        2.401 2.401         VMZ_120x400_1201V_2401H_ARRAY_2x1
   VIA   vmz   1.201 1.201        3.98 3.98           VMZ_120x400_1201V_3980H_ARRAY_2x3
   VIA   vmz   2.401 2.401        0.54 0.54           VMZ_120x400_2401V_540H_ARRAY_6x1
   VIA   vmz   2.401 2.401        0.721 0.721         VMZ_120x400_2401V_721H_ARRAY_6x1
   VIA   vmz   2.401 2.401        1.08 1.08           VMZ_120x400_2401V_1080H_ARRAY_6x1
   VIA   vmz   2.401 2.401        1.201 1.201         VMZ_120x400_2401V_1201H_ARRAY_6x1
   VIA   vmz   2.401 2.401        2.13 2.13           VMZ_120x400_2401V_2130H_ARRAY_6x2
   VIA   vmz   2.401 2.401        2.401 2.401         VMZ_120x400_2401V_2401H_ARRAY_6x1
   VIA   vmz   2.401 2.401        3.98 3.98           VMZ_120x400_2401V_3980H_ARRAY_6x3
   VIA   vmz   0.54 0.721         0.54 0.54           VMZ_120X400_540H_540V PGVIA
   VIA   vmz   0.54 1.201         0.721 1.08          VMZ_120X400_540H_721V PGVIA
   VIA   vmz   0.54 1.201         1.201 1.201         VMZ_120X400_540H_1201V PGVIA
   VIA   vmz   0.54 0.54          2.13 2.13           VMZ_120x400_540H_2130V_ARRAY_3x1 PGVIA
   VIA   vmz   0.54 1.201         2.401 2.401         VMZ_120X400_540H_2401V PGVIA
   VIA   vmz   0.54 0.54          3.98 3.98           VMZ_120x400_540H_3980V_ARRAY_5x1 PGVIA
   VIA   vmz   0.721 0.721        2.13 2.13           VMZ_120x400_721H_2130V_ARRAY_3x1 PGVIA
   VIA   vmz   0.721 0.721        3.98 3.98           VMZ_120x400_721H_3980V_ARRAY_5x1 PGVIA
   VIA   vmz   1.201 1.201        0.54 0.54           VMZ_120x400_1201H_540V_ARRAY_1x2 PGVIA
   VIA   vmz   1.201 1.201        2.13 2.13           VMZ_120x400_1201H_2130V_ARRAY_3x1 PGVIA
   VIA   vmz   1.201 1.201        3.98 3.98           VMZ_120x400_1201H_3980V_ARRAY_5x1 PGVIA
   VIA   vmz   2.401 2.401        0.54 0.54           VMZ_120x400_2401H_540V_ARRAY_1x3 PGVIA
   VIA   vmz   2.401 2.401        0.721 0.721         VMZ_120x400_2401H_721V_ARRAY_1x3 PGVIA
   VIA   vmz   2.401 2.401        1.08 1.08           VMZ_120x400_2401H_1080V_ARRAY_1x3 PGVIA
   VIA   vmz   2.401 2.401        1.201 1.201         VMZ_120x400_2401H_1201V_ARRAY_1x3 PGVIA
   VIA   vmz   2.401 2.401        2.13 2.13           VMZ_120x400_2401H_2130V_ARRAY_3x3 PGVIA
   VIA   vmz   2.401 2.401        2.401 2.401         VMZ_120x400_2401H_2401V_ARRAY_1x3 PGVIA
   VIA   vmz   2.401 2.401        3.98 3.98           VMZ_120x400_2401H_3980V_ARRAY_5x3 PGVIA
   VIA   vmz   0.54 0.721         0.54 0.54           VMZ_120X400_540H_540H PGVIA
   VIA   vmz   0.54 0.54          0.721 0.721         VMZ_120x400_540H_721V_ARRAY_2x1 PGVIA
   VIA   vmz   0.54 0.54          1.08 1.08           VMZ_120x400_540H_1080V_ARRAY_3x1 PGVIA
   VIA   vmz   0.54 0.54          1.201 1.201         VMZ_120x400_540H_1201V_ARRAY_3x1 PGVIA
   VIA   vmz   0.54 0.54          2.13 2.13           VMZ_120x400_540H_2130V_ARRAY_5x1 PGVIA
   VIA   vmz   0.54 0.54          2.401 2.401         VMZ_120x400_540H_2401V_ARRAY_6x1 PGVIA
   VIA   vmz   0.54 0.54          3.98 3.98           VMZ_120x400_540H_3980V_ARRAY_10x1 PGVIA
   VIA   vmz   0.721 0.721        0.721 0.721         VMZ_120x400_721H_721V_ARRAY_2x1 PGVIA
   VIA   vmz   0.721 0.721        1.08 1.08           VMZ_120x400_721H_1080V_ARRAY_3x1 PGVIA
   VIA   vmz   0.721 0.721        1.201 1.201         VMZ_120x400_721H_1201V_ARRAY_3x1 PGVIA
   VIA   vmz   0.721 0.721        2.13 2.13           VMZ_120x400_721H_2130V_ARRAY_5x1 PGVIA
   VIA   vmz   0.721 0.721        2.401 2.401         VMZ_120x400_721H_2401V_ARRAY_6x1 PGVIA
   VIA   vmz   0.721 0.721        3.98 3.98           VMZ_120x400_721H_3980V_ARRAY_10x1 PGVIA
   VIA   vmz   1.201 1.201        0.721 0.721         VMZ_120x400_1201H_721V_ARRAY_2x1 PGVIA
   VIA   vmz   1.201 1.201        1.08 1.08           VMZ_120x400_1201H_1080V_ARRAY_3x1 PGVIA
   VIA   vmz   1.201 1.201        1.201 1.201         VMZ_120x400_1201H_1201V_ARRAY_3x1 PGVIA
   VIA   vmz   1.201 1.201        2.13 2.13           VMZ_120x400_1201H_2130V_ARRAY_5x1 PGVIA
   VIA   vmz   1.201 1.201        2.401 2.401         VMZ_120x400_1201H_2401V_ARRAY_6x1 PGVIA
   VIA   vmz   1.201 1.201        3.98 3.98           VMZ_120x400_1201H_3980V_ARRAY_10x1 PGVIA
   VIA   vmz   2.401 2.401        0.721 0.721         VMZ_120x400_2401H_721V_ARRAY_2x3 PGVIA
   VIA   vmz   2.401 2.401        1.08 1.08           VMZ_120x400_2401H_1080V_ARRAY_3x3 PGVIA
   VIA   vmz   2.401 2.401        1.201 1.201         VMZ_120x400_2401H_1201V_ARRAY_3x2 PGVIA
   VIA   vmz   2.401 2.401        2.13 2.13           VMZ_120x400_2401H_2130V_ARRAY_5x2 PGVIA
   VIA   vmz   2.401 2.401        2.401 2.401         VMZ_120x400_2401H_2401V_ARRAY_6x1 PGVIA
   VIA   vmz   2.401 2.401        3.98 3.98           VMZ_120x400_2401H_3980V_ARRAY_10x1 PGVIA
   VIA   vmz   0.54 0.721         0.54 0.54           VMZ_120X400_540V_540V PGVIA
   VIA   vmz   0.54 0.721         0.721 1.08          VMZ_120X400_540V_721V PGVIA
   VIA   vmz   0.54 1.201         1.201 1.201         VMZ_120X400_540V_1201V PGVIA
   VIA   vmz   0.54 0.54          2.13 2.13           VMZ_120x400_540V_2130H_ARRAY_1x3 PGVIA
   VIA   vmz   0.54 0.54          2.401 2.401         VMZ_120x400_540V_2401H_ARRAY_1x3 PGVIA
   VIA   vmz   0.54 0.54          3.98 3.98           VMZ_120x400_540V_3980H_ARRAY_1x6 PGVIA
   VIA   vmz   0.721 0.721        2.13 2.13           VMZ_120x400_721V_2130H_ARRAY_1x3 PGVIA
   VIA   vmz   0.721 0.721        2.401 2.401         VMZ_120x400_721V_2401H_ARRAY_1x3 PGVIA
   VIA   vmz   0.721 0.721        3.98 3.98           VMZ_120x400_721V_3980H_ARRAY_1x6 PGVIA
   VIA   vmz   1.201 1.201        2.13 2.13           VMZ_120x400_1201V_2130H_ARRAY_1x3 PGVIA
   VIA   vmz   1.201 1.201        2.401 2.401         VMZ_120x400_1201V_2401H_ARRAY_2x3 PGVIA
   VIA   vmz   1.201 1.201        3.98 3.98           VMZ_120x400_1201V_3980H_ARRAY_2x6 PGVIA
   VIA   vmz   2.401 2.401        0.721 0.721         VMZ_120x400_2401V_721H_ARRAY_5x1 PGVIA
   VIA   vmz   2.401 2.401        1.08 1.08           VMZ_120x400_2401V_1080H_ARRAY_5x1 PGVIA
   VIA   vmz   2.401 2.401        1.201 1.201         VMZ_120x400_2401V_1201H_ARRAY_4x1 PGVIA
   VIA   vmz   2.401 2.401        2.13 2.13           VMZ_120x400_2401V_2130H_ARRAY_4x3 PGVIA
   VIA   vmz   2.401 2.401        2.401 2.401         VMZ_120x400_2401V_2401H_ARRAY_1x3 PGVIA
   VIA   vmz   2.401 2.401        3.98 3.98           VMZ_120x400_2401V_3980H_ARRAY_1x6 PGVIA
   VIA   gv0   0.54 7.000         1.0 4.0             GV0_1850X800_1080H_3050V
   VIA   gv0   0.54 7.000         4.00 8.60           GV0_3700X800_1080H_4900V
   VIA   gv0   0.54 7.000         8.6 12.0            GV0_7400X800_1080H_8600V
   VIA   gv0   0.54 7.000         1.0 4.0             GV0_1850X800_1080H_3050V PGVIA
   VIA   gv0   0.54 7.000         4.00 8.60           GV0_3700X800_1080H_4900V PGVIA
   VIA   gv0   0.54 7.000         8.6 12.0            GV0_7400X800_1080H_8600V PGVIA
   VIA   gv0   0.54 7.000         1.0 4.0             GV0_800X1850_1080V_3050H PGVIA
   VIA   gv0   0.54 7.000         4.00 8.60           GV0_800X3700_1080V_4900H PGVIA
   VIA   gv0   0.54 7.000         8.6 12.0            GV0_800X7400_1080V_8600H PGVIA
   VIA   gv0   0.54 7.00          1.0 12.0            GV0_7400X800_1080H_2000H PGVIA
   VIA   gv0   0.54 7.00          1.0 12.0            GV0_800X7400_1080V_2000V PGVIA
   ;
 " ;
END PROPERTYDEFINITIONS




#################################################
# Site Definitions
#################################################
SITE core
 CLASS CORE ;
 SIZE 0.1080 BY 0.6300 ;
 SYMMETRY X Y ;
END core

SITE core2h
 CLASS CORE ;
 SIZE 0.1080 BY 1.2600 ;
 SYMMETRY X Y ;
END core2h

SITE bonuscore
 CLASS CORE ;
 SIZE 0.4320 BY 0.6300 ;
 SYMMETRY X Y ;
END bonuscore


END LIBRARY
