module ring_terminator_n1 ();
endmodule

module sup1v8_n1 ();
endmodule