VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO uni_2x2sub4x4_gpio_top_lef_LEFT_SIDE
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN uni_2x2sub4x4_gpio_top_lef_LEFT_SIDE 0 0 ;
  SIZE 623.808 BY 911.933 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN dq[40]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 616.446 776.48 616.626 778.68 ;
    END
  END dq[40]
  PIN dq[41]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 473.886 776.48 474.066 778.68 ;
    END
  END dq[41]
  PIN dq[42]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 612.126 776.48 612.306 778.68 ;
    END
  END dq[42]
  PIN dq[43]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 478.206 776.48 478.386 778.68 ;
    END
  END dq[43]
  PIN dq[44]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 549.846 776.48 550.026 778.68 ;
    END
  END dq[44]
  PIN dq[45]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 536.166 776.48 536.346 778.68 ;
    END
  END dq[45]
  PIN dq[46]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 581.886 776.48 582.066 778.68 ;
    END
  END dq[46]
  PIN dq[47]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 503.046 776.48 503.226 778.68 ;
    END
  END dq[47]
  PIN dq[48]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 460.494 776.48 460.674 778.68 ;
    END
  END dq[48]
  PIN dq[49]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 317.934 776.48 318.114 778.68 ;
    END
  END dq[49]
  PIN dq[50]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 456.174 776.48 456.354 778.68 ;
    END
  END dq[50]
  PIN dq[51]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 322.254 776.48 322.434 778.68 ;
    END
  END dq[51]
  PIN dq[52]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 393.894 776.48 394.074 778.68 ;
    END
  END dq[52]
  PIN dq[53]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 380.214 776.48 380.394 778.68 ;
    END
  END dq[53]
  PIN dq[54]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 425.934 776.48 426.114 778.68 ;
    END
  END dq[54]
  PIN dq[55]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 347.094 776.48 347.274 778.68 ;
    END
  END dq[55]
  PIN dq[56]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 304.542 776.48 304.722 778.68 ;
    END
  END dq[56]
  PIN dq[57]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 161.982 776.48 162.162 778.68 ;
    END
  END dq[57]
  PIN dq[58]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 300.222 776.48 300.402 778.68 ;
    END
  END dq[58]
  PIN dq[59]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 166.302 776.48 166.482 778.68 ;
    END
  END dq[59]
  PIN dq[60]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 237.942 776.48 238.122 778.68 ;
    END
  END dq[60]
  PIN dq[61]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 224.262 776.48 224.442 778.68 ;
    END
  END dq[61]
  PIN dq[62]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 269.982 776.48 270.162 778.68 ;
    END
  END dq[62]
  PIN dq[63]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 191.142 776.48 191.322 778.68 ;
    END
  END dq[63]
  PIN dq[64]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 148.59 776.48 148.77 778.68 ;
    END
  END dq[64]
  PIN dq[65]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 6.03 776.48 6.21 778.68 ;
    END
  END dq[65]
  PIN dq[66]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 144.27 776.48 144.45 778.68 ;
    END
  END dq[66]
  PIN dq[67]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 10.35 776.48 10.53 778.68 ;
    END
  END dq[67]
  PIN dq[68]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 81.99 776.48 82.17 778.68 ;
    END
  END dq[68]
  PIN dq[69]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 68.31 776.48 68.49 778.68 ;
    END
  END dq[69]
  PIN dq[70]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 114.03 776.48 114.21 778.68 ;
    END
  END dq[70]
  PIN dq[71]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 35.19 776.48 35.37 778.68 ;
    END
  END dq[71]
  PIN drv0[5]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 622.926 776.48 623.106 778.68 ;
    END
  END drv0[5]
  PIN drv0[6]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 466.974 776.48 467.154 778.68 ;
    END
  END drv0[6]
  PIN drv0[7]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 311.022 776.48 311.202 778.68 ;
    END
  END drv0[7]
  PIN drv0[8]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 155.07 776.48 155.25 778.68 ;
    END
  END drv0[8]
  PIN drv1[5]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 621.846 776.48 622.026 778.68 ;
    END
  END drv1[5]
  PIN drv1[6]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 465.894 776.48 466.074 778.68 ;
    END
  END drv1[6]
  PIN drv1[7]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 309.942 776.48 310.122 778.68 ;
    END
  END drv1[7]
  PIN drv1[8]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 153.99 776.48 154.17 778.68 ;
    END
  END drv1[8]
  PIN drv2[5]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 620.766 776.48 620.946 778.68 ;
    END
  END drv2[5]
  PIN drv2[6]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 464.814 776.48 464.994 778.68 ;
    END
  END drv2[6]
  PIN drv2[7]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 308.862 776.48 309.042 778.68 ;
    END
  END drv2[7]
  PIN drv2[8]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 152.91 776.48 153.09 778.68 ;
    END
  END drv2[8]
  PIN enabq[40]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 615.366 776.48 615.546 778.68 ;
    END
  END enabq[40]
  PIN enabq[41]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 474.966 776.48 475.146 778.68 ;
    END
  END enabq[41]
  PIN enabq[42]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 613.206 776.48 613.386 778.68 ;
    END
  END enabq[42]
  PIN enabq[43]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 477.126 776.48 477.306 778.68 ;
    END
  END enabq[43]
  PIN enabq[44]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 556.326 776.48 556.506 778.68 ;
    END
  END enabq[44]
  PIN enabq[45]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 542.646 776.48 542.826 778.68 ;
    END
  END enabq[45]
  PIN enabq[46]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 588.366 776.48 588.546 778.68 ;
    END
  END enabq[46]
  PIN enabq[47]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 509.526 776.48 509.706 778.68 ;
    END
  END enabq[47]
  PIN enabq[48]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 459.414 776.48 459.594 778.68 ;
    END
  END enabq[48]
  PIN enabq[49]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 319.014 776.48 319.194 778.68 ;
    END
  END enabq[49]
  PIN enabq[50]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 457.254 776.48 457.434 778.68 ;
    END
  END enabq[50]
  PIN enabq[51]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 321.174 776.48 321.354 778.68 ;
    END
  END enabq[51]
  PIN enabq[52]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 400.374 776.48 400.554 778.68 ;
    END
  END enabq[52]
  PIN enabq[53]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 386.694 776.48 386.874 778.68 ;
    END
  END enabq[53]
  PIN enabq[54]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 432.414 776.48 432.594 778.68 ;
    END
  END enabq[54]
  PIN enabq[55]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 353.574 776.48 353.754 778.68 ;
    END
  END enabq[55]
  PIN enabq[56]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 303.462 776.48 303.642 778.68 ;
    END
  END enabq[56]
  PIN enabq[57]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 163.062 776.48 163.242 778.68 ;
    END
  END enabq[57]
  PIN enabq[58]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 301.302 776.48 301.482 778.68 ;
    END
  END enabq[58]
  PIN enabq[59]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 165.222 776.48 165.402 778.68 ;
    END
  END enabq[59]
  PIN enabq[60]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 244.422 776.48 244.602 778.68 ;
    END
  END enabq[60]
  PIN enabq[61]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 230.742 776.48 230.922 778.68 ;
    END
  END enabq[61]
  PIN enabq[62]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 276.462 776.48 276.642 778.68 ;
    END
  END enabq[62]
  PIN enabq[63]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 197.622 776.48 197.802 778.68 ;
    END
  END enabq[63]
  PIN enabq[64]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 147.51 776.48 147.69 778.68 ;
    END
  END enabq[64]
  PIN enabq[65]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 7.11 776.48 7.29 778.68 ;
    END
  END enabq[65]
  PIN enabq[66]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 145.35 776.48 145.53 778.68 ;
    END
  END enabq[66]
  PIN enabq[67]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 9.27 776.48 9.45 778.68 ;
    END
  END enabq[67]
  PIN enabq[68]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 88.47 776.48 88.65 778.68 ;
    END
  END enabq[68]
  PIN enabq[69]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 74.79 776.48 74.97 778.68 ;
    END
  END enabq[69]
  PIN enabq[70]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 120.51 776.48 120.69 778.68 ;
    END
  END enabq[70]
  PIN enabq[71]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 41.67 776.48 41.85 778.68 ;
    END
  END enabq[71]
  PIN enq[40]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 614.646 776.48 614.826 778.68 ;
    END
  END enq[40]
  PIN enq[41]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 475.686 776.48 475.866 778.68 ;
    END
  END enq[41]
  PIN enq[42]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 613.926 776.48 614.106 778.68 ;
    END
  END enq[42]
  PIN enq[43]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 476.406 776.48 476.586 778.68 ;
    END
  END enq[43]
  PIN enq[44]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 554.166 776.48 554.346 778.68 ;
    END
  END enq[44]
  PIN enq[45]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 540.486 776.48 540.666 778.68 ;
    END
  END enq[45]
  PIN enq[46]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 586.206 776.48 586.386 778.68 ;
    END
  END enq[46]
  PIN enq[47]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 507.366 776.48 507.546 778.68 ;
    END
  END enq[47]
  PIN enq[48]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 458.694 776.48 458.874 778.68 ;
    END
  END enq[48]
  PIN enq[49]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 319.734 776.48 319.914 778.68 ;
    END
  END enq[49]
  PIN enq[50]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 457.974 776.48 458.154 778.68 ;
    END
  END enq[50]
  PIN enq[51]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 320.454 776.48 320.634 778.68 ;
    END
  END enq[51]
  PIN enq[52]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 398.214 776.48 398.394 778.68 ;
    END
  END enq[52]
  PIN enq[53]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 384.534 776.48 384.714 778.68 ;
    END
  END enq[53]
  PIN enq[54]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 430.254 776.48 430.434 778.68 ;
    END
  END enq[54]
  PIN enq[55]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 351.414 776.48 351.594 778.68 ;
    END
  END enq[55]
  PIN enq[56]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 302.742 776.48 302.922 778.68 ;
    END
  END enq[56]
  PIN enq[57]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 163.782 776.48 163.962 778.68 ;
    END
  END enq[57]
  PIN enq[58]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 302.022 776.48 302.202 778.68 ;
    END
  END enq[58]
  PIN enq[59]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 164.502 776.48 164.682 778.68 ;
    END
  END enq[59]
  PIN enq[60]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 242.262 776.48 242.442 778.68 ;
    END
  END enq[60]
  PIN enq[61]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 228.582 776.48 228.762 778.68 ;
    END
  END enq[61]
  PIN enq[62]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 274.302 776.48 274.482 778.68 ;
    END
  END enq[62]
  PIN enq[63]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 195.462 776.48 195.642 778.68 ;
    END
  END enq[63]
  PIN enq[64]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 146.79 776.48 146.97 778.68 ;
    END
  END enq[64]
  PIN enq[65]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 7.83 776.48 8.01 778.68 ;
    END
  END enq[65]
  PIN enq[66]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 146.07 776.48 146.25 778.68 ;
    END
  END enq[66]
  PIN enq[67]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 8.55 776.48 8.73 778.68 ;
    END
  END enq[67]
  PIN enq[68]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 86.31 776.48 86.49 778.68 ;
    END
  END enq[68]
  PIN enq[69]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 72.63 776.48 72.81 778.68 ;
    END
  END enq[69]
  PIN enq[70]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 118.35 776.48 118.53 778.68 ;
    END
  END enq[70]
  PIN enq[71]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 39.51 776.48 39.69 778.68 ;
    END
  END enq[71]
  PIN outi[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 617.526 776.48 617.706 778.68 ;
    END
  END outi[40]
  PIN outi[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 472.806 776.48 472.986 778.68 ;
    END
  END outi[41]
  PIN outi[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 611.046 776.48 611.226 778.68 ;
    END
  END outi[42]
  PIN outi[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 479.286 776.48 479.466 778.68 ;
    END
  END outi[43]
  PIN outi[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 552.006 776.48 552.186 778.68 ;
    END
  END outi[44]
  PIN outi[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 538.326 776.48 538.506 778.68 ;
    END
  END outi[45]
  PIN outi[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 584.046 776.48 584.226 778.68 ;
    END
  END outi[46]
  PIN outi[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 505.206 776.48 505.386 778.68 ;
    END
  END outi[47]
  PIN outi[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 461.574 776.48 461.754 778.68 ;
    END
  END outi[48]
  PIN outi[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 316.854 776.48 317.034 778.68 ;
    END
  END outi[49]
  PIN outi[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 455.094 776.48 455.274 778.68 ;
    END
  END outi[50]
  PIN outi[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 323.334 776.48 323.514 778.68 ;
    END
  END outi[51]
  PIN outi[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 396.054 776.48 396.234 778.68 ;
    END
  END outi[52]
  PIN outi[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 382.374 776.48 382.554 778.68 ;
    END
  END outi[53]
  PIN outi[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 428.094 776.48 428.274 778.68 ;
    END
  END outi[54]
  PIN outi[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 349.254 776.48 349.434 778.68 ;
    END
  END outi[55]
  PIN outi[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 305.622 776.48 305.802 778.68 ;
    END
  END outi[56]
  PIN outi[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 160.902 776.48 161.082 778.68 ;
    END
  END outi[57]
  PIN outi[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 299.142 776.48 299.322 778.68 ;
    END
  END outi[58]
  PIN outi[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 167.382 776.48 167.562 778.68 ;
    END
  END outi[59]
  PIN outi[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 240.102 776.48 240.282 778.68 ;
    END
  END outi[60]
  PIN outi[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 226.422 776.48 226.602 778.68 ;
    END
  END outi[61]
  PIN outi[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 272.142 776.48 272.322 778.68 ;
    END
  END outi[62]
  PIN outi[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 193.302 776.48 193.482 778.68 ;
    END
  END outi[63]
  PIN outi[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 149.67 776.48 149.85 778.68 ;
    END
  END outi[64]
  PIN outi[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 4.95 776.48 5.13 778.68 ;
    END
  END outi[65]
  PIN outi[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 143.19 776.48 143.37 778.68 ;
    END
  END outi[66]
  PIN outi[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 11.43 776.48 11.61 778.68 ;
    END
  END outi[67]
  PIN outi[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 84.15 776.48 84.33 778.68 ;
    END
  END outi[68]
  PIN outi[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 70.47 776.48 70.65 778.68 ;
    END
  END outi[69]
  PIN outi[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 116.19 776.48 116.37 778.68 ;
    END
  END outi[70]
  PIN outi[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m7 ;
        RECT 37.35 776.48 37.53 778.68 ;
    END
  END outi[71]
  PIN pd[5]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 619.686 776.48 619.866 778.68 ;
    END
  END pd[5]
  PIN pd[6]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 463.734 776.48 463.914 778.68 ;
    END
  END pd[6]
  PIN pd[7]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 307.782 776.48 307.962 778.68 ;
    END
  END pd[7]
  PIN pd[8]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 151.83 776.48 152.01 778.68 ;
    END
  END pd[8]
  PIN ppen[5]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 469.566 776.48 469.746 778.68 ;
    END
  END ppen[5]
  PIN ppen[6]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 313.614 776.48 313.794 778.68 ;
    END
  END ppen[6]
  PIN ppen[7]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 157.662 776.48 157.842 778.68 ;
    END
  END ppen[7]
  PIN ppen[8]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 1.71 776.48 1.89 778.68 ;
    END
  END ppen[8]
  PIN prg_slew[5]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 468.486 776.48 468.666 778.68 ;
    END
  END prg_slew[5]
  PIN prg_slew[6]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 312.534 776.48 312.714 778.68 ;
    END
  END prg_slew[6]
  PIN prg_slew[7]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 156.582 776.48 156.762 778.68 ;
    END
  END prg_slew[7]
  PIN prg_slew[8]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 0.63 776.48 0.81 778.68 ;
    END
  END prg_slew[8]
  PIN puq[5]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 618.606 776.48 618.786 778.68 ;
    END
  END puq[5]
  PIN puq[6]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 462.654 776.48 462.834 778.68 ;
    END
  END puq[6]
  PIN puq[7]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 306.702 776.48 306.882 778.68 ;
    END
  END puq[7]
  PIN puq[8]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 150.75 776.48 150.93 778.68 ;
    END
  END puq[8]
  PIN pwrup_pull_en[5]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 470.646 776.48 470.826 778.68 ;
    END
  END pwrup_pull_en[5]
  PIN pwrup_pull_en[6]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 314.694 776.48 314.874 778.68 ;
    END
  END pwrup_pull_en[6]
  PIN pwrup_pull_en[7]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 158.742 776.48 158.922 778.68 ;
    END
  END pwrup_pull_en[7]
  PIN pwrup_pull_en[8]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 2.79 776.48 2.97 778.68 ;
    END
  END pwrup_pull_en[8]
  PIN pwrupzhl[5]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 471.726 776.48 471.906 778.68 ;
    END
  END pwrupzhl[5]
  PIN pwrupzhl[6]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 315.774 776.48 315.954 778.68 ;
    END
  END pwrupzhl[6]
  PIN pwrupzhl[7]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 159.822 776.48 160.002 778.68 ;
    END
  END pwrupzhl[7]
  PIN pwrupzhl[8]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m7 ;
        RECT 3.87 776.48 4.05 778.68 ;
    END
  END pwrupzhl[8]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER gmz ;
        RECT 327.959 783.5175 330.409 910.004 ;
    END
    PORT
      LAYER gmz ;
        RECT 604.871 783.5175 607.321 910.004 ;
        RECT 587.591 783.5175 590.041 910.004 ;
        RECT 570.311 783.5175 572.761 910.004 ;
        RECT 553.031 783.5175 555.481 910.004 ;
        RECT 535.751 783.5175 538.201 910.004 ;
        RECT 518.471 783.5175 520.921 910.004 ;
        RECT 501.191 783.5175 503.641 910.004 ;
        RECT 483.911 783.5175 486.361 910.004 ;
        RECT 448.919 783.5175 451.369 910.004 ;
        RECT 431.639 783.5175 434.089 910.004 ;
        RECT 414.359 783.5175 416.809 910.004 ;
        RECT 397.079 783.5175 399.529 910.004 ;
        RECT 379.799 783.5175 382.249 910.004 ;
        RECT 362.519 783.5175 364.969 910.004 ;
        RECT 345.239 783.5175 347.689 910.004 ;
        RECT 292.967 783.5175 295.417 910.004 ;
        RECT 275.687 783.5175 278.137 910.004 ;
        RECT 258.407 783.5175 260.857 910.004 ;
        RECT 241.127 783.5175 243.577 910.004 ;
        RECT 223.847 783.5175 226.297 910.004 ;
        RECT 206.567 783.5175 209.017 910.004 ;
        RECT 189.287 783.5175 191.737 910.004 ;
        RECT 172.007 783.5175 174.457 910.004 ;
        RECT 137.015 783.5175 139.465 910.004 ;
        RECT 119.735 783.5175 122.185 910.004 ;
        RECT 102.455 783.5175 104.905 910.004 ;
        RECT 85.175 783.5175 87.625 910.004 ;
        RECT 67.895 783.5175 70.345 910.004 ;
        RECT 50.615 783.5175 53.065 910.004 ;
        RECT 33.335 783.5175 35.785 910.004 ;
        RECT 16.055 783.5175 18.505 910.004 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER gmz ;
        RECT 613.511 783.5175 615.961 910.004 ;
        RECT 596.231 783.5175 598.681 910.004 ;
        RECT 578.951 783.5175 581.401 910.004 ;
        RECT 561.671 783.5175 564.121 910.004 ;
        RECT 544.391 783.5175 546.841 910.004 ;
        RECT 527.111 783.5175 529.561 910.004 ;
        RECT 509.831 783.5175 512.281 910.004 ;
        RECT 492.551 783.5175 495.001 910.004 ;
        RECT 475.271 783.5175 477.721 910.004 ;
        RECT 457.559 783.5175 460.009 910.004 ;
        RECT 440.279 783.5175 442.729 910.004 ;
        RECT 422.999 783.5175 425.449 910.004 ;
        RECT 405.719 783.5175 408.169 910.004 ;
        RECT 388.439 783.5175 390.889 910.004 ;
        RECT 371.159 783.5175 373.609 910.004 ;
        RECT 353.879 783.5175 356.329 910.004 ;
        RECT 336.599 783.5175 339.049 910.004 ;
        RECT 319.319 783.5175 321.769 910.004 ;
        RECT 301.607 783.5175 304.057 910.004 ;
        RECT 284.327 783.5175 286.777 910.004 ;
        RECT 267.047 783.5175 269.497 910.004 ;
        RECT 249.767 783.5175 252.217 910.004 ;
        RECT 232.487 783.5175 234.937 910.004 ;
        RECT 215.207 783.5175 217.657 910.004 ;
        RECT 197.927 783.5175 200.377 910.004 ;
        RECT 180.647 783.5175 183.097 910.004 ;
        RECT 163.367 783.5175 165.817 910.004 ;
        RECT 145.655 783.5175 148.105 910.004 ;
        RECT 128.375 783.5175 130.825 910.004 ;
        RECT 111.095 783.5175 113.545 910.004 ;
        RECT 93.815 783.5175 96.265 910.004 ;
        RECT 76.535 783.5175 78.985 910.004 ;
        RECT 59.255 783.5175 61.705 910.004 ;
        RECT 41.975 783.5175 44.425 910.004 ;
        RECT 24.695 783.5175 27.145 910.004 ;
        RECT 7.415 783.5175 9.865 910.004 ;
    END
  END vss
  OBS
    LAYER m1 SPACING 0.04 ;
      RECT 0 0 623.808 911.933 ;
    LAYER m5 SPACING 0.046 ;
      RECT 0 0 623.808 911.933 ;
    LAYER m2 SPACING 0.046 ;
      RECT 0 0 623.808 911.933 ;
    LAYER m3 SPACING 0.046 ;
      RECT 0 0 623.808 911.933 ;
    LAYER m4 SPACING 0.046 ;
      RECT 0 0 623.808 911.933 ;
    LAYER m8 SPACING 0.18 ;
      RECT 0 779.56 623.808 911.933 ;
      RECT 589.426 0 610.166 911.933 ;
      RECT 587.266 0 587.486 911.933 ;
      RECT 585.106 0 585.326 911.933 ;
      RECT 582.946 0 583.166 911.933 ;
      RECT 557.386 0 581.006 911.933 ;
      RECT 555.226 0 555.446 911.933 ;
      RECT 553.066 0 553.286 911.933 ;
      RECT 550.906 0 551.126 911.933 ;
      RECT 543.706 0 548.966 911.933 ;
      RECT 541.546 0 541.766 911.933 ;
      RECT 539.386 0 539.606 911.933 ;
      RECT 537.226 0 537.446 911.933 ;
      RECT 510.586 0 535.286 911.933 ;
      RECT 508.426 0 508.646 911.933 ;
      RECT 506.266 0 506.486 911.933 ;
      RECT 504.106 0 504.326 911.933 ;
      RECT 480.346 0 502.166 911.933 ;
      RECT 433.474 0 454.214 911.933 ;
      RECT 431.314 0 431.534 911.933 ;
      RECT 429.154 0 429.374 911.933 ;
      RECT 426.994 0 427.214 911.933 ;
      RECT 401.434 0 425.054 911.933 ;
      RECT 399.274 0 399.494 911.933 ;
      RECT 397.114 0 397.334 911.933 ;
      RECT 394.954 0 395.174 911.933 ;
      RECT 387.754 0 393.014 911.933 ;
      RECT 385.594 0 385.814 911.933 ;
      RECT 383.434 0 383.654 911.933 ;
      RECT 381.274 0 381.494 911.933 ;
      RECT 354.634 0 379.334 911.933 ;
      RECT 352.474 0 352.694 911.933 ;
      RECT 350.314 0 350.534 911.933 ;
      RECT 348.154 0 348.374 911.933 ;
      RECT 324.394 0 346.214 911.933 ;
      RECT 277.522 0 298.262 911.933 ;
      RECT 275.362 0 275.582 911.933 ;
      RECT 273.202 0 273.422 911.933 ;
      RECT 271.042 0 271.262 911.933 ;
      RECT 245.482 0 269.102 911.933 ;
      RECT 243.322 0 243.542 911.933 ;
      RECT 241.162 0 241.382 911.933 ;
      RECT 239.002 0 239.222 911.933 ;
      RECT 231.802 0 237.062 911.933 ;
      RECT 229.642 0 229.862 911.933 ;
      RECT 227.482 0 227.702 911.933 ;
      RECT 225.322 0 225.542 911.933 ;
      RECT 198.682 0 223.382 911.933 ;
      RECT 196.522 0 196.742 911.933 ;
      RECT 194.362 0 194.582 911.933 ;
      RECT 192.202 0 192.422 911.933 ;
      RECT 168.442 0 190.262 911.933 ;
      RECT 121.57 0 142.31 911.933 ;
      RECT 119.41 0 119.63 911.933 ;
      RECT 117.25 0 117.47 911.933 ;
      RECT 115.09 0 115.31 911.933 ;
      RECT 89.53 0 113.15 911.933 ;
      RECT 87.37 0 87.59 911.933 ;
      RECT 85.21 0 85.43 911.933 ;
      RECT 83.05 0 83.27 911.933 ;
      RECT 75.85 0 81.11 911.933 ;
      RECT 73.69 0 73.91 911.933 ;
      RECT 71.53 0 71.75 911.933 ;
      RECT 69.37 0 69.59 911.933 ;
      RECT 42.73 0 67.43 911.933 ;
      RECT 40.57 0 40.79 911.933 ;
      RECT 38.41 0 38.63 911.933 ;
      RECT 36.25 0 36.47 911.933 ;
      RECT 12.49 0 34.31 911.933 ;
      RECT 0 0 623.808 775.6 ;
    LAYER m6 SPACING 0.046 ;
      RECT 0 0 623.808 911.933 ;
    LAYER m7 SPACING 0.18 ;
      RECT 0 779.1 623.808 911.933 ;
      RECT 623.526 0 623.808 911.933 ;
      RECT 588.966 0 610.626 911.933 ;
      RECT 586.806 0 587.946 911.933 ;
      RECT 584.646 0 585.786 911.933 ;
      RECT 582.486 0 583.626 911.933 ;
      RECT 556.926 0 581.466 911.933 ;
      RECT 554.766 0 555.906 911.933 ;
      RECT 552.606 0 553.746 911.933 ;
      RECT 550.446 0 551.586 911.933 ;
      RECT 543.246 0 549.426 911.933 ;
      RECT 541.086 0 542.226 911.933 ;
      RECT 538.926 0 540.066 911.933 ;
      RECT 536.766 0 537.906 911.933 ;
      RECT 510.126 0 535.746 911.933 ;
      RECT 507.966 0 509.106 911.933 ;
      RECT 505.806 0 506.946 911.933 ;
      RECT 503.646 0 504.786 911.933 ;
      RECT 479.886 0 502.626 911.933 ;
      RECT 467.574 0 468.066 911.933 ;
      RECT 433.014 0 454.674 911.933 ;
      RECT 430.854 0 431.994 911.933 ;
      RECT 428.694 0 429.834 911.933 ;
      RECT 426.534 0 427.674 911.933 ;
      RECT 400.974 0 425.514 911.933 ;
      RECT 398.814 0 399.954 911.933 ;
      RECT 396.654 0 397.794 911.933 ;
      RECT 394.494 0 395.634 911.933 ;
      RECT 387.294 0 393.474 911.933 ;
      RECT 385.134 0 386.274 911.933 ;
      RECT 382.974 0 384.114 911.933 ;
      RECT 380.814 0 381.954 911.933 ;
      RECT 354.174 0 379.794 911.933 ;
      RECT 352.014 0 353.154 911.933 ;
      RECT 349.854 0 350.994 911.933 ;
      RECT 347.694 0 348.834 911.933 ;
      RECT 323.934 0 346.674 911.933 ;
      RECT 311.622 0 312.114 911.933 ;
      RECT 277.062 0 298.722 911.933 ;
      RECT 274.902 0 276.042 911.933 ;
      RECT 272.742 0 273.882 911.933 ;
      RECT 270.582 0 271.722 911.933 ;
      RECT 245.022 0 269.562 911.933 ;
      RECT 242.862 0 244.002 911.933 ;
      RECT 240.702 0 241.842 911.933 ;
      RECT 238.542 0 239.682 911.933 ;
      RECT 231.342 0 237.522 911.933 ;
      RECT 229.182 0 230.322 911.933 ;
      RECT 227.022 0 228.162 911.933 ;
      RECT 224.862 0 226.002 911.933 ;
      RECT 198.222 0 223.842 911.933 ;
      RECT 196.062 0 197.202 911.933 ;
      RECT 193.902 0 195.042 911.933 ;
      RECT 191.742 0 192.882 911.933 ;
      RECT 167.982 0 190.722 911.933 ;
      RECT 155.67 0 156.162 911.933 ;
      RECT 121.11 0 142.77 911.933 ;
      RECT 118.95 0 120.09 911.933 ;
      RECT 116.79 0 117.93 911.933 ;
      RECT 114.63 0 115.77 911.933 ;
      RECT 89.07 0 113.61 911.933 ;
      RECT 86.91 0 88.05 911.933 ;
      RECT 84.75 0 85.89 911.933 ;
      RECT 82.59 0 83.73 911.933 ;
      RECT 75.39 0 81.57 911.933 ;
      RECT 73.23 0 74.37 911.933 ;
      RECT 71.07 0 72.21 911.933 ;
      RECT 68.91 0 70.05 911.933 ;
      RECT 42.27 0 67.89 911.933 ;
      RECT 40.11 0 41.25 911.933 ;
      RECT 37.95 0 39.09 911.933 ;
      RECT 35.79 0 36.93 911.933 ;
      RECT 12.03 0 34.77 911.933 ;
      RECT 0 0 0.21 911.933 ;
      RECT 0 0 623.808 776.06 ;
    LAYER c4 SPACING 49.3 ;
      RECT 0 0 623.808 911.933 ;
    LAYER c4emib SPACING 35 ;
      RECT 0 0 623.808 911.933 ;
    LAYER gm0 SPACING 0.54 ;
      RECT 0 910.644 623.808 911.933 ;
      RECT 616.601 0 623.808 911.933 ;
      RECT 607.961 0 612.871 911.933 ;
      RECT 599.321 0 604.231 911.933 ;
      RECT 590.681 0 595.591 911.933 ;
      RECT 582.041 0 586.951 911.933 ;
      RECT 573.401 0 578.311 911.933 ;
      RECT 564.761 0 569.671 911.933 ;
      RECT 556.121 0 561.031 911.933 ;
      RECT 547.481 0 552.391 911.933 ;
      RECT 538.841 0 543.751 911.933 ;
      RECT 530.201 0 535.111 911.933 ;
      RECT 521.561 0 526.471 911.933 ;
      RECT 512.921 0 517.831 911.933 ;
      RECT 504.281 0 509.191 911.933 ;
      RECT 495.641 0 500.551 911.933 ;
      RECT 487.001 0 491.911 911.933 ;
      RECT 478.361 0 483.271 911.933 ;
      RECT 460.649 0 474.631 911.933 ;
      RECT 452.009 0 456.919 911.933 ;
      RECT 443.369 0 448.279 911.933 ;
      RECT 434.729 0 439.639 911.933 ;
      RECT 426.089 0 430.999 911.933 ;
      RECT 417.449 0 422.359 911.933 ;
      RECT 408.809 0 413.719 911.933 ;
      RECT 400.169 0 405.079 911.933 ;
      RECT 391.529 0 396.439 911.933 ;
      RECT 382.889 0 387.799 911.933 ;
      RECT 374.249 0 379.159 911.933 ;
      RECT 365.609 0 370.519 911.933 ;
      RECT 356.969 0 361.879 911.933 ;
      RECT 348.329 0 353.239 911.933 ;
      RECT 339.689 0 344.599 911.933 ;
      RECT 331.049 0 335.959 911.933 ;
      RECT 322.409 0 327.319 911.933 ;
      RECT 304.697 0 318.679 911.933 ;
      RECT 296.057 0 300.967 911.933 ;
      RECT 287.417 0 292.327 911.933 ;
      RECT 278.777 0 283.687 911.933 ;
      RECT 270.137 0 275.047 911.933 ;
      RECT 261.497 0 266.407 911.933 ;
      RECT 252.857 0 257.767 911.933 ;
      RECT 244.217 0 249.127 911.933 ;
      RECT 235.577 0 240.487 911.933 ;
      RECT 226.937 0 231.847 911.933 ;
      RECT 218.297 0 223.207 911.933 ;
      RECT 209.657 0 214.567 911.933 ;
      RECT 201.017 0 205.927 911.933 ;
      RECT 192.377 0 197.287 911.933 ;
      RECT 183.737 0 188.647 911.933 ;
      RECT 175.097 0 180.007 911.933 ;
      RECT 166.457 0 171.367 911.933 ;
      RECT 148.745 0 162.727 911.933 ;
      RECT 140.105 0 145.015 911.933 ;
      RECT 131.465 0 136.375 911.933 ;
      RECT 122.825 0 127.735 911.933 ;
      RECT 114.185 0 119.095 911.933 ;
      RECT 105.545 0 110.455 911.933 ;
      RECT 96.905 0 101.815 911.933 ;
      RECT 88.265 0 93.175 911.933 ;
      RECT 79.625 0 84.535 911.933 ;
      RECT 70.985 0 75.895 911.933 ;
      RECT 62.345 0 67.255 911.933 ;
      RECT 53.705 0 58.615 911.933 ;
      RECT 45.065 0 49.975 911.933 ;
      RECT 36.425 0 41.335 911.933 ;
      RECT 27.785 0 32.695 911.933 ;
      RECT 19.145 0 24.055 911.933 ;
      RECT 10.505 0 15.415 911.933 ;
      RECT 0 0 6.775 911.933 ;
      RECT 0 0 623.808 782.8775 ;
    LAYER gmz SPACING 0.54 ;
      RECT 0 910.644 623.808 911.933 ;
      RECT 616.601 0 623.808 911.933 ;
      RECT 607.961 0 612.871 911.933 ;
      RECT 599.321 0 604.231 911.933 ;
      RECT 590.681 0 595.591 911.933 ;
      RECT 582.041 0 586.951 911.933 ;
      RECT 573.401 0 578.311 911.933 ;
      RECT 564.761 0 569.671 911.933 ;
      RECT 556.121 0 561.031 911.933 ;
      RECT 547.481 0 552.391 911.933 ;
      RECT 538.841 0 543.751 911.933 ;
      RECT 530.201 0 535.111 911.933 ;
      RECT 521.561 0 526.471 911.933 ;
      RECT 512.921 0 517.831 911.933 ;
      RECT 504.281 0 509.191 911.933 ;
      RECT 495.641 0 500.551 911.933 ;
      RECT 487.001 0 491.911 911.933 ;
      RECT 478.361 0 483.271 911.933 ;
      RECT 460.649 0 474.631 911.933 ;
      RECT 452.009 0 456.919 911.933 ;
      RECT 443.369 0 448.279 911.933 ;
      RECT 434.729 0 439.639 911.933 ;
      RECT 426.089 0 430.999 911.933 ;
      RECT 417.449 0 422.359 911.933 ;
      RECT 408.809 0 413.719 911.933 ;
      RECT 400.169 0 405.079 911.933 ;
      RECT 391.529 0 396.439 911.933 ;
      RECT 382.889 0 387.799 911.933 ;
      RECT 374.249 0 379.159 911.933 ;
      RECT 365.609 0 370.519 911.933 ;
      RECT 356.969 0 361.879 911.933 ;
      RECT 348.329 0 353.239 911.933 ;
      RECT 339.689 0 344.599 911.933 ;
      RECT 331.049 0 335.959 911.933 ;
      RECT 322.409 0 327.319 911.933 ;
      RECT 304.697 0 318.679 911.933 ;
      RECT 296.057 0 300.967 911.933 ;
      RECT 287.417 0 292.327 911.933 ;
      RECT 278.777 0 283.687 911.933 ;
      RECT 270.137 0 275.047 911.933 ;
      RECT 261.497 0 266.407 911.933 ;
      RECT 252.857 0 257.767 911.933 ;
      RECT 244.217 0 249.127 911.933 ;
      RECT 235.577 0 240.487 911.933 ;
      RECT 226.937 0 231.847 911.933 ;
      RECT 218.297 0 223.207 911.933 ;
      RECT 209.657 0 214.567 911.933 ;
      RECT 201.017 0 205.927 911.933 ;
      RECT 192.377 0 197.287 911.933 ;
      RECT 183.737 0 188.647 911.933 ;
      RECT 175.097 0 180.007 911.933 ;
      RECT 166.457 0 171.367 911.933 ;
      RECT 148.745 0 162.727 911.933 ;
      RECT 140.105 0 145.015 911.933 ;
      RECT 131.465 0 136.375 911.933 ;
      RECT 122.825 0 127.735 911.933 ;
      RECT 114.185 0 119.095 911.933 ;
      RECT 105.545 0 110.455 911.933 ;
      RECT 96.905 0 101.815 911.933 ;
      RECT 88.265 0 93.175 911.933 ;
      RECT 79.625 0 84.535 911.933 ;
      RECT 70.985 0 75.895 911.933 ;
      RECT 62.345 0 67.255 911.933 ;
      RECT 53.705 0 58.615 911.933 ;
      RECT 45.065 0 49.975 911.933 ;
      RECT 36.425 0 41.335 911.933 ;
      RECT 27.785 0 32.695 911.933 ;
      RECT 19.145 0 24.055 911.933 ;
      RECT 10.505 0 15.415 911.933 ;
      RECT 0 0 6.775 911.933 ;
      RECT 0 0 623.808 782.8775 ;
    LAYER gmb SPACING 1 ;
      RECT 0 0 623.808 911.933 ;
  END
END uni_2x2sub4x4_gpio_top_lef_LEFT_SIDE

END LIBRARY
