module mem_tlul (clk_i,
    rst_ni,
    en_ifetch_i,
    tl_i,
    tl_o);
 input clk_i;
 input rst_ni;
 input [3:0] en_ifetch_i;
 input [108:0] tl_i;
 output [65:0] tl_o;

 wire N1;
 wire n126;
 wire n131;
 wire n170;
 wire n175;
 wire n188;
 wire n189;
 wire n192;
 wire n197;
 wire n211;
 wire n322;
 wire n323;
 wire n324;
 wire n325;
 wire n326;
 wire n327;
 wire n328;
 wire n329;
 wire n330;
 wire n331;
 wire n332;
 wire n333;
 wire n334;
 wire n335;
 wire n336;
 wire n337;
 wire n338;
 wire n339;
 wire n340;
 wire n341;
 wire n342;
 wire n343;
 wire n344;
 wire n345;
 wire n346;
 wire n347;
 wire n348;
 wire n349;
 wire n350;
 wire n351;
 wire n352;
 wire n353;
 wire n354;
 wire n355;
 wire n356;
 wire n357;
 wire n358;
 wire n359;
 wire n360;
 wire n361;
 wire n362;
 wire n363;
 wire n364;
 wire n365;
 wire n366;
 wire n367;
 wire n368;
 wire n369;
 wire n370;
 wire n371;
 wire n372;
 wire n373;
 wire n374;
 wire n375;
 wire n376;
 wire n377;
 wire n378;
 wire n379;
 wire n380;
 wire n381;
 wire n382;
 wire n383;
 wire n384;
 wire n385;
 wire n386;
 wire n387;
 wire n388;
 wire n389;
 wire n390;
 wire n391;
 wire n392;
 wire n393;
 wire n394;
 wire n395;
 wire n396;
 wire n397;
 wire n401;
 wire n402;
 wire n403;
 wire n404;
 wire n405;
 wire n409;
 wire n410;
 wire n411;
 wire n412;
 wire n413;
 wire n414;
 wire n415;
 wire n416;
 wire n417;
 wire n418;
 wire n419;
 wire n420;
 wire n421;
 wire n424;
 wire n426;
 wire n427;
 wire n428;
 wire n429;
 wire n430;
 wire n431;
 wire n432;
 wire n433;
 wire n434;
 wire n438;
 wire n439;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire n_0_net_;
 wire clknet_0_clk_i;
 wire rvalid;
 wire u_tlul_adapter_sram_N210;
 wire u_tlul_adapter_sram_reqfifo_wdata_op__0_;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_rptr_1_;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_wptr_1_;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_rptr_value_0_;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N11;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N23;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N25;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst;
 wire u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_wptr_value_0_;
 wire u_tlul_adapter_sram_u_reqfifo_net644;
 wire u_tlul_adapter_sram_u_reqfifo_net650;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_rptr_1_;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_wptr_1_;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_rptr_value_0_;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N11;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N23;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N25;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst;
 wire u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_wptr_value_0_;
 wire u_tlul_adapter_sram_u_rspfifo_net616;
 wire u_tlul_adapter_sram_u_rspfifo_net622;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_rptr_1_;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_wptr_1_;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_rptr_value_0_;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N11;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N23;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N25;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst;
 wire u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_wptr_value_0_;
 wire wen;
 wire net285;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_1_1__leaf_clk_i;
 wire clknet_0_u_tlul_adapter_sram_u_rspfifo_net616;
 wire clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net616;
 wire clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net616;
 wire clknet_0_u_tlul_adapter_sram_u_rspfifo_net622;
 wire clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622;
 wire clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622;
 wire clknet_0_u_tlul_adapter_sram_u_reqfifo_net644;
 wire clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net644;
 wire clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net644;
 wire clknet_0_u_tlul_adapter_sram_u_reqfifo_net650;
 wire clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net650;
 wire clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net650;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire [10:0] addr;
 wire [31:0] rdata;
 wire [31:0] u_tlul_adapter_sram_rdata_tlword;
 wire [16:0] u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata;
 wire [39:0] u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata;
 wire [4:0] u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata;
 wire [31:0] wdata;

 b15inv000as1n80x5 U430 (.a(net12),
    .o1(n328));
 b15nonb02aq1n16x5 U431 (.a(net57),
    .b(net172),
    .out0(addr[2]));
 b15nonb02aq1n03x5 U432 (.a(net56),
    .b(net171),
    .out0(addr[1]));
 b15nonb02as1n16x5 U433 (.a(net55),
    .b(net171),
    .out0(addr[0]));
 b15nonb02an1n16x5 U434 (.a(net59),
    .b(net172),
    .out0(addr[4]));
 b15nonb02as1n16x5 U435 (.a(net174),
    .b(net172),
    .out0(addr[3]));
 b15nonb02as1n16x5 U436 (.a(net61),
    .b(net172),
    .out0(addr[6]));
 b15nonb02ah1n16x5 U437 (.a(net63),
    .b(net172),
    .out0(addr[8]));
 b15nonb02ah1n16x5 U438 (.a(net60),
    .b(net172),
    .out0(addr[5]));
 b15nonb02aq1n16x5 U439 (.a(net65),
    .b(net172),
    .out0(addr[10]));
 b15nonb02as1n16x5 U440 (.a(net64),
    .b(net172),
    .out0(addr[9]));
 b15nonb02ah1n16x5 U441 (.a(net62),
    .b(net172),
    .out0(addr[7]));
 b15norp03as1n24x5 U442 (.a(net11),
    .b(net10),
    .c(n328),
    .o1(wen));
 b15nandp2an1n24x5 U443 (.a(net177),
    .b(net157),
    .o1(n322));
 b15nonb02ar1n12x5 U444 (.a(net21),
    .b(n322),
    .out0(wdata[4]));
 b15nonb02an1n08x5 U445 (.a(net20),
    .b(n322),
    .out0(wdata[3]));
 b15nonb02ah1n06x5 U446 (.a(net19),
    .b(n322),
    .out0(wdata[2]));
 b15nonb02al1n08x5 U447 (.a(net18),
    .b(n322),
    .out0(wdata[1]));
 b15nonb02al1n12x5 U448 (.a(net23),
    .b(n322),
    .out0(wdata[6]));
 b15nonb02ar1n12x5 U449 (.a(net22),
    .b(n322),
    .out0(wdata[5]));
 b15nonb02aq1n06x5 U450 (.a(net17),
    .b(n322),
    .out0(wdata[0]));
 b15nand02ah1n48x5 U451 (.a(net175),
    .b(net157),
    .o1(n323));
 b15nonb02an1n12x5 U452 (.a(net25),
    .b(n323),
    .out0(wdata[8]));
 b15nonb02ah1n08x5 U453 (.a(net24),
    .b(n322),
    .out0(wdata[7]));
 b15nonb02aq1n12x5 U454 (.a(net26),
    .b(n323),
    .out0(wdata[9]));
 b15nonb02al1n16x5 U455 (.a(net27),
    .b(n323),
    .out0(wdata[10]));
 b15nonb02as1n12x5 U456 (.a(net28),
    .b(n323),
    .out0(wdata[11]));
 b15nonb02aq1n16x5 U457 (.a(net29),
    .b(n323),
    .out0(wdata[12]));
 b15nonb02aq1n16x5 U458 (.a(net30),
    .b(n323),
    .out0(wdata[13]));
 b15nonb02aq1n16x5 U459 (.a(net31),
    .b(n323),
    .out0(wdata[14]));
 b15nonb02ah1n16x5 U460 (.a(net32),
    .b(n323),
    .out0(wdata[15]));
 b15inv040as1n12x5 U461 (.a(net157),
    .o1(n_0_net_));
 b15inv040ah1n12x5 U462 (.a(net52),
    .o1(n347));
 b15norp02an1n48x5 U463 (.a(n347),
    .b(net144),
    .o1(n324));
 b15and002an1n08x5 U464 (.a(n324),
    .b(net48),
    .o(wdata[31]));
 b15and002an1n08x5 U465 (.a(n324),
    .b(net47),
    .o(wdata[30]));
 b15and002an1n08x5 U466 (.a(n324),
    .b(net46),
    .o(wdata[29]));
 b15and002an1n08x5 U467 (.a(n324),
    .b(net45),
    .o(wdata[28]));
 b15and002an1n08x5 U468 (.a(n324),
    .b(net44),
    .o(wdata[27]));
 b15and002ar1n12x5 U469 (.a(n324),
    .b(net43),
    .o(wdata[26]));
 b15and002al1n08x5 U470 (.a(n324),
    .b(net42),
    .o(wdata[25]));
 b15and002ah1n08x5 U471 (.a(n324),
    .b(net41),
    .o(wdata[24]));
 b15inv000ah1n12x5 U472 (.a(net51),
    .o1(n345));
 b15norp02aq1n48x5 U473 (.a(n345),
    .b(net144),
    .o1(n325));
 b15and002aq1n12x5 U474 (.a(n325),
    .b(net40),
    .o(wdata[23]));
 b15and002al1n16x5 U475 (.a(n325),
    .b(net39),
    .o(wdata[22]));
 b15and002aq1n12x5 U476 (.a(n325),
    .b(net38),
    .o(wdata[21]));
 b15and002aq1n12x5 U477 (.a(n325),
    .b(net37),
    .o(wdata[20]));
 b15and002an1n12x5 U478 (.a(n325),
    .b(net36),
    .o(wdata[19]));
 b15and002ar1n16x5 U479 (.a(n325),
    .b(net35),
    .o(wdata[18]));
 b15and002aq1n12x5 U480 (.a(n325),
    .b(net34),
    .o(wdata[17]));
 b15and002al1n16x5 U481 (.a(n325),
    .b(net33),
    .o(wdata[16]));
 b15xor002an1n16x5 U482 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_wptr_1_),
    .b(net161),
    .out0(n360));
 b15inv040as1n12x5 U483 (.a(net164),
    .o1(n327));
 b15inv000ar1n20x5 U484 (.a(net163),
    .o1(n365));
 b15aoi022as1n48x5 U485 (.a(net162),
    .b(n327),
    .c(net164),
    .d(n365),
    .o1(n359));
 b15nanb02as1n24x5 U486 (.a(n360),
    .b(n359),
    .out0(n418));
 b15inv040aq1n05x5 U487 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst),
    .o1(n356));
 b15xor002as1n08x5 U488 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_rptr_value_0_),
    .b(net349),
    .out0(n358));
 b15inv000an1n03x5 U489 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_rptr_1_),
    .o1(n326));
 b15aboi22as1n12x5 U490 (.a(net369),
    .b(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_rptr_1_),
    .c(net369),
    .d(n326),
    .out0(n357));
 b15nanb02an1n16x5 U491 (.a(net350),
    .b(net370),
    .out0(n384));
 b15nandp2ah1n12x5 U492 (.a(n356),
    .b(net371),
    .o1(n374));
 b15inv040as1n05x5 U493 (.a(net372),
    .o1(n373));
 b15nand02ah1n12x5 U494 (.a(n373),
    .b(net363),
    .o1(n369));
 b15nonb03as1n12x5 U495 (.a(n418),
    .b(net159),
    .c(n369),
    .out0(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N23));
 b15nor002an1n16x5 U496 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .b(n327),
    .o1(n175));
 b15aoi112ar1n08x5 U497 (.a(net10),
    .b(n328),
    .c(net13),
    .d(net178),
    .o1(n355));
 b15norp02an1n02x5 U498 (.a(net52),
    .b(net50),
    .o1(n330));
 b15norp02ar1n02x5 U499 (.a(net51),
    .b(net49),
    .o1(n329));
 b15inv000as1n03x5 U500 (.a(net53),
    .o1(n343));
 b15aoi022an1n04x5 U501 (.a(net53),
    .b(n330),
    .c(n329),
    .d(n343),
    .o1(n331));
 b15aboi22aq1n02x5 U502 (.a(net173),
    .b(n331),
    .c(net49),
    .d(net50),
    .out0(n334));
 b15inv000al1n02x5 U503 (.a(net8),
    .o1(n332));
 b15aoai13al1n03x5 U504 (.a(net51),
    .b(n332),
    .c(net49),
    .d(net50),
    .o1(n333));
 b15oai022an1n08x5 U505 (.a(net8),
    .b(n334),
    .c(n333),
    .d(n347),
    .o1(n340));
 b15inv000an1n08x5 U506 (.a(net11),
    .o1(n439));
 b15inv020ah1n06x5 U507 (.a(net14),
    .o1(n336));
 b15nor004ah1n06x5 U508 (.a(net4),
    .b(net1),
    .c(n439),
    .d(n336),
    .o1(n335));
 b15aoi013al1n08x5 U509 (.a(net16),
    .b(net2),
    .c(net3),
    .d(n335),
    .o1(n338));
 b15obai22ar1n16x5 U510 (.a(net16),
    .b(net13),
    .c(net178),
    .d(n336),
    .out0(n337));
 b15aoi112aq1n02x5 U511 (.a(n338),
    .b(n337),
    .c(net173),
    .d(net53),
    .o1(n339));
 b15oai013as1n03x5 U512 (.a(n339),
    .b(n340),
    .c(net9),
    .d(net11),
    .o1(n341));
 b15aoi012al1n06x5 U513 (.a(n341),
    .b(net9),
    .c(net11),
    .o1(n354));
 b15aoi022an1n04x5 U514 (.a(net53),
    .b(net49),
    .c(net50),
    .d(n343),
    .o1(n344));
 b15nor002an1n06x5 U515 (.a(net54),
    .b(net51),
    .o1(n348));
 b15inv000ah1n04x5 U516 (.a(net54),
    .o1(n342));
 b15norp03ah1n12x5 U517 (.a(net49),
    .b(net50),
    .c(n342),
    .o1(n346));
 b15aoi022as1n06x5 U518 (.a(n344),
    .b(n348),
    .c(n346),
    .d(n343),
    .o1(n351));
 b15aoi013al1n06x5 U519 (.a(net8),
    .b(net53),
    .c(n346),
    .d(n345),
    .o1(n350));
 b15aoai13an1n06x5 U520 (.a(net173),
    .b(n346),
    .c(n348),
    .d(n347),
    .o1(n349));
 b15oai112as1n16x5 U521 (.a(n350),
    .b(n349),
    .c(net52),
    .d(n351),
    .o1(n353));
 b15oai013an1n08x5 U522 (.a(net8),
    .b(net54),
    .c(net53),
    .d(net173),
    .o1(n352));
 b15nand04as1n16x5 U523 (.a(n355),
    .b(n354),
    .c(n353),
    .d(n352),
    .o1(u_tlul_adapter_sram_N210));
 b15oai012aq1n16x5 U524 (.a(n356),
    .b(net350),
    .c(n357),
    .o1(n361));
 b15norp03as1n24x5 U525 (.a(wen),
    .b(n361),
    .c(u_tlul_adapter_sram_N210),
    .o1(N1));
 b15aoi012ar1n16x5 U526 (.a(net159),
    .b(n360),
    .c(n359),
    .o1(n362));
 b15nand02ar1n24x5 U527 (.a(n362),
    .b(N1),
    .o1(n364));
 b15norp02ar1n08x5 U528 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_wptr_1_),
    .b(n364),
    .o1(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N11));
 b15nonb02ah1n06x5 U529 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .b(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_rptr_1_),
    .out0(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N25));
 b15nonb02ah1n12x5 U530 (.a(net552),
    .b(net351),
    .out0(net74));
 b15nandp2al1n16x5 U531 (.a(net12),
    .b(net74),
    .o1(n363));
 b15qgbno2an1n10x5 U532 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_wptr_1_),
    .b(n363),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N11));
 b15inv020ar1n40x5 U533 (.a(n363),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9));
 b15nonb02as1n12x5 U534 (.a(net169),
    .b(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .out0(n170));
 b15inv000aq1n40x5 U535 (.a(n364),
    .o1(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9));
 b15norp02an1n16x5 U536 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .b(n365),
    .o1(n192));
 b15nonb02aq1n16x5 U537 (.a(n188),
    .b(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .out0(n189));
 b15inv000an1n08x5 U538 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_rptr_1_),
    .o1(n372));
 b15obai22aq1n24x5 U539 (.a(net384),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_rptr_1_),
    .c(n372),
    .d(net384),
    .out0(n367));
 b15inv000ar1n16x5 U540 (.a(net355),
    .o1(n366));
 b15inv000al1n10x5 U541 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_rptr_value_0_),
    .o1(n370));
 b15aoi022aq1n32x5 U542 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_rptr_value_0_),
    .b(n366),
    .c(net355),
    .d(n370),
    .o1(n368));
 b15aoi112as1n08x5 U543 (.a(net165),
    .b(n369),
    .c(n367),
    .d(n368),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9));
 b15qgbno2an1n10x5 U544 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .b(n366),
    .o1(n126));
 b15nonb02as1n16x5 U545 (.a(net356),
    .b(net385),
    .out0(n380));
 b15inv040ah1n16x5 U546 (.a(net357),
    .o1(n386));
 b15ao0012aq1n08x5 U547 (.a(net165),
    .b(net364),
    .c(net357),
    .o(n375));
 b15nanb02as1n24x5 U548 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[16]),
    .b(net379),
    .out0(n379));
 b15nor004as1n12x5 U549 (.a(net365),
    .b(n379),
    .c(n374),
    .d(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[14]),
    .o1(n385));
 b15aob012as1n24x5 U550 (.a(net374),
    .b(net377),
    .c(net358),
    .out0(net125));
 b15aob012as1n24x5 U551 (.a(net366),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[2]),
    .c(net358),
    .out0(net101));
 b15aob012as1n24x5 U552 (.a(net374),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[4]),
    .c(net358),
    .out0(net121));
 b15nonb02aq1n08x5 U553 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .b(net167),
    .out0(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N11));
 b15inv000al1n24x5 U554 (.a(net366),
    .o1(n382));
 b15nonb02as1n16x5 U555 (.a(net6),
    .b(n382),
    .out0(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N23));
 b15nor002an1n12x5 U556 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .b(n370),
    .o1(n131));
 b15norp02an1n16x5 U557 (.a(net357),
    .b(n382),
    .o1(n371));
 b15and002aq1n16x5 U558 (.a(n371),
    .b(net391),
    .o(net111));
 b15and002ar1n24x5 U559 (.a(n371),
    .b(net403),
    .o(net90));
 b15and002aq1n16x5 U560 (.a(n371),
    .b(net389),
    .o(net126));
 b15and002aq1n16x5 U561 (.a(n371),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[5]),
    .o(net124));
 b15and002al1n08x5 U562 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .b(n372),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N25));
 b15nand02ah1n16x5 U563 (.a(n373),
    .b(net380),
    .o1(net122));
 b15inv020aq1n05x5 U564 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[14]),
    .o1(n377));
 b15aoai13as1n08x5 U565 (.a(net381),
    .b(net372),
    .c(n377),
    .d(net365),
    .o1(net123));
 b15inv040as1n36x5 U566 (.a(net395),
    .o1(n376));
 b15nonb02al1n12x5 U567 (.a(net500),
    .b(n376),
    .out0(net119));
 b15nonb02al1n08x5 U568 (.a(net486),
    .b(n376),
    .out0(net113));
 b15nonb02ah1n08x5 U569 (.a(net523),
    .b(n376),
    .out0(net118));
 b15nonb02al1n08x5 U570 (.a(net483),
    .b(n376),
    .out0(net117));
 b15nonb02ah1n08x5 U571 (.a(net397),
    .b(n376),
    .out0(net115));
 b15nonb02ah1n08x5 U572 (.a(net405),
    .b(n376),
    .out0(net116));
 b15nonb02ah1n08x5 U573 (.a(net400),
    .b(n376),
    .out0(net110));
 b15nonb02ah1n08x5 U574 (.a(net520),
    .b(n376),
    .out0(net114));
 b15nonb02ah1n08x5 U575 (.a(net529),
    .b(n376),
    .out0(net120));
 b15nonb02ah1n08x5 U576 (.a(net408),
    .b(n376),
    .out0(net112));
 b15nonb02as1n16x5 U577 (.a(net6),
    .b(n376),
    .out0(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N23));
 b15nonb02ah1n12x5 U578 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_rptr_value_0_),
    .b(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .out0(n197));
 b15nonb02aq1n08x5 U579 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .b(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_rptr_1_),
    .out0(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N25));
 b15nand02aq1n16x5 U580 (.a(net155),
    .b(net358),
    .o1(n378));
 b15oaoi13as1n08x5 U581 (.a(n376),
    .b(n377),
    .c(net380),
    .d(net359),
    .o1(net79));
 b15nand02ar1n16x5 U582 (.a(net532),
    .b(n418),
    .o1(n397));
 b15nonb02al1n12x5 U583 (.a(rdata[26]),
    .b(net143),
    .out0(u_tlul_adapter_sram_rdata_tlword[26]));
 b15norp03as1n24x5 U584 (.a(net357),
    .b(net155),
    .c(n382),
    .o1(n381));
 b15inv000ar1n03x5 U585 (.a(net285),
    .o1(tl_o[9]));
 b15nor002an1n32x5 U587 (.a(net358),
    .b(n382),
    .o1(n383));
 b15inv000ar1n03x5 U588 (.a(net286),
    .o1(tl_o[10]));
 b15aoi022ah1n12x5 U590 (.a(net133),
    .b(net417),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[26]),
    .o1(n390));
 b15nandp3aq1n24x5 U591 (.a(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[12]),
    .b(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[11]),
    .c(net371),
    .o1(n388));
 b15aob012aq1n06x5 U592 (.a(net366),
    .b(net155),
    .c(net358),
    .out0(n387));
 b15oai013as1n12x5 U593 (.a(n387),
    .b(net429),
    .c(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[10]),
    .d(n388),
    .o1(n389));
 b15inv000ar1n03x5 U594 (.a(net287),
    .o1(tl_o[11]));
 b15nandp2ah1n04x5 U596 (.a(net418),
    .b(net127),
    .o1(net104));
 b15nonb02as1n16x5 U597 (.a(rdata[27]),
    .b(net534),
    .out0(u_tlul_adapter_sram_rdata_tlword[27]));
 b15aoi022al1n08x5 U598 (.a(net135),
    .b(net546),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[27]),
    .o1(n391));
 b15nandp2ar1n12x5 U599 (.a(net547),
    .b(net127),
    .o1(net105));
 b15nonb02aq1n12x5 U600 (.a(rdata[24]),
    .b(net534),
    .out0(u_tlul_adapter_sram_rdata_tlword[24]));
 b15aoi022aq1n12x5 U601 (.a(net133),
    .b(net537),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[24]),
    .o1(n392));
 b15inv000ar1n03x5 U602 (.a(net288),
    .o1(tl_o[12]));
 b15nand02as1n04x5 U603 (.a(net538),
    .b(net127),
    .o1(net102));
 b15nonb02aq1n12x5 U604 (.a(rdata[25]),
    .b(net143),
    .out0(u_tlul_adapter_sram_rdata_tlword[25]));
 b15aoi022aq1n12x5 U605 (.a(net133),
    .b(net526),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[25]),
    .o1(n393));
 b15qgbna2an1n05x5 U606 (.o1(net103),
    .a(net527),
    .b(net127));
 b15nonb02aq1n16x5 U607 (.a(rdata[30]),
    .b(net143),
    .out0(u_tlul_adapter_sram_rdata_tlword[30]));
 b15aoi022ar1n24x5 U608 (.a(net133),
    .b(net543),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[30]),
    .o1(n394));
 b15nand02an1n16x5 U609 (.a(net544),
    .b(net127),
    .o1(net108));
 b15nonb02aq1n16x5 U610 (.a(rdata[31]),
    .b(net143),
    .out0(u_tlul_adapter_sram_rdata_tlword[31]));
 b15aoi022an1n12x5 U611 (.a(net133),
    .b(net489),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[31]),
    .o1(n395));
 b15nand02ah1n04x5 U612 (.a(net490),
    .b(net127),
    .o1(net109));
 b15nonb02ah1n16x5 U613 (.a(rdata[28]),
    .b(net534),
    .out0(u_tlul_adapter_sram_rdata_tlword[28]));
 b15aoi022aq1n08x5 U614 (.a(net133),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[36]),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[28]),
    .o1(n396));
 b15nand02al1n06x5 U615 (.a(net535),
    .b(net129),
    .o1(net106));
 b15nonb02al1n16x5 U616 (.a(rdata[29]),
    .b(net143),
    .out0(u_tlul_adapter_sram_rdata_tlword[29]));
 b15aoi022al1n16x5 U617 (.a(net133),
    .b(net503),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[29]),
    .o1(n401));
 b15nand02aq1n12x5 U618 (.a(net504),
    .b(net127),
    .o1(net107));
 b15nand02aq1n08x5 U619 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[3]),
    .b(n418),
    .o1(n434));
 b15nonb02as1n12x5 U620 (.a(rdata[20]),
    .b(net142),
    .out0(u_tlul_adapter_sram_rdata_tlword[20]));
 b15inv000ar1n03x5 U622 (.a(net289),
    .o1(tl_o[13]));
 b15aoi022al1n12x5 U623 (.a(net135),
    .b(net496),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[20]),
    .o1(n402));
 b15nand02al1n08x5 U624 (.a(net497),
    .b(net129),
    .o1(net97));
 b15nonb02ah1n12x5 U625 (.a(rdata[21]),
    .b(net142),
    .out0(u_tlul_adapter_sram_rdata_tlword[21]));
 b15aoi022an1n16x5 U626 (.a(net133),
    .b(net450),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[21]),
    .o1(n403));
 b15nandp2an1n05x5 U627 (.a(net451),
    .b(net127),
    .o1(net98));
 b15nonb02aq1n16x5 U628 (.a(rdata[22]),
    .b(net142),
    .out0(u_tlul_adapter_sram_rdata_tlword[22]));
 b15aoi022an1n16x5 U629 (.a(net133),
    .b(net513),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[22]),
    .o1(n404));
 b15nandp2ah1n08x5 U630 (.a(net514),
    .b(net127),
    .o1(net99));
 b15nonb02ah1n16x5 U631 (.a(rdata[23]),
    .b(net142),
    .out0(u_tlul_adapter_sram_rdata_tlword[23]));
 b15aoi022aq1n12x5 U632 (.a(net133),
    .b(net421),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[23]),
    .o1(n405));
 b15nandp2ah1n05x5 U633 (.a(net422),
    .b(net127),
    .o1(net100));
 b15nandp2an1n48x5 U634 (.a(net411),
    .b(n418),
    .o1(n416));
 b15nonb02an1n04x5 U635 (.a(rdata[0]),
    .b(net412),
    .out0(u_tlul_adapter_sram_rdata_tlword[0]));
 b15inv000ar1n03x5 U637 (.a(net290),
    .o1(tl_o[14]));
 b15aoi022ah1n48x5 U638 (.a(net134),
    .b(net493),
    .c(net132),
    .d(net141),
    .o1(n409));
 b15nand02al1n06x5 U640 (.a(net494),
    .b(net431),
    .o1(net75));
 b15nonb02as1n16x5 U641 (.a(rdata[1]),
    .b(net412),
    .out0(u_tlul_adapter_sram_rdata_tlword[1]));
 b15aoi022aq1n48x5 U642 (.a(net134),
    .b(net443),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[1]),
    .o1(n410));
 b15nand02ah1n04x5 U643 (.a(net444),
    .b(net431),
    .o1(net76));
 b15nonb02an1n04x5 U644 (.a(rdata[2]),
    .b(net412),
    .out0(u_tlul_adapter_sram_rdata_tlword[2]));
 b15aoi022ah1n48x5 U645 (.a(net134),
    .b(net517),
    .c(net132),
    .d(net140),
    .o1(n411));
 b15nandp2ar1n05x5 U646 (.a(net518),
    .b(net431),
    .o1(net77));
 b15nonb02as1n16x5 U647 (.a(rdata[3]),
    .b(net412),
    .out0(u_tlul_adapter_sram_rdata_tlword[3]));
 b15aoi022aq1n48x5 U648 (.a(net134),
    .b(net458),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[3]),
    .o1(n412));
 b15nand02al1n06x5 U649 (.a(net459),
    .b(net431),
    .o1(net78));
 b15nonb02aq1n03x5 U650 (.a(rdata[4]),
    .b(net412),
    .out0(u_tlul_adapter_sram_rdata_tlword[4]));
 b15aoi022ah1n12x5 U651 (.a(net134),
    .b(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[12]),
    .c(net132),
    .d(net139),
    .o1(n413));
 b15nandp2ah1n16x5 U652 (.a(n413),
    .b(net128),
    .o1(net80));
 b15nonb02as1n16x5 U653 (.a(rdata[5]),
    .b(net412),
    .out0(u_tlul_adapter_sram_rdata_tlword[5]));
 b15aoi022as1n16x5 U654 (.a(net134),
    .b(net477),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[5]),
    .o1(n414));
 b15nand02ar1n32x5 U655 (.a(net478),
    .b(net128),
    .o1(net81));
 b15nonb02as1n16x5 U656 (.a(rdata[6]),
    .b(net412),
    .out0(u_tlul_adapter_sram_rdata_tlword[6]));
 b15aoi022an1n48x5 U657 (.a(net134),
    .b(net462),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[6]),
    .o1(n415));
 b15nandp2aq1n04x5 U658 (.a(net463),
    .b(net431),
    .o1(net82));
 b15nonb02as1n16x5 U659 (.a(rdata[7]),
    .b(net412),
    .out0(u_tlul_adapter_sram_rdata_tlword[7]));
 b15aoi022aq1n48x5 U660 (.a(net134),
    .b(net151),
    .c(net132),
    .d(net413),
    .o1(n417));
 b15nand02ah1n04x5 U661 (.a(net414),
    .b(net130),
    .o1(net83));
 b15nandp2ah1n48x5 U662 (.a(net437),
    .b(n418),
    .o1(n429));
 b15nonb02as1n16x5 U663 (.a(rdata[8]),
    .b(net438),
    .out0(u_tlul_adapter_sram_rdata_tlword[8]));
 b15aoi022as1n48x5 U664 (.a(net134),
    .b(net447),
    .c(n383),
    .d(u_tlul_adapter_sram_rdata_tlword[8]),
    .o1(n419));
 b15nand02aq1n12x5 U665 (.a(net448),
    .b(net431),
    .o1(net84));
 b15nonb02as1n16x5 U666 (.a(rdata[9]),
    .b(net438),
    .out0(u_tlul_adapter_sram_rdata_tlword[9]));
 b15aoi022aq1n48x5 U667 (.a(net134),
    .b(net474),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[9]),
    .o1(n420));
 b15nand02aq1n12x5 U668 (.a(net475),
    .b(net431),
    .o1(net85));
 b15nonb02aq1n03x5 U669 (.a(rdata[10]),
    .b(net438),
    .out0(u_tlul_adapter_sram_rdata_tlword[10]));
 b15aoi022as1n08x5 U670 (.a(net135),
    .b(net540),
    .c(net132),
    .d(net138),
    .o1(n421));
 b15nandp2ar1n08x5 U671 (.a(net541),
    .b(net129),
    .o1(net86));
 b15nonb02as1n16x5 U672 (.a(rdata[11]),
    .b(net438),
    .out0(u_tlul_adapter_sram_rdata_tlword[11]));
 b15aoi022aq1n48x5 U673 (.a(n381),
    .b(net148),
    .c(net132),
    .d(net439),
    .o1(n424));
 b15nand02ar1n16x5 U674 (.a(net440),
    .b(net431),
    .o1(net87));
 b15nonb02aq1n03x5 U675 (.a(rdata[12]),
    .b(n429),
    .out0(u_tlul_adapter_sram_rdata_tlword[12]));
 b15aoi022aq1n08x5 U676 (.a(net135),
    .b(net434),
    .c(net132),
    .d(net137),
    .o1(n426));
 b15nandp2ah1n05x5 U677 (.a(net435),
    .b(net127),
    .o1(net88));
 b15nonb02as1n16x5 U678 (.a(rdata[13]),
    .b(n429),
    .out0(u_tlul_adapter_sram_rdata_tlword[13]));
 b15aoi022aq1n12x5 U679 (.a(net133),
    .b(net425),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[13]),
    .o1(n427));
 b15nand02ah1n06x5 U680 (.a(net426),
    .b(net127),
    .o1(net89));
 b15nonb02as1n16x5 U681 (.a(rdata[14]),
    .b(net438),
    .out0(u_tlul_adapter_sram_rdata_tlword[14]));
 b15aoi022aq1n08x5 U682 (.a(net135),
    .b(net454),
    .c(net132),
    .d(u_tlul_adapter_sram_rdata_tlword[14]),
    .o1(n428));
 b15nand02an1n08x5 U683 (.a(net455),
    .b(net127),
    .o1(net91));
 b15nonb02as1n16x5 U684 (.a(net179),
    .b(net438),
    .out0(u_tlul_adapter_sram_rdata_tlword[15]));
 b15aoi022an1n08x5 U685 (.a(net133),
    .b(net480),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[15]),
    .o1(n430));
 b15nandp2al1n08x5 U686 (.a(net481),
    .b(net127),
    .o1(net92));
 b15nonb02as1n08x5 U687 (.a(rdata[16]),
    .b(net142),
    .out0(u_tlul_adapter_sram_rdata_tlword[16]));
 b15aoi022as1n12x5 U688 (.a(net133),
    .b(net469),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[16]),
    .o1(n431));
 b15nand02al1n12x5 U689 (.a(net470),
    .b(net127),
    .o1(net93));
 b15nonb02al1n12x5 U690 (.a(rdata[17]),
    .b(net142),
    .out0(u_tlul_adapter_sram_rdata_tlword[17]));
 b15aoi022an1n06x5 U691 (.a(net133),
    .b(net506),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[17]),
    .o1(n432));
 b15nandp2ar1n08x5 U692 (.a(net507),
    .b(net129),
    .o1(net94));
 b15nonb02ah1n16x5 U693 (.a(rdata[18]),
    .b(net142),
    .out0(u_tlul_adapter_sram_rdata_tlword[18]));
 b15aoi022al1n16x5 U694 (.a(net133),
    .b(net509),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[18]),
    .o1(n433));
 b15nandp2as1n03x5 U695 (.a(net510),
    .b(net127),
    .o1(net95));
 b15nonb02aq1n12x5 U696 (.a(rdata[19]),
    .b(net142),
    .out0(u_tlul_adapter_sram_rdata_tlword[19]));
 b15aoi022aq1n08x5 U697 (.a(net133),
    .b(net465),
    .c(net131),
    .d(u_tlul_adapter_sram_rdata_tlword[19]),
    .o1(n438));
 b15nandp2ah1n04x5 U698 (.a(net466),
    .b(net129),
    .o1(net96));
 b15norp03as1n24x5 U700 (.a(net9),
    .b(net10),
    .c(n439),
    .o1(u_tlul_adapter_sram_reqfifo_wdata_op__0_));
 b15inv000ar1n03x5 U702 (.a(net291),
    .o1(tl_o[15]));
 b15inv000ar1n03x5 U704 (.a(net292),
    .o1(tl_o[48]));
 b15inv000ar1n03x5 U706 (.a(net293),
    .o1(tl_o[59]));
 b15inv000ar1n03x5 U708 (.a(net294),
    .o1(tl_o[60]));
 b15inv000ar1n03x5 U710 (.a(net295),
    .o1(tl_o[61]));
 b15inv000ar1n03x5 U712 (.a(net296),
    .o1(tl_o[63]));
 b15inv000ar1n03x5 U714 (.a(net297),
    .o1(tl_o[64]));
 b15ztpn00an1n08x5 PHY_5 ();
 b15ztpn00an1n08x5 PHY_4 ();
 b15ztpn00an1n08x5 PHY_3 ();
 b15ztpn00an1n08x5 PHY_2 ();
 b15ztpn00an1n08x5 PHY_1 ();
 b15ztpn00an1n08x5 PHY_0 ();
 b15fqy203ar1n02x5 rvalid_reg_u_tlul_adapter_sram_intg_error_q_reg (.rb(net176),
    .clk(clknet_1_1__leaf_clk_i),
    .d1(N1),
    .d2(net549),
    .o1(rvalid),
    .o2(n211),
    .si1(net180),
    .si2(net181),
    .ssb(net298));
 ip224uhdlp1p11rf_2048x32m8b2c1s0_t0r0p0d0a1m1h u_sram (.clkbyp(net182),
    .fwen(net183),
    .mcen(net187),
    .ren(net145),
    .wen(net158),
    .wpulseen(net299),
    .clk(clknet_1_1__leaf_clk_i),
    .adr({addr[10],
    addr[9],
    addr[8],
    addr[7],
    addr[6],
    addr[5],
    addr[4],
    addr[3],
    addr[2],
    addr[1],
    addr[0]}),
    .din({wdata[31],
    wdata[30],
    wdata[29],
    wdata[28],
    wdata[27],
    wdata[26],
    wdata[25],
    wdata[24],
    wdata[23],
    wdata[22],
    wdata[21],
    wdata[20],
    wdata[19],
    wdata[18],
    wdata[17],
    wdata[16],
    wdata[15],
    wdata[14],
    wdata[13],
    wdata[12],
    wdata[11],
    wdata[10],
    wdata[9],
    wdata[8],
    wdata[7],
    wdata[6],
    wdata[5],
    wdata[4],
    wdata[3],
    wdata[2],
    wdata[1],
    wdata[0]}),
    .mc({net186,
    net185,
    net184}),
    .q({rdata[31],
    rdata[30],
    rdata[29],
    rdata[28],
    rdata[27],
    rdata[26],
    rdata[25],
    rdata[24],
    rdata[23],
    rdata[22],
    rdata[21],
    rdata[20],
    rdata[19],
    rdata[18],
    rdata[17],
    rdata[16],
    rdata[15],
    rdata[14],
    rdata[13],
    rdata[12],
    rdata[11],
    rdata[10],
    rdata[9],
    rdata[8],
    rdata[7],
    rdata[6],
    rdata[5],
    rdata[4],
    rdata[3],
    rdata[2],
    rdata[1],
    rdata[0]}),
    .wa({net189,
    net188}),
    .wpulse({net191,
    net190}));
 b15cilb05ah1n02x3 u_tlul_adapter_sram_u_reqfifo_clk_gate_gen_normal_fifo_storage_reg_0__0_latch (.clk(clknet_1_0__leaf_clk_i),
    .clkout(u_tlul_adapter_sram_u_reqfifo_net650),
    .en(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .te(net192));
 b15cilb05ah1n02x3 u_tlul_adapter_sram_u_reqfifo_clk_gate_gen_normal_fifo_storage_reg_0__latch (.clk(clknet_1_0__leaf_clk_i),
    .clkout(u_tlul_adapter_sram_u_reqfifo_net644),
    .en(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .te(net193));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__1_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net644),
    .d1(net66),
    .d2(net67),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[0]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[1]),
    .si1(net194),
    .si2(net195),
    .ssb(net300));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__11__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__12_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net650),
    .d1(net14),
    .d2(net178),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[11]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[12]),
    .si1(net196),
    .si2(net197),
    .ssb(net301));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__13__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__14_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net650),
    .d1(net16),
    .d2(u_tlul_adapter_sram_N210),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[13]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[14]),
    .si1(net198),
    .si2(net199),
    .ssb(net302));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__15__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__16_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net650),
    .d1(u_tlul_adapter_sram_reqfifo_wdata_op__0_),
    .d2(net200),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[15]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[16]),
    .si1(net201),
    .si2(net202),
    .ssb(net303));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__3_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net644),
    .d1(net68),
    .d2(net69),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[2]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[3]),
    .si1(net203),
    .si2(net204),
    .ssb(net304));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__5_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net644),
    .d1(net70),
    .d2(net71),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[4]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[5]),
    .si1(net205),
    .si2(net206),
    .ssb(net305));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__7_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net644),
    .d1(net72),
    .d2(net73),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[6]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[7]),
    .si1(net207),
    .si2(net208),
    .ssb(net306));
 b15fpy000ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__8_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net644),
    .d(net173),
    .o(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[8]),
    .si(net209),
    .ssb(net307));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__9__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__10_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net650),
    .d1(net8),
    .d2(net13),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[9]),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[10]),
    .si1(net210),
    .si2(net211),
    .ssb(net308));
 b15fqy203ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0_ (.rb(net176),
    .clk(clknet_1_0__leaf_clk_i),
    .d1(n197),
    .d2(n170),
    .o1(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_rptr_value_0_),
    .o2(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_wptr_value_0_),
    .si1(net212),
    .si2(net213),
    .ssb(net309));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N25),
    .den(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .o(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_rptr_1_),
    .rb(net5),
    .si(net214),
    .ssb(net310));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N11),
    .den(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .o(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_wptr_1_),
    .rb(net5),
    .si(net215),
    .ssb(net311));
 b15fqy00car1n02x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst_reg (.clk(clknet_1_1__leaf_clk_i),
    .d(net216),
    .o(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst),
    .psb(net176),
    .si(net217),
    .ssb(net312));
 b15cilb05ah1n02x3 u_tlul_adapter_sram_u_rspfifo_clk_gate_gen_normal_fifo_storage_reg_0__0_latch (.clk(clknet_1_0__leaf_clk_i),
    .clkout(u_tlul_adapter_sram_u_rspfifo_net622),
    .en(net136),
    .te(net218));
 b15cilb05ah1n02x3 u_tlul_adapter_sram_u_rspfifo_clk_gate_gen_normal_fifo_storage_reg_0__latch (.clk(clknet_1_0__leaf_clk_i),
    .clkout(u_tlul_adapter_sram_u_rspfifo_net616),
    .en(net136),
    .te(net219));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(net220),
    .d2(net221),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[0]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[1]),
    .si1(net222),
    .si2(net223),
    .ssb(net313));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__10__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__11_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(net140),
    .d2(u_tlul_adapter_sram_rdata_tlword[3]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[10]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[11]),
    .si1(net224),
    .si2(net225),
    .ssb(net314));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__12__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__13_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(net139),
    .d2(u_tlul_adapter_sram_rdata_tlword[5]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[12]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[13]),
    .si1(net226),
    .si2(net227),
    .ssb(net315));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__14__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__15_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[6]),
    .d2(u_tlul_adapter_sram_rdata_tlword[7]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[14]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[15]),
    .si1(net228),
    .si2(net229),
    .ssb(net316));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__16__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__17_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[8]),
    .d2(u_tlul_adapter_sram_rdata_tlword[9]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[16]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[17]),
    .si1(net230),
    .si2(net231),
    .ssb(net317));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__18__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__19_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(net138),
    .d2(u_tlul_adapter_sram_rdata_tlword[11]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[18]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[19]),
    .si1(net232),
    .si2(net233),
    .ssb(net318));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__20__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__21_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(net137),
    .d2(u_tlul_adapter_sram_rdata_tlword[13]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[20]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[21]),
    .si1(net234),
    .si2(net235),
    .ssb(net319));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__22__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__23_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[14]),
    .d2(u_tlul_adapter_sram_rdata_tlword[15]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[22]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[23]),
    .si1(net236),
    .si2(net237),
    .ssb(net320));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__24__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__25_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[16]),
    .d2(u_tlul_adapter_sram_rdata_tlword[17]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[24]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[25]),
    .si1(net238),
    .si2(net239),
    .ssb(net321));
 b15fpy000ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__26_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d(u_tlul_adapter_sram_rdata_tlword[18]),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[26]),
    .si(net240),
    .ssb(net322));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__27__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__28_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[19]),
    .d2(u_tlul_adapter_sram_rdata_tlword[20]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[27]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[28]),
    .si1(net241),
    .si2(net242),
    .ssb(net323));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__29__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__30_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[21]),
    .d2(u_tlul_adapter_sram_rdata_tlword[22]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[29]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[30]),
    .si1(net243),
    .si2(net244),
    .ssb(net324));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(net245),
    .d2(net246),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[2]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[3]),
    .si1(net247),
    .si2(net248),
    .ssb(net325));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__31__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__32_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[23]),
    .d2(u_tlul_adapter_sram_rdata_tlword[24]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[31]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[32]),
    .si1(net249),
    .si2(net250),
    .ssb(net326));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__33__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__34_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[25]),
    .d2(u_tlul_adapter_sram_rdata_tlword[26]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[33]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[34]),
    .si1(net251),
    .si2(net252),
    .ssb(net327));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__35__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__36_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[27]),
    .d2(u_tlul_adapter_sram_rdata_tlword[28]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[35]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[36]),
    .si1(net253),
    .si2(net254),
    .ssb(net328));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__37__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__38_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d1(u_tlul_adapter_sram_rdata_tlword[29]),
    .d2(u_tlul_adapter_sram_rdata_tlword[30]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[37]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[38]),
    .si1(net255),
    .si2(net256),
    .ssb(net329));
 b15fpy000ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__39_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622),
    .d(u_tlul_adapter_sram_rdata_tlword[31]),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[39]),
    .si(net257),
    .ssb(net330));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(net258),
    .d2(net259),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[4]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[5]),
    .si1(net260),
    .si2(net261),
    .ssb(net331));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7_ (.clk(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(net262),
    .d2(net263),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[6]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[7]),
    .si1(net264),
    .si2(net265),
    .ssb(net332));
 b15fpy200ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__8__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__9_ (.clk(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net616),
    .d1(net141),
    .d2(u_tlul_adapter_sram_rdata_tlword[1]),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[8]),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[9]),
    .si1(net266),
    .si2(net267),
    .ssb(net333));
 b15fqy203ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0_ (.rb(net176),
    .clk(clknet_1_1__leaf_clk_i),
    .d1(n131),
    .d2(n126),
    .o1(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_rptr_value_0_),
    .o2(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_wptr_value_0_),
    .si1(net268),
    .si2(net269),
    .ssb(net334));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N25),
    .den(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_rptr_1_),
    .rb(net5),
    .si(net270),
    .ssb(net335));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N11),
    .den(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_wptr_1_),
    .rb(net5),
    .si(net271),
    .ssb(net336));
 b15fqy00car1n02x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst_reg (.clk(clknet_1_1__leaf_clk_i),
    .d(net272),
    .o(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst),
    .psb(net176),
    .si(net273),
    .ssb(net337));
 b15fpy000ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__0_ (.clk(clknet_1_1__leaf_clk_i),
    .d(n189),
    .o(n188),
    .si(net274),
    .ssb(net338));
 b15fpy040ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__1_ (.clk(clknet_1_1__leaf_clk_i),
    .d(net177),
    .den(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[1]),
    .si(net275),
    .ssb(net339));
 b15fpy040ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__2_ (.clk(clknet_1_1__leaf_clk_i),
    .d(net175),
    .den(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[2]),
    .si(net276),
    .ssb(net340));
 b15fpy040ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__3_ (.clk(clknet_1_1__leaf_clk_i),
    .d(net51),
    .den(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[3]),
    .si(net277),
    .ssb(net341));
 b15fpy040ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__4_ (.clk(clknet_1_1__leaf_clk_i),
    .d(net52),
    .den(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[4]),
    .si(net278),
    .ssb(net342));
 b15fqy203ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0_ (.rb(net176),
    .clk(clknet_1_0__leaf_clk_i),
    .d1(n175),
    .d2(n192),
    .o1(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_rptr_value_0_),
    .o2(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_wptr_value_0_),
    .si1(net279),
    .si2(net280),
    .ssb(net343));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N25),
    .den(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N23),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_rptr_1_),
    .rb(net5),
    .si(net281),
    .ssb(net344));
 b15fqy043ar1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1_ (.clk(clknet_1_0__leaf_clk_i),
    .d(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N11),
    .den(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_wptr_1_),
    .rb(net5),
    .si(net282),
    .ssb(net345));
 b15fqy00car1n02x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst_reg (.clk(clknet_1_1__leaf_clk_i),
    .d(net283),
    .o(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst),
    .psb(net176),
    .si(net284),
    .ssb(net346));
 b15tihi00an1n03x5 U585_285 (.o(net285));
 b15cbf000an1n16x5 clkbuf_0_clk_i (.clk(net347),
    .clkout(clknet_0_clk_i));
 b15ztpn00an1n08x5 PHY_6 ();
 b15ztpn00an1n08x5 PHY_7 ();
 b15ztpn00an1n08x5 PHY_8 ();
 b15ztpn00an1n08x5 PHY_9 ();
 b15ztpn00an1n08x5 PHY_10 ();
 b15ztpn00an1n08x5 PHY_11 ();
 b15ztpn00an1n08x5 PHY_12 ();
 b15ztpn00an1n08x5 PHY_13 ();
 b15ztpn00an1n08x5 PHY_14 ();
 b15ztpn00an1n08x5 PHY_15 ();
 b15ztpn00an1n08x5 PHY_16 ();
 b15ztpn00an1n08x5 PHY_17 ();
 b15ztpn00an1n08x5 PHY_18 ();
 b15ztpn00an1n08x5 PHY_19 ();
 b15ztpn00an1n08x5 PHY_20 ();
 b15ztpn00an1n08x5 PHY_21 ();
 b15ztpn00an1n08x5 PHY_22 ();
 b15ztpn00an1n08x5 PHY_23 ();
 b15ztpn00an1n08x5 PHY_24 ();
 b15ztpn00an1n08x5 PHY_25 ();
 b15ztpn00an1n08x5 PHY_26 ();
 b15ztpn00an1n08x5 PHY_27 ();
 b15ztpn00an1n08x5 PHY_28 ();
 b15ztpn00an1n08x5 PHY_29 ();
 b15ztpn00an1n08x5 PHY_30 ();
 b15ztpn00an1n08x5 PHY_31 ();
 b15ztpn00an1n08x5 PHY_32 ();
 b15ztpn00an1n08x5 PHY_33 ();
 b15ztpn00an1n08x5 PHY_34 ();
 b15ztpn00an1n08x5 PHY_35 ();
 b15ztpn00an1n08x5 PHY_36 ();
 b15ztpn00an1n08x5 PHY_37 ();
 b15ztpn00an1n08x5 PHY_38 ();
 b15ztpn00an1n08x5 PHY_39 ();
 b15ztpn00an1n08x5 PHY_40 ();
 b15ztpn00an1n08x5 PHY_41 ();
 b15ztpn00an1n08x5 PHY_42 ();
 b15ztpn00an1n08x5 PHY_43 ();
 b15ztpn00an1n08x5 PHY_44 ();
 b15ztpn00an1n08x5 PHY_45 ();
 b15ztpn00an1n08x5 PHY_46 ();
 b15ztpn00an1n08x5 PHY_47 ();
 b15ztpn00an1n08x5 PHY_48 ();
 b15ztpn00an1n08x5 PHY_49 ();
 b15ztpn00an1n08x5 PHY_50 ();
 b15ztpn00an1n08x5 PHY_51 ();
 b15ztpn00an1n08x5 PHY_52 ();
 b15ztpn00an1n08x5 PHY_53 ();
 b15ztpn00an1n08x5 PHY_54 ();
 b15ztpn00an1n08x5 PHY_55 ();
 b15ztpn00an1n08x5 PHY_56 ();
 b15ztpn00an1n08x5 PHY_57 ();
 b15ztpn00an1n08x5 PHY_58 ();
 b15ztpn00an1n08x5 PHY_59 ();
 b15ztpn00an1n08x5 PHY_60 ();
 b15ztpn00an1n08x5 PHY_61 ();
 b15ztpn00an1n08x5 PHY_62 ();
 b15ztpn00an1n08x5 PHY_63 ();
 b15ztpn00an1n08x5 PHY_64 ();
 b15ztpn00an1n08x5 PHY_65 ();
 b15ztpn00an1n08x5 PHY_66 ();
 b15ztpn00an1n08x5 PHY_67 ();
 b15ztpn00an1n08x5 PHY_68 ();
 b15ztpn00an1n08x5 PHY_69 ();
 b15ztpn00an1n08x5 PHY_70 ();
 b15ztpn00an1n08x5 PHY_71 ();
 b15ztpn00an1n08x5 PHY_72 ();
 b15ztpn00an1n08x5 PHY_73 ();
 b15ztpn00an1n08x5 PHY_74 ();
 b15ztpn00an1n08x5 PHY_75 ();
 b15ztpn00an1n08x5 PHY_76 ();
 b15ztpn00an1n08x5 PHY_77 ();
 b15ztpn00an1n08x5 PHY_78 ();
 b15ztpn00an1n08x5 PHY_79 ();
 b15ztpn00an1n08x5 PHY_80 ();
 b15ztpn00an1n08x5 PHY_81 ();
 b15ztpn00an1n08x5 PHY_82 ();
 b15ztpn00an1n08x5 PHY_83 ();
 b15ztpn00an1n08x5 PHY_84 ();
 b15ztpn00an1n08x5 PHY_85 ();
 b15ztpn00an1n08x5 PHY_86 ();
 b15ztpn00an1n08x5 PHY_87 ();
 b15ztpn00an1n08x5 PHY_88 ();
 b15ztpn00an1n08x5 PHY_89 ();
 b15ztpn00an1n08x5 PHY_90 ();
 b15ztpn00an1n08x5 PHY_91 ();
 b15ztpn00an1n08x5 PHY_92 ();
 b15ztpn00an1n08x5 PHY_93 ();
 b15ztpn00an1n08x5 PHY_94 ();
 b15ztpn00an1n08x5 PHY_95 ();
 b15ztpn00an1n08x5 PHY_96 ();
 b15ztpn00an1n08x5 PHY_97 ();
 b15ztpn00an1n08x5 PHY_98 ();
 b15ztpn00an1n08x5 PHY_99 ();
 b15ztpn00an1n08x5 PHY_100 ();
 b15ztpn00an1n08x5 PHY_101 ();
 b15ztpn00an1n08x5 PHY_102 ();
 b15ztpn00an1n08x5 PHY_103 ();
 b15ztpn00an1n08x5 PHY_104 ();
 b15ztpn00an1n08x5 PHY_105 ();
 b15ztpn00an1n08x5 PHY_106 ();
 b15ztpn00an1n08x5 PHY_107 ();
 b15ztpn00an1n08x5 PHY_108 ();
 b15ztpn00an1n08x5 PHY_109 ();
 b15ztpn00an1n08x5 PHY_110 ();
 b15ztpn00an1n08x5 PHY_111 ();
 b15ztpn00an1n08x5 PHY_112 ();
 b15ztpn00an1n08x5 PHY_113 ();
 b15ztpn00an1n08x5 PHY_114 ();
 b15ztpn00an1n08x5 PHY_115 ();
 b15ztpn00an1n08x5 PHY_116 ();
 b15ztpn00an1n08x5 PHY_117 ();
 b15ztpn00an1n08x5 PHY_118 ();
 b15ztpn00an1n08x5 PHY_119 ();
 b15ztpn00an1n08x5 PHY_120 ();
 b15ztpn00an1n08x5 PHY_121 ();
 b15ztpn00an1n08x5 PHY_122 ();
 b15ztpn00an1n08x5 PHY_123 ();
 b15ztpn00an1n08x5 PHY_124 ();
 b15ztpn00an1n08x5 PHY_125 ();
 b15ztpn00an1n08x5 PHY_126 ();
 b15ztpn00an1n08x5 PHY_127 ();
 b15ztpn00an1n08x5 PHY_128 ();
 b15ztpn00an1n08x5 PHY_129 ();
 b15ztpn00an1n08x5 PHY_130 ();
 b15ztpn00an1n08x5 PHY_131 ();
 b15ztpn00an1n08x5 PHY_132 ();
 b15ztpn00an1n08x5 PHY_133 ();
 b15ztpn00an1n08x5 PHY_134 ();
 b15ztpn00an1n08x5 PHY_135 ();
 b15ztpn00an1n08x5 PHY_136 ();
 b15ztpn00an1n08x5 PHY_137 ();
 b15ztpn00an1n08x5 PHY_138 ();
 b15ztpn00an1n08x5 PHY_139 ();
 b15ztpn00an1n08x5 PHY_140 ();
 b15ztpn00an1n08x5 PHY_141 ();
 b15ztpn00an1n08x5 PHY_142 ();
 b15ztpn00an1n08x5 PHY_143 ();
 b15ztpn00an1n08x5 PHY_144 ();
 b15ztpn00an1n08x5 PHY_145 ();
 b15ztpn00an1n08x5 PHY_146 ();
 b15ztpn00an1n08x5 PHY_147 ();
 b15ztpn00an1n08x5 PHY_148 ();
 b15ztpn00an1n08x5 PHY_149 ();
 b15ztpn00an1n08x5 PHY_150 ();
 b15ztpn00an1n08x5 PHY_151 ();
 b15ztpn00an1n08x5 PHY_152 ();
 b15ztpn00an1n08x5 PHY_153 ();
 b15ztpn00an1n08x5 PHY_154 ();
 b15ztpn00an1n08x5 PHY_155 ();
 b15ztpn00an1n08x5 PHY_156 ();
 b15ztpn00an1n08x5 PHY_157 ();
 b15ztpn00an1n08x5 PHY_158 ();
 b15ztpn00an1n08x5 PHY_159 ();
 b15ztpn00an1n08x5 PHY_160 ();
 b15ztpn00an1n08x5 PHY_161 ();
 b15ztpn00an1n08x5 PHY_162 ();
 b15ztpn00an1n08x5 PHY_163 ();
 b15ztpn00an1n08x5 PHY_164 ();
 b15ztpn00an1n08x5 PHY_165 ();
 b15ztpn00an1n08x5 PHY_166 ();
 b15ztpn00an1n08x5 PHY_167 ();
 b15ztpn00an1n08x5 PHY_168 ();
 b15ztpn00an1n08x5 PHY_169 ();
 b15ztpn00an1n08x5 PHY_170 ();
 b15ztpn00an1n08x5 PHY_171 ();
 b15ztpn00an1n08x5 PHY_172 ();
 b15ztpn00an1n08x5 PHY_173 ();
 b15ztpn00an1n08x5 PHY_174 ();
 b15ztpn00an1n08x5 PHY_175 ();
 b15ztpn00an1n08x5 PHY_176 ();
 b15ztpn00an1n08x5 PHY_177 ();
 b15ztpn00an1n08x5 PHY_178 ();
 b15ztpn00an1n08x5 PHY_179 ();
 b15ztpn00an1n08x5 PHY_180 ();
 b15ztpn00an1n08x5 PHY_181 ();
 b15ztpn00an1n08x5 PHY_182 ();
 b15ztpn00an1n08x5 PHY_183 ();
 b15ztpn00an1n08x5 PHY_184 ();
 b15ztpn00an1n08x5 PHY_185 ();
 b15ztpn00an1n08x5 PHY_186 ();
 b15ztpn00an1n08x5 PHY_187 ();
 b15ztpn00an1n08x5 PHY_188 ();
 b15ztpn00an1n08x5 PHY_189 ();
 b15ztpn00an1n08x5 PHY_190 ();
 b15ztpn00an1n08x5 PHY_191 ();
 b15ztpn00an1n08x5 PHY_192 ();
 b15ztpn00an1n08x5 PHY_193 ();
 b15ztpn00an1n08x5 PHY_194 ();
 b15ztpn00an1n08x5 PHY_195 ();
 b15ztpn00an1n08x5 PHY_196 ();
 b15ztpn00an1n08x5 PHY_197 ();
 b15ztpn00an1n08x5 PHY_198 ();
 b15ztpn00an1n08x5 PHY_199 ();
 b15ztpn00an1n08x5 PHY_200 ();
 b15ztpn00an1n08x5 PHY_201 ();
 b15ztpn00an1n08x5 PHY_202 ();
 b15ztpn00an1n08x5 PHY_203 ();
 b15ztpn00an1n08x5 PHY_204 ();
 b15ztpn00an1n08x5 PHY_205 ();
 b15ztpn00an1n08x5 PHY_206 ();
 b15ztpn00an1n08x5 PHY_207 ();
 b15ztpn00an1n08x5 PHY_208 ();
 b15ztpn00an1n08x5 PHY_209 ();
 b15ztpn00an1n08x5 PHY_210 ();
 b15ztpn00an1n08x5 PHY_211 ();
 b15ztpn00an1n08x5 PHY_212 ();
 b15ztpn00an1n08x5 PHY_213 ();
 b15ztpn00an1n08x5 PHY_214 ();
 b15ztpn00an1n08x5 PHY_215 ();
 b15ztpn00an1n08x5 PHY_216 ();
 b15ztpn00an1n08x5 PHY_217 ();
 b15ztpn00an1n08x5 PHY_218 ();
 b15ztpn00an1n08x5 PHY_219 ();
 b15ztpn00an1n08x5 PHY_220 ();
 b15ztpn00an1n08x5 PHY_221 ();
 b15ztpn00an1n08x5 PHY_222 ();
 b15ztpn00an1n08x5 PHY_223 ();
 b15ztpn00an1n08x5 PHY_224 ();
 b15ztpn00an1n08x5 PHY_225 ();
 b15ztpn00an1n08x5 PHY_226 ();
 b15ztpn00an1n08x5 PHY_227 ();
 b15ztpn00an1n08x5 PHY_228 ();
 b15ztpn00an1n08x5 PHY_229 ();
 b15ztpn00an1n08x5 PHY_230 ();
 b15ztpn00an1n08x5 PHY_231 ();
 b15ztpn00an1n08x5 PHY_232 ();
 b15ztpn00an1n08x5 PHY_233 ();
 b15ztpn00an1n08x5 PHY_234 ();
 b15ztpn00an1n08x5 PHY_235 ();
 b15ztpn00an1n08x5 PHY_236 ();
 b15ztpn00an1n08x5 PHY_237 ();
 b15ztpn00an1n08x5 PHY_238 ();
 b15ztpn00an1n08x5 PHY_239 ();
 b15ztpn00an1n08x5 PHY_240 ();
 b15ztpn00an1n08x5 PHY_241 ();
 b15ztpn00an1n08x5 PHY_242 ();
 b15ztpn00an1n08x5 PHY_243 ();
 b15ztpn00an1n08x5 PHY_244 ();
 b15ztpn00an1n08x5 PHY_245 ();
 b15ztpn00an1n08x5 PHY_246 ();
 b15ztpn00an1n08x5 PHY_247 ();
 b15ztpn00an1n08x5 PHY_248 ();
 b15ztpn00an1n08x5 PHY_249 ();
 b15ztpn00an1n08x5 PHY_250 ();
 b15ztpn00an1n08x5 PHY_251 ();
 b15ztpn00an1n08x5 PHY_252 ();
 b15ztpn00an1n08x5 PHY_253 ();
 b15ztpn00an1n08x5 PHY_254 ();
 b15ztpn00an1n08x5 PHY_255 ();
 b15ztpn00an1n08x5 PHY_256 ();
 b15ztpn00an1n08x5 PHY_257 ();
 b15ztpn00an1n08x5 PHY_258 ();
 b15ztpn00an1n08x5 PHY_259 ();
 b15ztpn00an1n08x5 PHY_260 ();
 b15ztpn00an1n08x5 PHY_261 ();
 b15ztpn00an1n08x5 PHY_262 ();
 b15ztpn00an1n08x5 PHY_263 ();
 b15ztpn00an1n08x5 PHY_264 ();
 b15ztpn00an1n08x5 PHY_265 ();
 b15ztpn00an1n08x5 PHY_266 ();
 b15ztpn00an1n08x5 PHY_267 ();
 b15ztpn00an1n08x5 PHY_268 ();
 b15ztpn00an1n08x5 PHY_269 ();
 b15ztpn00an1n08x5 PHY_270 ();
 b15ztpn00an1n08x5 PHY_271 ();
 b15ztpn00an1n08x5 PHY_272 ();
 b15ztpn00an1n08x5 PHY_273 ();
 b15ztpn00an1n08x5 PHY_274 ();
 b15ztpn00an1n08x5 PHY_275 ();
 b15ztpn00an1n08x5 PHY_276 ();
 b15ztpn00an1n08x5 PHY_277 ();
 b15ztpn00an1n08x5 PHY_278 ();
 b15ztpn00an1n08x5 PHY_279 ();
 b15ztpn00an1n08x5 PHY_280 ();
 b15ztpn00an1n08x5 PHY_281 ();
 b15ztpn00an1n08x5 PHY_282 ();
 b15ztpn00an1n08x5 PHY_283 ();
 b15ztpn00an1n08x5 PHY_284 ();
 b15ztpn00an1n08x5 PHY_285 ();
 b15ztpn00an1n08x5 PHY_286 ();
 b15ztpn00an1n08x5 PHY_287 ();
 b15ztpn00an1n08x5 PHY_288 ();
 b15ztpn00an1n08x5 PHY_289 ();
 b15ztpn00an1n08x5 PHY_290 ();
 b15ztpn00an1n08x5 PHY_291 ();
 b15ztpn00an1n08x5 PHY_292 ();
 b15ztpn00an1n08x5 PHY_293 ();
 b15ztpn00an1n08x5 PHY_294 ();
 b15ztpn00an1n08x5 PHY_295 ();
 b15ztpn00an1n08x5 PHY_296 ();
 b15ztpn00an1n08x5 PHY_297 ();
 b15ztpn00an1n08x5 PHY_298 ();
 b15ztpn00an1n08x5 PHY_299 ();
 b15ztpn00an1n08x5 PHY_300 ();
 b15ztpn00an1n08x5 PHY_301 ();
 b15ztpn00an1n08x5 PHY_302 ();
 b15ztpn00an1n08x5 PHY_303 ();
 b15ztpn00an1n08x5 PHY_304 ();
 b15ztpn00an1n08x5 PHY_305 ();
 b15ztpn00an1n08x5 PHY_306 ();
 b15ztpn00an1n08x5 PHY_307 ();
 b15ztpn00an1n08x5 PHY_308 ();
 b15ztpn00an1n08x5 PHY_309 ();
 b15ztpn00an1n08x5 PHY_310 ();
 b15ztpn00an1n08x5 PHY_311 ();
 b15ztpn00an1n08x5 PHY_312 ();
 b15ztpn00an1n08x5 PHY_313 ();
 b15ztpn00an1n08x5 PHY_314 ();
 b15ztpn00an1n08x5 PHY_315 ();
 b15ztpn00an1n08x5 PHY_316 ();
 b15ztpn00an1n08x5 PHY_317 ();
 b15ztpn00an1n08x5 PHY_318 ();
 b15ztpn00an1n08x5 PHY_319 ();
 b15ztpn00an1n08x5 PHY_320 ();
 b15ztpn00an1n08x5 PHY_321 ();
 b15ztpn00an1n08x5 PHY_322 ();
 b15ztpn00an1n08x5 PHY_323 ();
 b15ztpn00an1n08x5 PHY_324 ();
 b15ztpn00an1n08x5 PHY_325 ();
 b15ztpn00an1n08x5 PHY_326 ();
 b15ztpn00an1n08x5 PHY_327 ();
 b15ztpn00an1n08x5 PHY_328 ();
 b15ztpn00an1n08x5 PHY_329 ();
 b15ztpn00an1n08x5 PHY_330 ();
 b15ztpn00an1n08x5 PHY_331 ();
 b15ztpn00an1n08x5 PHY_332 ();
 b15ztpn00an1n08x5 PHY_333 ();
 b15ztpn00an1n08x5 PHY_334 ();
 b15ztpn00an1n08x5 PHY_335 ();
 b15ztpn00an1n08x5 PHY_336 ();
 b15ztpn00an1n08x5 PHY_337 ();
 b15ztpn00an1n08x5 PHY_338 ();
 b15ztpn00an1n08x5 PHY_339 ();
 b15ztpn00an1n08x5 PHY_340 ();
 b15ztpn00an1n08x5 PHY_341 ();
 b15ztpn00an1n08x5 PHY_342 ();
 b15ztpn00an1n08x5 PHY_343 ();
 b15ztpn00an1n08x5 PHY_344 ();
 b15ztpn00an1n08x5 PHY_345 ();
 b15ztpn00an1n08x5 PHY_346 ();
 b15ztpn00an1n08x5 PHY_347 ();
 b15ztpn00an1n08x5 PHY_348 ();
 b15ztpn00an1n08x5 PHY_349 ();
 b15ztpn00an1n08x5 PHY_350 ();
 b15ztpn00an1n08x5 PHY_351 ();
 b15ztpn00an1n08x5 PHY_352 ();
 b15ztpn00an1n08x5 PHY_353 ();
 b15ztpn00an1n08x5 PHY_354 ();
 b15ztpn00an1n08x5 PHY_355 ();
 b15ztpn00an1n08x5 PHY_356 ();
 b15ztpn00an1n08x5 PHY_357 ();
 b15ztpn00an1n08x5 PHY_358 ();
 b15ztpn00an1n08x5 PHY_359 ();
 b15ztpn00an1n08x5 PHY_360 ();
 b15ztpn00an1n08x5 PHY_361 ();
 b15ztpn00an1n08x5 PHY_362 ();
 b15ztpn00an1n08x5 PHY_363 ();
 b15ztpn00an1n08x5 PHY_364 ();
 b15ztpn00an1n08x5 PHY_365 ();
 b15ztpn00an1n08x5 PHY_366 ();
 b15ztpn00an1n08x5 PHY_367 ();
 b15ztpn00an1n08x5 PHY_368 ();
 b15ztpn00an1n08x5 PHY_369 ();
 b15ztpn00an1n08x5 PHY_370 ();
 b15ztpn00an1n08x5 PHY_371 ();
 b15ztpn00an1n08x5 PHY_372 ();
 b15ztpn00an1n08x5 PHY_373 ();
 b15ztpn00an1n08x5 PHY_374 ();
 b15ztpn00an1n08x5 PHY_375 ();
 b15ztpn00an1n08x5 PHY_376 ();
 b15ztpn00an1n08x5 PHY_377 ();
 b15ztpn00an1n08x5 PHY_378 ();
 b15ztpn00an1n08x5 PHY_379 ();
 b15ztpn00an1n08x5 PHY_380 ();
 b15ztpn00an1n08x5 PHY_381 ();
 b15ztpn00an1n08x5 PHY_382 ();
 b15ztpn00an1n08x5 PHY_383 ();
 b15ztpn00an1n08x5 PHY_384 ();
 b15ztpn00an1n08x5 PHY_385 ();
 b15ztpn00an1n08x5 PHY_386 ();
 b15ztpn00an1n08x5 PHY_387 ();
 b15ztpn00an1n08x5 PHY_388 ();
 b15ztpn00an1n08x5 PHY_389 ();
 b15ztpn00an1n08x5 PHY_390 ();
 b15ztpn00an1n08x5 PHY_391 ();
 b15ztpn00an1n08x5 PHY_392 ();
 b15ztpn00an1n08x5 PHY_393 ();
 b15ztpn00an1n08x5 PHY_394 ();
 b15ztpn00an1n08x5 PHY_395 ();
 b15ztpn00an1n08x5 PHY_396 ();
 b15ztpn00an1n08x5 PHY_397 ();
 b15ztpn00an1n08x5 PHY_398 ();
 b15ztpn00an1n08x5 PHY_399 ();
 b15ztpn00an1n08x5 PHY_400 ();
 b15ztpn00an1n08x5 PHY_401 ();
 b15ztpn00an1n08x5 PHY_402 ();
 b15ztpn00an1n08x5 PHY_403 ();
 b15ztpn00an1n08x5 PHY_404 ();
 b15ztpn00an1n08x5 PHY_405 ();
 b15ztpn00an1n08x5 PHY_406 ();
 b15ztpn00an1n08x5 PHY_407 ();
 b15ztpn00an1n08x5 PHY_408 ();
 b15ztpn00an1n08x5 PHY_409 ();
 b15ztpn00an1n08x5 PHY_410 ();
 b15ztpn00an1n08x5 PHY_411 ();
 b15ztpn00an1n08x5 PHY_412 ();
 b15ztpn00an1n08x5 PHY_413 ();
 b15ztpn00an1n08x5 PHY_414 ();
 b15ztpn00an1n08x5 PHY_415 ();
 b15ztpn00an1n08x5 PHY_416 ();
 b15ztpn00an1n08x5 PHY_417 ();
 b15ztpn00an1n08x5 PHY_418 ();
 b15ztpn00an1n08x5 PHY_419 ();
 b15ztpn00an1n08x5 PHY_420 ();
 b15ztpn00an1n08x5 PHY_421 ();
 b15ztpn00an1n08x5 PHY_422 ();
 b15ztpn00an1n08x5 PHY_423 ();
 b15ztpn00an1n08x5 PHY_424 ();
 b15ztpn00an1n08x5 PHY_425 ();
 b15ztpn00an1n08x5 PHY_426 ();
 b15ztpn00an1n08x5 PHY_427 ();
 b15ztpn00an1n08x5 PHY_428 ();
 b15ztpn00an1n08x5 PHY_429 ();
 b15ztpn00an1n08x5 PHY_430 ();
 b15ztpn00an1n08x5 PHY_431 ();
 b15ztpn00an1n08x5 PHY_432 ();
 b15ztpn00an1n08x5 PHY_433 ();
 b15ztpn00an1n08x5 PHY_434 ();
 b15ztpn00an1n08x5 PHY_435 ();
 b15ztpn00an1n08x5 PHY_436 ();
 b15ztpn00an1n08x5 PHY_437 ();
 b15ztpn00an1n08x5 PHY_438 ();
 b15ztpn00an1n08x5 PHY_439 ();
 b15ztpn00an1n08x5 PHY_440 ();
 b15ztpn00an1n08x5 PHY_441 ();
 b15ztpn00an1n08x5 PHY_442 ();
 b15ztpn00an1n08x5 PHY_443 ();
 b15ztpn00an1n08x5 PHY_444 ();
 b15ztpn00an1n08x5 PHY_445 ();
 b15ztpn00an1n08x5 PHY_446 ();
 b15ztpn00an1n08x5 PHY_447 ();
 b15ztpn00an1n08x5 PHY_448 ();
 b15ztpn00an1n08x5 PHY_449 ();
 b15ztpn00an1n08x5 PHY_450 ();
 b15ztpn00an1n08x5 PHY_451 ();
 b15ztpn00an1n08x5 PHY_452 ();
 b15ztpn00an1n08x5 PHY_453 ();
 b15ztpn00an1n08x5 PHY_454 ();
 b15ztpn00an1n08x5 PHY_455 ();
 b15ztpn00an1n08x5 PHY_456 ();
 b15ztpn00an1n08x5 PHY_457 ();
 b15ztpn00an1n08x5 PHY_458 ();
 b15ztpn00an1n08x5 PHY_459 ();
 b15ztpn00an1n08x5 PHY_460 ();
 b15ztpn00an1n08x5 PHY_461 ();
 b15ztpn00an1n08x5 PHY_462 ();
 b15ztpn00an1n08x5 PHY_463 ();
 b15ztpn00an1n08x5 PHY_464 ();
 b15ztpn00an1n08x5 PHY_465 ();
 b15ztpn00an1n08x5 PHY_466 ();
 b15ztpn00an1n08x5 PHY_467 ();
 b15ztpn00an1n08x5 PHY_468 ();
 b15ztpn00an1n08x5 PHY_469 ();
 b15ztpn00an1n08x5 PHY_470 ();
 b15ztpn00an1n08x5 PHY_471 ();
 b15ztpn00an1n08x5 PHY_472 ();
 b15ztpn00an1n08x5 PHY_473 ();
 b15ztpn00an1n08x5 PHY_474 ();
 b15ztpn00an1n08x5 PHY_475 ();
 b15ztpn00an1n08x5 PHY_476 ();
 b15ztpn00an1n08x5 PHY_477 ();
 b15ztpn00an1n08x5 PHY_478 ();
 b15ztpn00an1n08x5 PHY_479 ();
 b15ztpn00an1n08x5 PHY_480 ();
 b15ztpn00an1n08x5 PHY_481 ();
 b15ztpn00an1n08x5 PHY_482 ();
 b15ztpn00an1n08x5 PHY_483 ();
 b15ztpn00an1n08x5 PHY_484 ();
 b15ztpn00an1n08x5 PHY_485 ();
 b15ztpn00an1n08x5 PHY_486 ();
 b15ztpn00an1n08x5 PHY_487 ();
 b15ztpn00an1n08x5 PHY_488 ();
 b15ztpn00an1n08x5 PHY_489 ();
 b15ztpn00an1n08x5 PHY_490 ();
 b15ztpn00an1n08x5 PHY_491 ();
 b15ztpn00an1n08x5 PHY_492 ();
 b15ztpn00an1n08x5 PHY_493 ();
 b15ztpn00an1n08x5 PHY_494 ();
 b15ztpn00an1n08x5 PHY_495 ();
 b15ztpn00an1n08x5 PHY_496 ();
 b15ztpn00an1n08x5 PHY_497 ();
 b15ztpn00an1n08x5 PHY_498 ();
 b15ztpn00an1n08x5 PHY_499 ();
 b15ztpn00an1n08x5 PHY_500 ();
 b15ztpn00an1n08x5 PHY_501 ();
 b15ztpn00an1n08x5 PHY_502 ();
 b15ztpn00an1n08x5 PHY_503 ();
 b15ztpn00an1n08x5 PHY_504 ();
 b15ztpn00an1n08x5 PHY_505 ();
 b15ztpn00an1n08x5 PHY_506 ();
 b15ztpn00an1n08x5 PHY_507 ();
 b15ztpn00an1n08x5 PHY_508 ();
 b15ztpn00an1n08x5 PHY_509 ();
 b15ztpn00an1n08x5 PHY_510 ();
 b15ztpn00an1n08x5 PHY_511 ();
 b15ztpn00an1n08x5 PHY_512 ();
 b15ztpn00an1n08x5 PHY_513 ();
 b15ztpn00an1n08x5 PHY_514 ();
 b15ztpn00an1n08x5 PHY_515 ();
 b15ztpn00an1n08x5 PHY_516 ();
 b15ztpn00an1n08x5 PHY_517 ();
 b15ztpn00an1n08x5 PHY_518 ();
 b15ztpn00an1n08x5 PHY_519 ();
 b15ztpn00an1n08x5 PHY_520 ();
 b15ztpn00an1n08x5 PHY_521 ();
 b15ztpn00an1n08x5 PHY_522 ();
 b15ztpn00an1n08x5 PHY_523 ();
 b15ztpn00an1n08x5 PHY_524 ();
 b15ztpn00an1n08x5 PHY_525 ();
 b15ztpn00an1n08x5 PHY_526 ();
 b15ztpn00an1n08x5 PHY_527 ();
 b15ztpn00an1n08x5 PHY_528 ();
 b15ztpn00an1n08x5 PHY_529 ();
 b15ztpn00an1n08x5 PHY_530 ();
 b15ztpn00an1n08x5 PHY_531 ();
 b15ztpn00an1n08x5 PHY_532 ();
 b15ztpn00an1n08x5 PHY_533 ();
 b15ztpn00an1n08x5 PHY_534 ();
 b15ztpn00an1n08x5 PHY_535 ();
 b15ztpn00an1n08x5 PHY_536 ();
 b15ztpn00an1n08x5 PHY_537 ();
 b15ztpn00an1n08x5 PHY_538 ();
 b15ztpn00an1n08x5 PHY_539 ();
 b15ztpn00an1n08x5 PHY_540 ();
 b15ztpn00an1n08x5 PHY_541 ();
 b15ztpn00an1n08x5 PHY_542 ();
 b15ztpn00an1n08x5 PHY_543 ();
 b15ztpn00an1n08x5 PHY_544 ();
 b15ztpn00an1n08x5 PHY_545 ();
 b15ztpn00an1n08x5 PHY_546 ();
 b15ztpn00an1n08x5 PHY_547 ();
 b15ztpn00an1n08x5 PHY_548 ();
 b15ztpn00an1n08x5 PHY_549 ();
 b15ztpn00an1n08x5 PHY_550 ();
 b15ztpn00an1n08x5 PHY_551 ();
 b15ztpn00an1n08x5 PHY_552 ();
 b15ztpn00an1n08x5 PHY_553 ();
 b15ztpn00an1n08x5 PHY_554 ();
 b15ztpn00an1n08x5 PHY_555 ();
 b15ztpn00an1n08x5 PHY_556 ();
 b15ztpn00an1n08x5 PHY_557 ();
 b15ztpn00an1n08x5 PHY_558 ();
 b15ztpn00an1n08x5 PHY_559 ();
 b15ztpn00an1n08x5 PHY_560 ();
 b15ztpn00an1n08x5 PHY_561 ();
 b15ztpn00an1n08x5 PHY_562 ();
 b15ztpn00an1n08x5 PHY_563 ();
 b15ztpn00an1n08x5 PHY_564 ();
 b15ztpn00an1n08x5 PHY_565 ();
 b15ztpn00an1n08x5 PHY_566 ();
 b15ztpn00an1n08x5 PHY_567 ();
 b15ztpn00an1n08x5 PHY_568 ();
 b15ztpn00an1n08x5 PHY_569 ();
 b15ztpn00an1n08x5 PHY_570 ();
 b15ztpn00an1n08x5 PHY_571 ();
 b15ztpn00an1n08x5 PHY_572 ();
 b15ztpn00an1n08x5 PHY_573 ();
 b15ztpn00an1n08x5 PHY_574 ();
 b15ztpn00an1n08x5 PHY_575 ();
 b15ztpn00an1n08x5 PHY_576 ();
 b15ztpn00an1n08x5 PHY_577 ();
 b15ztpn00an1n08x5 PHY_578 ();
 b15ztpn00an1n08x5 PHY_579 ();
 b15ztpn00an1n08x5 PHY_580 ();
 b15ztpn00an1n08x5 PHY_581 ();
 b15ztpn00an1n08x5 PHY_582 ();
 b15ztpn00an1n08x5 PHY_583 ();
 b15ztpn00an1n08x5 TAP_584 ();
 b15ztpn00an1n08x5 TAP_585 ();
 b15ztpn00an1n08x5 TAP_586 ();
 b15ztpn00an1n08x5 TAP_587 ();
 b15ztpn00an1n08x5 TAP_588 ();
 b15ztpn00an1n08x5 TAP_589 ();
 b15ztpn00an1n08x5 TAP_590 ();
 b15ztpn00an1n08x5 TAP_591 ();
 b15ztpn00an1n08x5 TAP_592 ();
 b15ztpn00an1n08x5 TAP_593 ();
 b15ztpn00an1n08x5 TAP_594 ();
 b15ztpn00an1n08x5 TAP_595 ();
 b15ztpn00an1n08x5 TAP_596 ();
 b15ztpn00an1n08x5 TAP_597 ();
 b15ztpn00an1n08x5 TAP_598 ();
 b15ztpn00an1n08x5 TAP_599 ();
 b15ztpn00an1n08x5 TAP_600 ();
 b15ztpn00an1n08x5 TAP_601 ();
 b15ztpn00an1n08x5 TAP_602 ();
 b15ztpn00an1n08x5 TAP_603 ();
 b15ztpn00an1n08x5 TAP_604 ();
 b15ztpn00an1n08x5 TAP_605 ();
 b15ztpn00an1n08x5 TAP_606 ();
 b15ztpn00an1n08x5 TAP_607 ();
 b15ztpn00an1n08x5 TAP_608 ();
 b15ztpn00an1n08x5 TAP_609 ();
 b15ztpn00an1n08x5 TAP_610 ();
 b15ztpn00an1n08x5 TAP_611 ();
 b15ztpn00an1n08x5 TAP_612 ();
 b15ztpn00an1n08x5 TAP_613 ();
 b15ztpn00an1n08x5 TAP_614 ();
 b15ztpn00an1n08x5 TAP_615 ();
 b15ztpn00an1n08x5 TAP_616 ();
 b15ztpn00an1n08x5 TAP_617 ();
 b15ztpn00an1n08x5 TAP_618 ();
 b15ztpn00an1n08x5 TAP_619 ();
 b15ztpn00an1n08x5 TAP_620 ();
 b15ztpn00an1n08x5 TAP_621 ();
 b15ztpn00an1n08x5 TAP_622 ();
 b15ztpn00an1n08x5 TAP_623 ();
 b15ztpn00an1n08x5 TAP_624 ();
 b15ztpn00an1n08x5 TAP_625 ();
 b15ztpn00an1n08x5 TAP_626 ();
 b15ztpn00an1n08x5 TAP_627 ();
 b15ztpn00an1n08x5 TAP_628 ();
 b15ztpn00an1n08x5 TAP_629 ();
 b15ztpn00an1n08x5 TAP_630 ();
 b15ztpn00an1n08x5 TAP_631 ();
 b15ztpn00an1n08x5 TAP_632 ();
 b15ztpn00an1n08x5 TAP_633 ();
 b15ztpn00an1n08x5 TAP_634 ();
 b15ztpn00an1n08x5 TAP_635 ();
 b15ztpn00an1n08x5 TAP_636 ();
 b15ztpn00an1n08x5 TAP_637 ();
 b15ztpn00an1n08x5 TAP_638 ();
 b15ztpn00an1n08x5 TAP_639 ();
 b15ztpn00an1n08x5 TAP_640 ();
 b15ztpn00an1n08x5 TAP_641 ();
 b15ztpn00an1n08x5 TAP_642 ();
 b15ztpn00an1n08x5 TAP_643 ();
 b15ztpn00an1n08x5 TAP_644 ();
 b15ztpn00an1n08x5 TAP_645 ();
 b15ztpn00an1n08x5 TAP_646 ();
 b15ztpn00an1n08x5 TAP_647 ();
 b15ztpn00an1n08x5 TAP_648 ();
 b15ztpn00an1n08x5 TAP_649 ();
 b15ztpn00an1n08x5 TAP_650 ();
 b15ztpn00an1n08x5 TAP_651 ();
 b15ztpn00an1n08x5 TAP_652 ();
 b15ztpn00an1n08x5 TAP_653 ();
 b15ztpn00an1n08x5 TAP_654 ();
 b15ztpn00an1n08x5 TAP_655 ();
 b15ztpn00an1n08x5 TAP_656 ();
 b15ztpn00an1n08x5 TAP_657 ();
 b15ztpn00an1n08x5 TAP_658 ();
 b15ztpn00an1n08x5 TAP_659 ();
 b15ztpn00an1n08x5 TAP_660 ();
 b15ztpn00an1n08x5 TAP_661 ();
 b15ztpn00an1n08x5 TAP_662 ();
 b15ztpn00an1n08x5 TAP_663 ();
 b15ztpn00an1n08x5 TAP_664 ();
 b15ztpn00an1n08x5 TAP_665 ();
 b15ztpn00an1n08x5 TAP_666 ();
 b15ztpn00an1n08x5 TAP_667 ();
 b15ztpn00an1n08x5 TAP_668 ();
 b15ztpn00an1n08x5 TAP_669 ();
 b15ztpn00an1n08x5 TAP_670 ();
 b15ztpn00an1n08x5 TAP_671 ();
 b15ztpn00an1n08x5 TAP_672 ();
 b15ztpn00an1n08x5 TAP_673 ();
 b15ztpn00an1n08x5 TAP_674 ();
 b15ztpn00an1n08x5 TAP_675 ();
 b15ztpn00an1n08x5 TAP_676 ();
 b15ztpn00an1n08x5 TAP_677 ();
 b15ztpn00an1n08x5 TAP_678 ();
 b15ztpn00an1n08x5 TAP_679 ();
 b15ztpn00an1n08x5 TAP_680 ();
 b15ztpn00an1n08x5 TAP_681 ();
 b15ztpn00an1n08x5 TAP_682 ();
 b15ztpn00an1n08x5 TAP_683 ();
 b15ztpn00an1n08x5 TAP_684 ();
 b15ztpn00an1n08x5 TAP_685 ();
 b15ztpn00an1n08x5 TAP_686 ();
 b15ztpn00an1n08x5 TAP_687 ();
 b15ztpn00an1n08x5 TAP_688 ();
 b15ztpn00an1n08x5 TAP_689 ();
 b15ztpn00an1n08x5 TAP_690 ();
 b15ztpn00an1n08x5 TAP_691 ();
 b15ztpn00an1n08x5 TAP_692 ();
 b15ztpn00an1n08x5 TAP_693 ();
 b15ztpn00an1n08x5 TAP_694 ();
 b15ztpn00an1n08x5 TAP_695 ();
 b15ztpn00an1n08x5 TAP_696 ();
 b15ztpn00an1n08x5 TAP_697 ();
 b15ztpn00an1n08x5 TAP_698 ();
 b15ztpn00an1n08x5 TAP_699 ();
 b15ztpn00an1n08x5 TAP_700 ();
 b15ztpn00an1n08x5 TAP_701 ();
 b15ztpn00an1n08x5 TAP_702 ();
 b15ztpn00an1n08x5 TAP_703 ();
 b15ztpn00an1n08x5 TAP_704 ();
 b15ztpn00an1n08x5 TAP_705 ();
 b15ztpn00an1n08x5 TAP_706 ();
 b15ztpn00an1n08x5 TAP_707 ();
 b15ztpn00an1n08x5 TAP_708 ();
 b15ztpn00an1n08x5 TAP_709 ();
 b15ztpn00an1n08x5 TAP_710 ();
 b15ztpn00an1n08x5 TAP_711 ();
 b15ztpn00an1n08x5 TAP_712 ();
 b15ztpn00an1n08x5 TAP_713 ();
 b15ztpn00an1n08x5 TAP_714 ();
 b15ztpn00an1n08x5 TAP_715 ();
 b15ztpn00an1n08x5 TAP_716 ();
 b15ztpn00an1n08x5 TAP_717 ();
 b15ztpn00an1n08x5 TAP_718 ();
 b15ztpn00an1n08x5 TAP_719 ();
 b15ztpn00an1n08x5 TAP_720 ();
 b15ztpn00an1n08x5 TAP_721 ();
 b15ztpn00an1n08x5 TAP_722 ();
 b15ztpn00an1n08x5 TAP_723 ();
 b15ztpn00an1n08x5 TAP_724 ();
 b15ztpn00an1n08x5 TAP_725 ();
 b15ztpn00an1n08x5 TAP_726 ();
 b15ztpn00an1n08x5 TAP_727 ();
 b15ztpn00an1n08x5 TAP_728 ();
 b15ztpn00an1n08x5 TAP_729 ();
 b15ztpn00an1n08x5 TAP_730 ();
 b15ztpn00an1n08x5 TAP_731 ();
 b15ztpn00an1n08x5 TAP_732 ();
 b15ztpn00an1n08x5 TAP_733 ();
 b15ztpn00an1n08x5 TAP_734 ();
 b15ztpn00an1n08x5 TAP_735 ();
 b15ztpn00an1n08x5 TAP_736 ();
 b15ztpn00an1n08x5 TAP_737 ();
 b15ztpn00an1n08x5 TAP_738 ();
 b15ztpn00an1n08x5 TAP_739 ();
 b15ztpn00an1n08x5 TAP_740 ();
 b15ztpn00an1n08x5 TAP_741 ();
 b15ztpn00an1n08x5 TAP_742 ();
 b15ztpn00an1n08x5 TAP_743 ();
 b15ztpn00an1n08x5 TAP_744 ();
 b15ztpn00an1n08x5 TAP_745 ();
 b15ztpn00an1n08x5 TAP_746 ();
 b15ztpn00an1n08x5 TAP_747 ();
 b15ztpn00an1n08x5 TAP_748 ();
 b15ztpn00an1n08x5 TAP_749 ();
 b15ztpn00an1n08x5 TAP_750 ();
 b15ztpn00an1n08x5 TAP_751 ();
 b15ztpn00an1n08x5 TAP_752 ();
 b15ztpn00an1n08x5 TAP_753 ();
 b15ztpn00an1n08x5 TAP_754 ();
 b15ztpn00an1n08x5 TAP_755 ();
 b15ztpn00an1n08x5 TAP_756 ();
 b15ztpn00an1n08x5 TAP_757 ();
 b15ztpn00an1n08x5 TAP_758 ();
 b15ztpn00an1n08x5 TAP_759 ();
 b15ztpn00an1n08x5 TAP_760 ();
 b15ztpn00an1n08x5 TAP_761 ();
 b15ztpn00an1n08x5 TAP_762 ();
 b15ztpn00an1n08x5 TAP_763 ();
 b15ztpn00an1n08x5 TAP_764 ();
 b15ztpn00an1n08x5 TAP_765 ();
 b15ztpn00an1n08x5 TAP_766 ();
 b15ztpn00an1n08x5 TAP_767 ();
 b15ztpn00an1n08x5 TAP_768 ();
 b15ztpn00an1n08x5 TAP_769 ();
 b15ztpn00an1n08x5 TAP_770 ();
 b15ztpn00an1n08x5 TAP_771 ();
 b15ztpn00an1n08x5 TAP_772 ();
 b15ztpn00an1n08x5 TAP_773 ();
 b15ztpn00an1n08x5 TAP_774 ();
 b15ztpn00an1n08x5 TAP_775 ();
 b15ztpn00an1n08x5 TAP_776 ();
 b15ztpn00an1n08x5 TAP_777 ();
 b15ztpn00an1n08x5 TAP_778 ();
 b15ztpn00an1n08x5 TAP_779 ();
 b15ztpn00an1n08x5 TAP_780 ();
 b15ztpn00an1n08x5 TAP_781 ();
 b15ztpn00an1n08x5 TAP_782 ();
 b15ztpn00an1n08x5 TAP_783 ();
 b15ztpn00an1n08x5 TAP_784 ();
 b15ztpn00an1n08x5 TAP_785 ();
 b15ztpn00an1n08x5 TAP_786 ();
 b15ztpn00an1n08x5 TAP_787 ();
 b15ztpn00an1n08x5 TAP_788 ();
 b15ztpn00an1n08x5 TAP_789 ();
 b15ztpn00an1n08x5 TAP_790 ();
 b15ztpn00an1n08x5 TAP_791 ();
 b15ztpn00an1n08x5 TAP_792 ();
 b15ztpn00an1n08x5 TAP_793 ();
 b15ztpn00an1n08x5 TAP_794 ();
 b15ztpn00an1n08x5 TAP_795 ();
 b15ztpn00an1n08x5 TAP_796 ();
 b15ztpn00an1n08x5 TAP_797 ();
 b15ztpn00an1n08x5 TAP_798 ();
 b15ztpn00an1n08x5 TAP_799 ();
 b15ztpn00an1n08x5 TAP_800 ();
 b15ztpn00an1n08x5 TAP_801 ();
 b15ztpn00an1n08x5 TAP_802 ();
 b15ztpn00an1n08x5 TAP_803 ();
 b15ztpn00an1n08x5 TAP_804 ();
 b15ztpn00an1n08x5 TAP_805 ();
 b15ztpn00an1n08x5 TAP_806 ();
 b15ztpn00an1n08x5 TAP_807 ();
 b15ztpn00an1n08x5 TAP_808 ();
 b15ztpn00an1n08x5 TAP_809 ();
 b15ztpn00an1n08x5 TAP_810 ();
 b15ztpn00an1n08x5 TAP_811 ();
 b15ztpn00an1n08x5 TAP_812 ();
 b15ztpn00an1n08x5 TAP_813 ();
 b15ztpn00an1n08x5 TAP_814 ();
 b15ztpn00an1n08x5 TAP_815 ();
 b15ztpn00an1n08x5 TAP_816 ();
 b15ztpn00an1n08x5 TAP_817 ();
 b15ztpn00an1n08x5 TAP_818 ();
 b15ztpn00an1n08x5 TAP_819 ();
 b15ztpn00an1n08x5 TAP_820 ();
 b15ztpn00an1n08x5 TAP_821 ();
 b15ztpn00an1n08x5 TAP_822 ();
 b15ztpn00an1n08x5 TAP_823 ();
 b15ztpn00an1n08x5 TAP_824 ();
 b15ztpn00an1n08x5 TAP_825 ();
 b15ztpn00an1n08x5 TAP_826 ();
 b15ztpn00an1n08x5 TAP_827 ();
 b15ztpn00an1n08x5 TAP_828 ();
 b15ztpn00an1n08x5 TAP_829 ();
 b15ztpn00an1n08x5 TAP_830 ();
 b15ztpn00an1n08x5 TAP_831 ();
 b15ztpn00an1n08x5 TAP_832 ();
 b15ztpn00an1n08x5 TAP_833 ();
 b15ztpn00an1n08x5 TAP_834 ();
 b15ztpn00an1n08x5 TAP_835 ();
 b15ztpn00an1n08x5 TAP_836 ();
 b15ztpn00an1n08x5 TAP_837 ();
 b15ztpn00an1n08x5 TAP_838 ();
 b15ztpn00an1n08x5 TAP_839 ();
 b15ztpn00an1n08x5 TAP_840 ();
 b15ztpn00an1n08x5 TAP_841 ();
 b15ztpn00an1n08x5 TAP_842 ();
 b15ztpn00an1n08x5 TAP_843 ();
 b15ztpn00an1n08x5 TAP_844 ();
 b15ztpn00an1n08x5 TAP_845 ();
 b15ztpn00an1n08x5 TAP_846 ();
 b15ztpn00an1n08x5 TAP_847 ();
 b15ztpn00an1n08x5 TAP_848 ();
 b15ztpn00an1n08x5 TAP_849 ();
 b15ztpn00an1n08x5 TAP_850 ();
 b15ztpn00an1n08x5 TAP_851 ();
 b15ztpn00an1n08x5 TAP_852 ();
 b15ztpn00an1n08x5 TAP_853 ();
 b15ztpn00an1n08x5 TAP_854 ();
 b15ztpn00an1n08x5 TAP_855 ();
 b15ztpn00an1n08x5 TAP_856 ();
 b15ztpn00an1n08x5 TAP_857 ();
 b15ztpn00an1n08x5 TAP_858 ();
 b15ztpn00an1n08x5 TAP_859 ();
 b15ztpn00an1n08x5 TAP_860 ();
 b15ztpn00an1n08x5 TAP_861 ();
 b15ztpn00an1n08x5 TAP_862 ();
 b15ztpn00an1n08x5 TAP_863 ();
 b15ztpn00an1n08x5 TAP_864 ();
 b15ztpn00an1n08x5 TAP_865 ();
 b15ztpn00an1n08x5 TAP_866 ();
 b15ztpn00an1n08x5 TAP_867 ();
 b15ztpn00an1n08x5 TAP_868 ();
 b15ztpn00an1n08x5 TAP_869 ();
 b15ztpn00an1n08x5 TAP_870 ();
 b15ztpn00an1n08x5 TAP_871 ();
 b15ztpn00an1n08x5 TAP_872 ();
 b15ztpn00an1n08x5 TAP_873 ();
 b15ztpn00an1n08x5 TAP_874 ();
 b15ztpn00an1n08x5 TAP_875 ();
 b15ztpn00an1n08x5 TAP_876 ();
 b15ztpn00an1n08x5 TAP_877 ();
 b15ztpn00an1n08x5 TAP_878 ();
 b15bfn000ah1n04x5 input1 (.a(en_ifetch_i[0]),
    .o(net1));
 b15bfn000as1n04x5 input2 (.a(en_ifetch_i[1]),
    .o(net2));
 b15bfn000as1n04x5 input3 (.a(en_ifetch_i[2]),
    .o(net3));
 b15bfn000ah1n04x5 input4 (.a(en_ifetch_i[3]),
    .o(net4));
 b15bfn001as1n48x5 input5 (.a(rst_ni),
    .o(net5));
 b15bfn000ah1n24x5 input6 (.a(tl_i[0]),
    .o(net6));
 b15bfn001as1n12x5 input7 (.a(tl_i[100]),
    .o(net7));
 b15bfn001as1n24x5 input8 (.a(tl_i[101]),
    .o(net8));
 b15bfn001as1n12x5 input9 (.a(tl_i[105]),
    .o(net9));
 b15bfn001as1n16x5 input10 (.a(tl_i[106]),
    .o(net10));
 b15bfn001ah1n16x5 input11 (.a(tl_i[107]),
    .o(net11));
 b15bfn001ah1n24x5 input12 (.a(tl_i[108]),
    .o(net12));
 b15bfn001ah1n24x5 input13 (.a(tl_i[15]),
    .o(net13));
 b15bfn001ah1n24x5 input14 (.a(tl_i[16]),
    .o(net14));
 b15bfn001as1n12x5 input15 (.a(tl_i[17]),
    .o(net15));
 b15bfn001ah1n24x5 input16 (.a(tl_i[18]),
    .o(net16));
 b15bfn000ah1n06x5 input17 (.a(tl_i[24]),
    .o(net17));
 b15bfn001as1n06x5 input18 (.a(tl_i[25]),
    .o(net18));
 b15bfn000as1n06x5 input19 (.a(tl_i[26]),
    .o(net19));
 b15bfn001as1n06x5 input20 (.a(tl_i[27]),
    .o(net20));
 b15bfn001as1n06x5 input21 (.a(tl_i[28]),
    .o(net21));
 b15bfn001as1n06x5 input22 (.a(tl_i[29]),
    .o(net22));
 b15bfn001as1n06x5 input23 (.a(tl_i[30]),
    .o(net23));
 b15bfn001as1n06x5 input24 (.a(tl_i[31]),
    .o(net24));
 b15bfn001as1n08x5 input25 (.a(tl_i[32]),
    .o(net25));
 b15bfn001as1n08x5 input26 (.a(tl_i[33]),
    .o(net26));
 b15bfn001as1n08x5 input27 (.a(tl_i[34]),
    .o(net27));
 b15bfn001as1n08x5 input28 (.a(tl_i[35]),
    .o(net28));
 b15bfn001ah1n08x5 input29 (.a(tl_i[36]),
    .o(net29));
 b15bfn001as1n08x5 input30 (.a(tl_i[37]),
    .o(net30));
 b15bfn001as1n08x5 input31 (.a(tl_i[38]),
    .o(net31));
 b15bfn001ah1n12x5 input32 (.a(tl_i[39]),
    .o(net32));
 b15bfn001as1n06x5 input33 (.a(tl_i[40]),
    .o(net33));
 b15bfn001ah1n08x5 input34 (.a(tl_i[41]),
    .o(net34));
 b15bfn001ah1n08x5 input35 (.a(tl_i[42]),
    .o(net35));
 b15bfn001ah1n08x5 input36 (.a(tl_i[43]),
    .o(net36));
 b15bfn001as1n08x5 input37 (.a(tl_i[44]),
    .o(net37));
 b15bfn001ah1n08x5 input38 (.a(tl_i[45]),
    .o(net38));
 b15bfn001ah1n08x5 input39 (.a(tl_i[46]),
    .o(net39));
 b15bfn001as1n06x5 input40 (.a(tl_i[47]),
    .o(net40));
 b15bfn000as1n02x5 input41 (.a(tl_i[48]),
    .o(net41));
 b15bfn000ah1n04x5 input42 (.a(tl_i[49]),
    .o(net42));
 b15bfn000as1n02x5 input43 (.a(tl_i[50]),
    .o(net43));
 b15bfn000ah1n03x5 input44 (.a(tl_i[51]),
    .o(net44));
 b15bfn000as1n02x5 input45 (.a(tl_i[52]),
    .o(net45));
 b15bfn000as1n02x5 input46 (.a(tl_i[53]),
    .o(net46));
 b15bfn000as1n02x5 input47 (.a(tl_i[54]),
    .o(net47));
 b15bfn000as1n02x5 input48 (.a(tl_i[55]),
    .o(net48));
 b15bfn001ah1n48x5 input49 (.a(tl_i[56]),
    .o(net49));
 b15bfn001ah1n48x5 input50 (.a(tl_i[57]),
    .o(net50));
 b15bfn000ah1n48x5 input51 (.a(tl_i[58]),
    .o(net51));
 b15bfn001ah1n48x5 input52 (.a(tl_i[59]),
    .o(net52));
 b15bfn001ah1n24x5 input53 (.a(tl_i[60]),
    .o(net53));
 b15bfn001ah1n24x5 input54 (.a(tl_i[61]),
    .o(net54));
 b15bfn001ah1n16x5 input55 (.a(tl_i[62]),
    .o(net55));
 b15bfn000as1n04x5 input56 (.a(tl_i[63]),
    .o(net56));
 b15bfn000ah1n03x5 input57 (.a(tl_i[64]),
    .o(net57));
 b15bfn001as1n12x5 input58 (.a(tl_i[65]),
    .o(net58));
 b15bfn001as1n16x5 input59 (.a(tl_i[66]),
    .o(net59));
 b15bfn001aq1n06x5 input60 (.a(tl_i[67]),
    .o(net60));
 b15bfn001as1n06x5 input61 (.a(tl_i[68]),
    .o(net61));
 b15bfn001aq1n06x5 input62 (.a(tl_i[69]),
    .o(net62));
 b15bfn001aq1n06x5 input63 (.a(tl_i[70]),
    .o(net63));
 b15bfn000as1n04x5 input64 (.a(tl_i[71]),
    .o(net64));
 b15bfn000ah1n03x5 input65 (.a(tl_i[72]),
    .o(net65));
 b15bfn001as1n12x5 input66 (.a(tl_i[92]),
    .o(net66));
 b15bfn001as1n12x5 input67 (.a(tl_i[93]),
    .o(net67));
 b15bfn001as1n12x5 input68 (.a(tl_i[94]),
    .o(net68));
 b15bfn001ah1n12x5 input69 (.a(tl_i[95]),
    .o(net69));
 b15bfn001as1n12x5 input70 (.a(tl_i[96]),
    .o(net70));
 b15bfn001as1n12x5 input71 (.a(tl_i[97]),
    .o(net71));
 b15bfn000as1n12x5 input72 (.a(tl_i[98]),
    .o(net72));
 b15bfn001ah1n12x5 input73 (.a(tl_i[99]),
    .o(net73));
 b15bfn000ah1n03x5 output74 (.a(net352),
    .o(net353));
 b15bfn000ah1n03x5 output75 (.a(net495),
    .o(tl_o[16]));
 b15bfn000ah1n03x5 output76 (.a(net445),
    .o(tl_o[17]));
 b15bfn000ah1n03x5 output77 (.a(net519),
    .o(tl_o[18]));
 b15bfn000ah1n03x5 output78 (.a(net460),
    .o(tl_o[19]));
 b15bfn000ah1n03x5 output79 (.a(net360),
    .o(net361));
 b15bfn000ah1n03x5 output80 (.a(net432),
    .o(net433));
 b15bfn000ah1n03x5 output81 (.a(net479),
    .o(tl_o[21]));
 b15bfn000ah1n03x5 output82 (.a(net464),
    .o(tl_o[22]));
 b15bfn000ah1n03x5 output83 (.a(net415),
    .o(net416));
 b15bfn000ah1n03x5 output84 (.a(net449),
    .o(tl_o[24]));
 b15bfn000ah1n03x5 output85 (.a(net476),
    .o(tl_o[25]));
 b15bfn000ah1n03x5 output86 (.a(net542),
    .o(tl_o[26]));
 b15bfn000ah1n03x5 output87 (.a(net441),
    .o(tl_o[27]));
 b15bfn000ah1n03x5 output88 (.a(net436),
    .o(tl_o[28]));
 b15bfn000ah1n03x5 output89 (.a(net427),
    .o(net428));
 b15bfn000ah1n03x5 output90 (.a(net404),
    .o(tl_o[2]));
 b15bfn000ah1n03x5 output91 (.a(net456),
    .o(tl_o[30]));
 b15bfn000ah1n03x5 output92 (.a(net482),
    .o(tl_o[31]));
 b15bfn000ah1n03x5 output93 (.a(net471),
    .o(net472));
 b15bfn000ah1n03x5 output94 (.a(net508),
    .o(tl_o[33]));
 b15bfn000ah1n03x5 output95 (.a(net511),
    .o(net512));
 b15bfn000ah1n03x5 output96 (.a(net467),
    .o(net468));
 b15bfn000ah1n03x5 output97 (.a(net498),
    .o(net499));
 b15bfn000ah1n03x5 output98 (.a(net452),
    .o(net453));
 b15bfn000ah1n03x5 output99 (.a(net515),
    .o(tl_o[38]));
 b15bfn000ah1n03x5 output100 (.a(net423),
    .o(net424));
 b15bfn000ah1n03x5 output101 (.a(net367),
    .o(net368));
 b15bfn000ah1n03x5 output102 (.a(net539),
    .o(tl_o[40]));
 b15bfn000ah1n03x5 output103 (.a(net528),
    .o(tl_o[41]));
 b15bfn000ah1n03x5 output104 (.a(net419),
    .o(net420));
 b15bfn000ah1n03x5 output105 (.a(net548),
    .o(tl_o[43]));
 b15bfn000ah1n03x5 output106 (.a(net536),
    .o(tl_o[44]));
 b15bfn000ah1n03x5 output107 (.a(net505),
    .o(tl_o[45]));
 b15bfn000ah1n03x5 output108 (.a(net545),
    .o(tl_o[46]));
 b15bfn000ah1n03x5 output109 (.a(net491),
    .o(tl_o[47]));
 b15bfn000ah1n03x5 output110 (.a(net401),
    .o(net402));
 b15bfn000ah1n03x5 output111 (.a(net392),
    .o(tl_o[4]));
 b15bfn000ah1n03x5 output112 (.a(net409),
    .o(net410));
 b15bfn000ah1n03x5 output113 (.a(net487),
    .o(net488));
 b15bfn000ah1n03x5 output114 (.a(net521),
    .o(net522));
 b15bfn000ah1n03x5 output115 (.a(net398),
    .o(net399));
 b15bfn000ah1n03x5 output116 (.a(net406),
    .o(net407));
 b15bfn000ah1n03x5 output117 (.a(net484),
    .o(net485));
 b15bfn000ah1n03x5 output118 (.a(net524),
    .o(net525));
 b15bfn000ah1n03x5 output119 (.a(net501),
    .o(net502));
 b15bfn000ah1n03x5 output120 (.a(net530),
    .o(net531));
 b15bfn000ah1n03x5 output121 (.a(net375),
    .o(net376));
 b15bfn000ah1n03x5 output122 (.a(net381),
    .o(net382));
 b15bfn000ah1n03x5 output123 (.a(net395),
    .o(net396));
 b15bfn000ah1n03x5 output124 (.a(net387),
    .o(net388));
 b15bfn000ah1n03x5 output125 (.a(net378),
    .o(tl_o[7]));
 b15bfn000ah1n03x5 output126 (.a(net390),
    .o(tl_o[8]));
 b15bfn001as1n24x5 fanout127 (.a(net129),
    .o(net127));
 b15bfn001as1n12x5 fanout128 (.a(net431),
    .o(net128));
 b15bfn001ah1n32x5 wire129 (.a(net128),
    .o(net129));
 b15bfn001as1n24x5 fanout130 (.a(net430),
    .o(net130));
 b15bfn001ah1n48x5 fanout131 (.a(net132),
    .o(net131));
 b15bfn001as1n80x5 fanout132 (.a(n383),
    .o(net132));
 b15bfn001as1n48x5 fanout133 (.a(net135),
    .o(net133));
 b15bfn001ah1n80x5 fanout134 (.a(n381),
    .o(net134));
 b15bfn000as1n32x5 wire135 (.a(net134),
    .o(net135));
 b15bfn001as1n16x5 max_length136 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_N9),
    .o(net136));
 b15bfn001ah1n24x5 wire137 (.a(u_tlul_adapter_sram_rdata_tlword[12]),
    .o(net137));
 b15bfn001ah1n24x5 wire138 (.a(u_tlul_adapter_sram_rdata_tlword[10]),
    .o(net138));
 b15bfn001ah1n24x5 wire139 (.a(u_tlul_adapter_sram_rdata_tlword[4]),
    .o(net139));
 b15bfn001ah1n32x5 wire140 (.a(u_tlul_adapter_sram_rdata_tlword[2]),
    .o(net140));
 b15bfn001ah1n32x5 wire141 (.a(u_tlul_adapter_sram_rdata_tlword[0]),
    .o(net141));
 b15bfn001ah1n48x5 wire142 (.a(n434),
    .o(net142));
 b15bfn001as1n48x5 wire143 (.a(net533),
    .o(net143));
 b15bfn001as1n32x5 wire144 (.a(net145),
    .o(net144));
 b15bfn001ah1n24x5 wire145 (.a(n_0_net_),
    .o(net145));
 b15bfn001ah1n16x5 wire146 (.a(net442),
    .o(net146));
 b15bfn000ah1n24x5 wire147 (.a(net492),
    .o(net147));
 b15bfn001as1n16x5 wire148 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[19]),
    .o(net148));
 b15bfn001as1n16x5 wire149 (.a(net473),
    .o(net149));
 b15bfn000ah1n24x5 wire150 (.a(net446),
    .o(net150));
 b15bfn001as1n16x5 wire151 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[15]),
    .o(net151));
 b15bfn001as1n16x5 wire152 (.a(net461),
    .o(net152));
 b15bfn001ah1n16x5 wire153 (.a(net457),
    .o(net153));
 b15bfn000ah1n24x5 wire154 (.a(net516),
    .o(net154));
 b15bfn001as1n24x5 wire155 (.a(net156),
    .o(net155));
 b15bfn001as1n12x5 wire156 (.a(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[0]),
    .o(net156));
 b15bfn000as1n32x5 wire157 (.a(net158),
    .o(net157));
 b15bfn001ah1n24x5 wire158 (.a(wen),
    .o(net158));
 b15bfn001as1n24x5 wire159 (.a(net551),
    .o(net159));
 b15bfn001ah1n16x5 wire160 (.a(net550),
    .o(net160));
 b15bfn001as1n12x5 max_cap161 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_fifo_rptr_1_),
    .o(net161));
 b15bfn001ah1n12x5 load_slew162 (.a(net163),
    .o(net162));
 b15bfn001as1n12x5 wire163 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_wptr_value_0_),
    .o(net163));
 b15bfn000ah1n24x5 wire164 (.a(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_rptr_value_0_),
    .o(net164));
 b15bfn000as1n24x5 wire165 (.a(net394),
    .o(net165));
 b15bfn001as1n08x5 wire166 (.a(net393),
    .o(net166));
 b15bfn001ah1n16x5 wire167 (.a(net383),
    .o(net167));
 b15bfn001ah1n16x5 wire168 (.a(net354),
    .o(net168));
 b15bfn001ah1n16x5 wire169 (.a(net348),
    .o(net169));
 b15bfn001as1n16x5 wire170 (.a(net362),
    .o(net170));
 b15bfn001ah1n32x5 wire171 (.a(net172),
    .o(net171));
 b15bfn001ah1n64x5 wire172 (.a(n328),
    .o(net172));
 b15bfn001ah1n24x5 wire173 (.a(net7),
    .o(net173));
 b15bfn001ah1n24x5 wire174 (.a(net58),
    .o(net174));
 b15bfn000ah1n48x5 wire175 (.a(net50),
    .o(net175));
 b15bfn001as1n32x5 wire176 (.a(net5),
    .o(net176));
 b15bfn001as1n32x5 wire177 (.a(net49),
    .o(net177));
 b15bfn001ah1n24x5 wire178 (.a(net15),
    .o(net178));
 b15bfn001ah1n24x5 wire179 (.a(rdata[15]),
    .o(net179));
 b15tilo00an1n03x5 rvalid_reg_u_tlul_adapter_sram_intg_error_q_reg_180 (.o(net180));
 b15tilo00an1n03x5 rvalid_reg_u_tlul_adapter_sram_intg_error_q_reg_181 (.o(net181));
 b15tilo00an1n03x5 u_sram_182 (.o(net182));
 b15tilo00an1n03x5 u_sram_183 (.o(net183));
 b15tilo00an1n03x5 u_sram_184 (.o(net184));
 b15tilo00an1n03x5 u_sram_185 (.o(net185));
 b15tilo00an1n03x5 u_sram_186 (.o(net186));
 b15tilo00an1n03x5 u_sram_187 (.o(net187));
 b15tilo00an1n03x5 u_sram_188 (.o(net188));
 b15tilo00an1n03x5 u_sram_189 (.o(net189));
 b15tilo00an1n03x5 u_sram_190 (.o(net190));
 b15tilo00an1n03x5 u_sram_191 (.o(net191));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_clk_gate_gen_normal_fifo_storage_reg_0__0_latch_192 (.o(net192));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_clk_gate_gen_normal_fifo_storage_reg_0__latch_193 (.o(net193));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__1__194 (.o(net194));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__1__195 (.o(net195));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__11__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__12__196 (.o(net196));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__11__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__12__197 (.o(net197));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__13__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__14__198 (.o(net198));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__13__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__14__199 (.o(net199));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__15__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__16__200 (.o(net200));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__15__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__16__201 (.o(net201));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__15__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__16__202 (.o(net202));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__3__203 (.o(net203));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__3__204 (.o(net204));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__5__205 (.o(net205));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__5__206 (.o(net206));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__7__207 (.o(net207));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__7__208 (.o(net208));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__8__209 (.o(net209));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__9__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__10__210 (.o(net210));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__9__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__10__211 (.o(net211));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__212 (.o(net212));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__213 (.o(net213));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__214 (.o(net214));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__215 (.o(net215));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst_reg_216 (.o(net216));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst_reg_217 (.o(net217));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_clk_gate_gen_normal_fifo_storage_reg_0__0_latch_218 (.o(net218));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_clk_gate_gen_normal_fifo_storage_reg_0__latch_219 (.o(net219));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1__220 (.o(net220));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1__221 (.o(net221));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1__222 (.o(net222));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1__223 (.o(net223));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__10__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__11__224 (.o(net224));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__10__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__11__225 (.o(net225));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__12__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__13__226 (.o(net226));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__12__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__13__227 (.o(net227));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__14__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__15__228 (.o(net228));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__14__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__15__229 (.o(net229));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__16__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__17__230 (.o(net230));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__16__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__17__231 (.o(net231));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__18__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__19__232 (.o(net232));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__18__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__19__233 (.o(net233));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__20__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__21__234 (.o(net234));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__20__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__21__235 (.o(net235));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__22__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__23__236 (.o(net236));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__22__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__23__237 (.o(net237));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__24__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__25__238 (.o(net238));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__24__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__25__239 (.o(net239));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__26__240 (.o(net240));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__27__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__28__241 (.o(net241));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__27__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__28__242 (.o(net242));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__29__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__30__243 (.o(net243));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__29__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__30__244 (.o(net244));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3__245 (.o(net245));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3__246 (.o(net246));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3__247 (.o(net247));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3__248 (.o(net248));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__31__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__32__249 (.o(net249));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__31__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__32__250 (.o(net250));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__33__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__34__251 (.o(net251));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__33__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__34__252 (.o(net252));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__35__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__36__253 (.o(net253));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__35__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__36__254 (.o(net254));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__37__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__38__255 (.o(net255));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__37__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__38__256 (.o(net256));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__39__257 (.o(net257));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5__258 (.o(net258));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5__259 (.o(net259));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5__260 (.o(net260));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5__261 (.o(net261));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7__262 (.o(net262));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7__263 (.o(net263));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7__264 (.o(net264));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7__265 (.o(net265));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__8__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__9__266 (.o(net266));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__8__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__9__267 (.o(net267));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__268 (.o(net268));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__269 (.o(net269));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__270 (.o(net270));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__271 (.o(net271));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst_reg_272 (.o(net272));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst_reg_273 (.o(net273));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__0__274 (.o(net274));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__1__275 (.o(net275));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__2__276 (.o(net276));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__3__277 (.o(net277));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__4__278 (.o(net278));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__279 (.o(net279));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__280 (.o(net280));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__281 (.o(net281));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__282 (.o(net282));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst_reg_283 (.o(net283));
 b15tilo00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst_reg_284 (.o(net284));
 b15tihi00an1n03x5 U588_286 (.o(net286));
 b15tihi00an1n03x5 U594_287 (.o(net287));
 b15tihi00an1n03x5 U602_288 (.o(net288));
 b15tihi00an1n03x5 U622_289 (.o(net289));
 b15tihi00an1n03x5 U637_290 (.o(net290));
 b15tihi00an1n03x5 U702_291 (.o(net291));
 b15tihi00an1n03x5 U704_292 (.o(net292));
 b15tihi00an1n03x5 U706_293 (.o(net293));
 b15tihi00an1n03x5 U708_294 (.o(net294));
 b15tihi00an1n03x5 U710_295 (.o(net295));
 b15tihi00an1n03x5 U712_296 (.o(net296));
 b15tihi00an1n03x5 U714_297 (.o(net297));
 b15tihi00an1n03x5 rvalid_reg_u_tlul_adapter_sram_intg_error_q_reg_298 (.o(net298));
 b15tihi00an1n03x5 u_sram_299 (.o(net299));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__1__300 (.o(net300));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__11__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__12__301 (.o(net301));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__13__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__14__302 (.o(net302));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__15__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__16__303 (.o(net303));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__3__304 (.o(net304));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__5__305 (.o(net305));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__7__306 (.o(net306));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__8__307 (.o(net307));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__9__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_reg_0__10__308 (.o(net308));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__309 (.o(net309));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__310 (.o(net310));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__311 (.o(net311));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_under_rst_reg_312 (.o(net312));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__1__313 (.o(net313));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__10__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__11__314 (.o(net314));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__12__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__13__315 (.o(net315));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__14__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__15__316 (.o(net316));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__16__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__17__317 (.o(net317));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__18__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__19__318 (.o(net318));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__20__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__21__319 (.o(net319));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__22__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__23__320 (.o(net320));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__24__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__25__321 (.o(net321));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__26__322 (.o(net322));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__27__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__28__323 (.o(net323));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__29__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__30__324 (.o(net324));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__2__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__3__325 (.o(net325));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__31__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__32__326 (.o(net326));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__33__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__34__327 (.o(net327));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__35__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__36__328 (.o(net328));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__37__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__38__329 (.o(net329));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__39__330 (.o(net330));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__4__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__5__331 (.o(net331));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__6__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__7__332 (.o(net332));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__8__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_reg_0__9__333 (.o(net333));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__334 (.o(net334));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__335 (.o(net335));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__336 (.o(net336));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst_reg_337 (.o(net337));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__0__338 (.o(net338));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__1__339 (.o(net339));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__2__340 (.o(net340));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__3__341 (.o(net341));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_reg_0__4__342 (.o(net342));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_0__u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_0__343 (.o(net343));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_rptr_o_reg_1__344 (.o(net344));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_u_fifo_cnt_wptr_o_reg_1__345 (.o(net345));
 b15tihi00an1n03x5 u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst_reg_346 (.o(net346));
 b15cbf000an1n16x5 clkbuf_1_0__f_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_1_0__leaf_clk_i));
 b15cbf000an1n16x5 clkbuf_1_1__f_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_1_1__leaf_clk_i));
 b15cbf000an1n16x5 clkbuf_0_u_tlul_adapter_sram_u_rspfifo_net616 (.clk(u_tlul_adapter_sram_u_rspfifo_net616),
    .clkout(clknet_0_u_tlul_adapter_sram_u_rspfifo_net616));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_tlul_adapter_sram_u_rspfifo_net616 (.clk(clknet_0_u_tlul_adapter_sram_u_rspfifo_net616),
    .clkout(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net616));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_tlul_adapter_sram_u_rspfifo_net616 (.clk(clknet_0_u_tlul_adapter_sram_u_rspfifo_net616),
    .clkout(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net616));
 b15cbf000an1n16x5 clkbuf_0_u_tlul_adapter_sram_u_rspfifo_net622 (.clk(u_tlul_adapter_sram_u_rspfifo_net622),
    .clkout(clknet_0_u_tlul_adapter_sram_u_rspfifo_net622));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_tlul_adapter_sram_u_rspfifo_net622 (.clk(clknet_0_u_tlul_adapter_sram_u_rspfifo_net622),
    .clkout(clknet_1_0__leaf_u_tlul_adapter_sram_u_rspfifo_net622));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_tlul_adapter_sram_u_rspfifo_net622 (.clk(clknet_0_u_tlul_adapter_sram_u_rspfifo_net622),
    .clkout(clknet_1_1__leaf_u_tlul_adapter_sram_u_rspfifo_net622));
 b15cbf000an1n16x5 clkbuf_0_u_tlul_adapter_sram_u_reqfifo_net644 (.clk(u_tlul_adapter_sram_u_reqfifo_net644),
    .clkout(clknet_0_u_tlul_adapter_sram_u_reqfifo_net644));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_tlul_adapter_sram_u_reqfifo_net644 (.clk(clknet_0_u_tlul_adapter_sram_u_reqfifo_net644),
    .clkout(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net644));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_tlul_adapter_sram_u_reqfifo_net644 (.clk(clknet_0_u_tlul_adapter_sram_u_reqfifo_net644),
    .clkout(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net644));
 b15cbf000an1n16x5 clkbuf_0_u_tlul_adapter_sram_u_reqfifo_net650 (.clk(u_tlul_adapter_sram_u_reqfifo_net650),
    .clkout(clknet_0_u_tlul_adapter_sram_u_reqfifo_net650));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_tlul_adapter_sram_u_reqfifo_net650 (.clk(clknet_0_u_tlul_adapter_sram_u_reqfifo_net650),
    .clkout(clknet_1_0__leaf_u_tlul_adapter_sram_u_reqfifo_net650));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_tlul_adapter_sram_u_reqfifo_net650 (.clk(clknet_0_u_tlul_adapter_sram_u_reqfifo_net650),
    .clkout(clknet_1_1__leaf_u_tlul_adapter_sram_u_reqfifo_net650));
 b15bfn001as1n16x5 wire1 (.a(clk_i),
    .o(net347));
 b15cbf034ar1n64x5 hold2 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_wptr_value_0_),
    .clkout(net348));
 b15cbf034ar1n64x5 hold3 (.clk(net169),
    .clkout(net349));
 b15cbf034ar1n64x5 hold4 (.clk(n358),
    .clkout(net350));
 b15cbf034ar1n64x5 hold5 (.clk(n361),
    .clkout(net351));
 b15cbf034ar1n64x5 hold6 (.clk(net74),
    .clkout(net352));
 b15cbf034ar1n64x5 hold7 (.clk(net353),
    .clkout(tl_o[0]));
 b15cbf034ar1n64x5 hold8 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_wptr_value_0_),
    .clkout(net354));
 b15cbf034ar1n64x5 hold9 (.clk(net168),
    .clkout(net355));
 b15cbf034ar1n64x5 hold10 (.clk(n368),
    .clkout(net356));
 b15cbf034ar1n64x5 hold11 (.clk(net386),
    .clkout(net357));
 b15cbf034ar1n64x5 hold12 (.clk(n386),
    .clkout(net358));
 b15cbf034ar1n64x5 hold13 (.clk(n378),
    .clkout(net359));
 b15cbf034ar1n64x5 hold14 (.clk(net79),
    .clkout(net360));
 b15cbf034ar1n64x5 hold15 (.clk(net361),
    .clkout(tl_o[1]));
 b15cbf034ar1n64x5 hold16 (.clk(rvalid),
    .clkout(net362));
 b15cbf034ar1n64x5 hold17 (.clk(net170),
    .clkout(net363));
 b15cbf034ar1n64x5 hold18 (.clk(n369),
    .clkout(net364));
 b15cbf034ar1n64x5 hold19 (.clk(n375),
    .clkout(net365));
 b15cbf034ar1n64x5 hold20 (.clk(net373),
    .clkout(net366));
 b15cbf034ar1n64x5 hold21 (.clk(net101),
    .clkout(net367));
 b15cbf034ar1n64x5 hold22 (.clk(net368),
    .clkout(tl_o[3]));
 b15cbf034ar1n64x5 hold23 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_fifo_wptr_1_),
    .clkout(net369));
 b15cbf034ar1n64x5 hold24 (.clk(n357),
    .clkout(net370));
 b15cbf034ar1n64x5 hold25 (.clk(n384),
    .clkout(net371));
 b15cbf034ar1n64x5 hold26 (.clk(n374),
    .clkout(net372));
 b15cbf034ar1n64x5 hold27 (.clk(n385),
    .clkout(net373));
 b15cbf034ar1n64x5 hold28 (.clk(net366),
    .clkout(net374));
 b15cbf034ar1n64x5 hold29 (.clk(net121),
    .clkout(net375));
 b15cbf034ar1n64x5 hold30 (.clk(net376),
    .clkout(tl_o[5]));
 b15cbf034ar1n64x5 hold31 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[6]),
    .clkout(net377));
 b15cbf034ar1n64x5 hold32 (.clk(net125),
    .clkout(net378));
 b15cbf034ar1n64x5 hold33 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[15]),
    .clkout(net379));
 b15cbf034ar1n64x5 hold34 (.clk(n379),
    .clkout(net380));
 b15cbf034ar1n64x5 hold35 (.clk(net122),
    .clkout(net381));
 b15cbf034ar1n64x5 hold36 (.clk(net382),
    .clkout(tl_o[62]));
 b15cbf034ar1n64x5 hold37 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_fifo_wptr_1_),
    .clkout(net383));
 b15cbf034ar1n64x5 hold38 (.clk(net167),
    .clkout(net384));
 b15cbf034ar1n64x5 hold39 (.clk(n367),
    .clkout(net385));
 b15cbf034ar1n64x5 hold40 (.clk(n380),
    .clkout(net386));
 b15cbf034ar1n64x5 hold41 (.clk(net124),
    .clkout(net387));
 b15cbf034ar1n64x5 hold42 (.clk(net388),
    .clkout(tl_o[6]));
 b15cbf034ar1n64x5 hold43 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[7]),
    .clkout(net389));
 b15cbf034ar1n64x5 hold44 (.clk(net126),
    .clkout(net390));
 b15cbf034ar1n64x5 hold45 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[3]),
    .clkout(net391));
 b15cbf034ar1n64x5 hold46 (.clk(net111),
    .clkout(net392));
 b15cbf034ar1n64x5 hold47 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_under_rst),
    .clkout(net393));
 b15cbf034ar1n64x5 hold48 (.clk(net166),
    .clkout(net394));
 b15cbf034ar1n64x5 hold49 (.clk(net123),
    .clkout(net395));
 b15cbf034ar1n64x5 hold50 (.clk(net396),
    .clkout(tl_o[65]));
 b15cbf034ar1n64x5 hold51 (.clk(net553),
    .clkout(net397));
 b15cbf034ar1n64x5 hold52 (.clk(net115),
    .clkout(net398));
 b15cbf034ar1n64x5 hold53 (.clk(net399),
    .clkout(tl_o[53]));
 b15cbf034ar1n64x5 hold54 (.clk(net554),
    .clkout(net400));
 b15cbf034ar1n64x5 hold55 (.clk(net110),
    .clkout(net401));
 b15cbf034ar1n64x5 hold56 (.clk(net402),
    .clkout(tl_o[49]));
 b15cbf034ar1n64x5 hold57 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[1]),
    .clkout(net403));
 b15cbf034ar1n64x5 hold58 (.clk(net90),
    .clkout(net404));
 b15cbf034ar1n64x5 hold59 (.clk(net555),
    .clkout(net405));
 b15cbf034ar1n64x5 hold60 (.clk(net116),
    .clkout(net406));
 b15cbf034ar1n64x5 hold61 (.clk(net407),
    .clkout(tl_o[54]));
 b15cbf034ar1n64x5 hold62 (.clk(net556),
    .clkout(net408));
 b15cbf034ar1n64x5 hold63 (.clk(net112),
    .clkout(net409));
 b15cbf034ar1n64x5 hold64 (.clk(net410),
    .clkout(tl_o[50]));
 b15cbf034ar1n64x5 hold65 (.clk(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[1]),
    .clkout(net411));
 b15cbf034ar1n64x5 hold66 (.clk(n416),
    .clkout(net412));
 b15cbf034ar1n64x5 hold67 (.clk(u_tlul_adapter_sram_rdata_tlword[7]),
    .clkout(net413));
 b15cbf034ar1n64x5 hold68 (.clk(n417),
    .clkout(net414));
 b15cbf034ar1n64x5 hold69 (.clk(net83),
    .clkout(net415));
 b15cbf034ar1n64x5 hold70 (.clk(net416),
    .clkout(tl_o[23]));
 b15cbf034ar1n64x5 hold71 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[34]),
    .clkout(net417));
 b15cbf034ar1n64x5 hold72 (.clk(n390),
    .clkout(net418));
 b15cbf034ar1n64x5 hold73 (.clk(net104),
    .clkout(net419));
 b15cbf034ar1n64x5 hold74 (.clk(net420),
    .clkout(tl_o[42]));
 b15cbf034ar1n64x5 hold75 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[31]),
    .clkout(net421));
 b15cbf034ar1n64x5 hold76 (.clk(n405),
    .clkout(net422));
 b15cbf034ar1n64x5 hold77 (.clk(net100),
    .clkout(net423));
 b15cbf034ar1n64x5 hold78 (.clk(net424),
    .clkout(tl_o[39]));
 b15cbf034ar1n64x5 hold79 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[21]),
    .clkout(net425));
 b15cbf034ar1n64x5 hold80 (.clk(n427),
    .clkout(net426));
 b15cbf034ar1n64x5 hold81 (.clk(net89),
    .clkout(net427));
 b15cbf034ar1n64x5 hold82 (.clk(net428),
    .clkout(tl_o[29]));
 b15cbf034ar1n64x5 hold83 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[13]),
    .clkout(net429));
 b15cbf034ar1n64x5 hold84 (.clk(n389),
    .clkout(net430));
 b15cbf034ar1n64x5 hold85 (.clk(net130),
    .clkout(net431));
 b15cbf034ar1n64x5 hold86 (.clk(net80),
    .clkout(net432));
 b15cbf034ar1n64x5 hold87 (.clk(net433),
    .clkout(tl_o[20]));
 b15cbf034ar1n64x5 hold88 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[20]),
    .clkout(net434));
 b15cbf034ar1n64x5 hold89 (.clk(n426),
    .clkout(net435));
 b15cbf034ar1n64x5 hold90 (.clk(net88),
    .clkout(net436));
 b15cbf034ar1n64x5 hold91 (.clk(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[2]),
    .clkout(net437));
 b15cbf034ar1n64x5 hold92 (.clk(n429),
    .clkout(net438));
 b15cbf034ar1n64x5 hold93 (.clk(u_tlul_adapter_sram_rdata_tlword[11]),
    .clkout(net439));
 b15cbf034ar1n64x5 hold94 (.clk(n424),
    .clkout(net440));
 b15cbf034ar1n64x5 hold95 (.clk(net87),
    .clkout(net441));
 b15cbf034ar1n64x5 hold96 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[9]),
    .clkout(net442));
 b15cbf034ar1n64x5 hold97 (.clk(net146),
    .clkout(net443));
 b15cbf034ar1n64x5 hold98 (.clk(n410),
    .clkout(net444));
 b15cbf034ar1n64x5 hold99 (.clk(net76),
    .clkout(net445));
 b15cbf034ar1n64x5 hold100 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[16]),
    .clkout(net446));
 b15cbf034ar1n64x5 hold101 (.clk(net150),
    .clkout(net447));
 b15cbf034ar1n64x5 hold102 (.clk(n419),
    .clkout(net448));
 b15cbf034ar1n64x5 hold103 (.clk(net84),
    .clkout(net449));
 b15cbf034ar1n64x5 hold104 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[29]),
    .clkout(net450));
 b15cbf034ar1n64x5 hold105 (.clk(n403),
    .clkout(net451));
 b15cbf034ar1n64x5 hold106 (.clk(net98),
    .clkout(net452));
 b15cbf034ar1n64x5 hold107 (.clk(net453),
    .clkout(tl_o[37]));
 b15cbf034ar1n64x5 hold108 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[22]),
    .clkout(net454));
 b15cbf034ar1n64x5 hold109 (.clk(n428),
    .clkout(net455));
 b15cbf034ar1n64x5 hold110 (.clk(net91),
    .clkout(net456));
 b15cbf034ar1n64x5 hold111 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[11]),
    .clkout(net457));
 b15cbf034ar1n64x5 hold112 (.clk(net153),
    .clkout(net458));
 b15cbf034ar1n64x5 hold113 (.clk(n412),
    .clkout(net459));
 b15cbf034ar1n64x5 hold114 (.clk(net78),
    .clkout(net460));
 b15cbf034ar1n64x5 hold115 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[14]),
    .clkout(net461));
 b15cbf034ar1n64x5 hold116 (.clk(net152),
    .clkout(net462));
 b15cbf034ar1n64x5 hold117 (.clk(n415),
    .clkout(net463));
 b15cbf034ar1n64x5 hold118 (.clk(net82),
    .clkout(net464));
 b15cbf034ar1n64x5 hold119 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[27]),
    .clkout(net465));
 b15cbf034ar1n64x5 hold120 (.clk(n438),
    .clkout(net466));
 b15cbf034ar1n64x5 hold121 (.clk(net96),
    .clkout(net467));
 b15cbf034ar1n64x5 hold122 (.clk(net468),
    .clkout(tl_o[35]));
 b15cbf034ar1n64x5 hold123 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[24]),
    .clkout(net469));
 b15cbf034ar1n64x5 hold124 (.clk(n431),
    .clkout(net470));
 b15cbf034ar1n64x5 hold125 (.clk(net93),
    .clkout(net471));
 b15cbf034ar1n64x5 hold126 (.clk(net472),
    .clkout(tl_o[32]));
 b15cbf034ar1n64x5 hold127 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[17]),
    .clkout(net473));
 b15cbf034ar1n64x5 hold128 (.clk(net149),
    .clkout(net474));
 b15cbf034ar1n64x5 hold129 (.clk(n420),
    .clkout(net475));
 b15cbf034ar1n64x5 hold130 (.clk(net85),
    .clkout(net476));
 b15cbf034ar1n64x5 hold131 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[13]),
    .clkout(net477));
 b15cbf034ar1n64x5 hold132 (.clk(n414),
    .clkout(net478));
 b15cbf034ar1n64x5 hold133 (.clk(net81),
    .clkout(net479));
 b15cbf034ar1n64x5 hold134 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[23]),
    .clkout(net480));
 b15cbf034ar1n64x5 hold135 (.clk(n430),
    .clkout(net481));
 b15cbf034ar1n64x5 hold136 (.clk(net92),
    .clkout(net482));
 b15cbf034ar1n64x5 hold137 (.clk(net557),
    .clkout(net483));
 b15cbf034ar1n64x5 hold138 (.clk(net117),
    .clkout(net484));
 b15cbf034ar1n64x5 hold139 (.clk(net485),
    .clkout(tl_o[55]));
 b15cbf034ar1n64x5 hold140 (.clk(net558),
    .clkout(net486));
 b15cbf034ar1n64x5 hold141 (.clk(net113),
    .clkout(net487));
 b15cbf034ar1n64x5 hold142 (.clk(net488),
    .clkout(tl_o[51]));
 b15cbf034ar1n64x5 hold143 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[39]),
    .clkout(net489));
 b15cbf034ar1n64x5 hold144 (.clk(n395),
    .clkout(net490));
 b15cbf034ar1n64x5 hold145 (.clk(net109),
    .clkout(net491));
 b15cbf034ar1n64x5 hold146 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[8]),
    .clkout(net492));
 b15cbf034ar1n64x5 hold147 (.clk(net147),
    .clkout(net493));
 b15cbf034ar1n64x5 hold148 (.clk(n409),
    .clkout(net494));
 b15cbf034ar1n64x5 hold149 (.clk(net75),
    .clkout(net495));
 b15cbf034ar1n64x5 hold150 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[28]),
    .clkout(net496));
 b15cbf034ar1n64x5 hold151 (.clk(n402),
    .clkout(net497));
 b15cbf034ar1n64x5 hold152 (.clk(net97),
    .clkout(net498));
 b15cbf034ar1n64x5 hold153 (.clk(net499),
    .clkout(tl_o[36]));
 b15cbf034ar1n64x5 hold154 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[8]),
    .clkout(net500));
 b15cbf034ar1n64x5 hold155 (.clk(net119),
    .clkout(net501));
 b15cbf034ar1n64x5 hold156 (.clk(net502),
    .clkout(tl_o[57]));
 b15cbf034ar1n64x5 hold157 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[37]),
    .clkout(net503));
 b15cbf034ar1n64x5 hold158 (.clk(n401),
    .clkout(net504));
 b15cbf034ar1n64x5 hold159 (.clk(net107),
    .clkout(net505));
 b15cbf034ar1n64x5 hold160 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[25]),
    .clkout(net506));
 b15cbf034ar1n64x5 hold161 (.clk(n432),
    .clkout(net507));
 b15cbf034ar1n64x5 hold162 (.clk(net94),
    .clkout(net508));
 b15cbf034ar1n64x5 hold163 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[26]),
    .clkout(net509));
 b15cbf034ar1n64x5 hold164 (.clk(n433),
    .clkout(net510));
 b15cbf034ar1n64x5 hold165 (.clk(net95),
    .clkout(net511));
 b15cbf034ar1n64x5 hold166 (.clk(net512),
    .clkout(tl_o[34]));
 b15cbf034ar1n64x5 hold167 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[30]),
    .clkout(net513));
 b15cbf034ar1n64x5 hold168 (.clk(n404),
    .clkout(net514));
 b15cbf034ar1n64x5 hold169 (.clk(net99),
    .clkout(net515));
 b15cbf034ar1n64x5 hold170 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[10]),
    .clkout(net516));
 b15cbf034ar1n64x5 hold171 (.clk(net154),
    .clkout(net517));
 b15cbf034ar1n64x5 hold172 (.clk(n411),
    .clkout(net518));
 b15cbf034ar1n64x5 hold173 (.clk(net77),
    .clkout(net519));
 b15cbf034ar1n64x5 hold174 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[3]),
    .clkout(net520));
 b15cbf034ar1n64x5 hold175 (.clk(net114),
    .clkout(net521));
 b15cbf034ar1n64x5 hold176 (.clk(net522),
    .clkout(tl_o[52]));
 b15cbf034ar1n64x5 hold177 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[7]),
    .clkout(net523));
 b15cbf034ar1n64x5 hold178 (.clk(net118),
    .clkout(net524));
 b15cbf034ar1n64x5 hold179 (.clk(net525),
    .clkout(tl_o[56]));
 b15cbf034ar1n64x5 hold180 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[33]),
    .clkout(net526));
 b15cbf034ar1n64x5 hold181 (.clk(n393),
    .clkout(net527));
 b15cbf034ar1n64x5 hold182 (.clk(net103),
    .clkout(net528));
 b15cbf034ar1n64x5 hold183 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[9]),
    .clkout(net529));
 b15cbf034ar1n64x5 hold184 (.clk(net120),
    .clkout(net530));
 b15cbf034ar1n64x5 hold185 (.clk(net531),
    .clkout(tl_o[58]));
 b15cbf034ar1n64x5 hold186 (.clk(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_storage_rdata[4]),
    .clkout(net532));
 b15cbf034ar1n64x5 hold187 (.clk(n397),
    .clkout(net533));
 b15cbf034ar1n64x5 hold188 (.clk(net143),
    .clkout(net534));
 b15cbf034ar1n64x5 hold189 (.clk(n396),
    .clkout(net535));
 b15cbf034ar1n64x5 hold190 (.clk(net106),
    .clkout(net536));
 b15cbf034ar1n64x5 hold191 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[32]),
    .clkout(net537));
 b15cbf034ar1n64x5 hold192 (.clk(n392),
    .clkout(net538));
 b15cbf034ar1n64x5 hold193 (.clk(net102),
    .clkout(net539));
 b15cbf034ar1n64x5 hold194 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[18]),
    .clkout(net540));
 b15cbf034ar1n64x5 hold195 (.clk(n421),
    .clkout(net541));
 b15cbf034ar1n64x5 hold196 (.clk(net86),
    .clkout(net542));
 b15cbf034ar1n64x5 hold197 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[38]),
    .clkout(net543));
 b15cbf034ar1n64x5 hold198 (.clk(n394),
    .clkout(net544));
 b15cbf034ar1n64x5 hold199 (.clk(net108),
    .clkout(net545));
 b15cbf034ar1n64x5 hold200 (.clk(u_tlul_adapter_sram_u_rspfifo_gen_normal_fifo_storage_rdata[35]),
    .clkout(net546));
 b15cbf034ar1n64x5 hold201 (.clk(n391),
    .clkout(net547));
 b15cbf034ar1n64x5 hold202 (.clk(net105),
    .clkout(net548));
 b15cbf034ar1n64x5 hold203 (.clk(n211),
    .clkout(net549));
 b15cbf034ar1n64x5 hold204 (.clk(u_tlul_adapter_sram_u_sramreqfifo_gen_normal_fifo_under_rst),
    .clkout(net550));
 b15cbf034ar1n64x5 hold205 (.clk(net160),
    .clkout(net551));
 b15cbf034ar1n64x5 hold206 (.clk(n362),
    .clkout(net552));
 b15cbf034ar1n64x5 hold207 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[4]),
    .clkout(net553));
 b15cbf034ar1n64x5 hold208 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[0]),
    .clkout(net554));
 b15cbf034ar1n64x5 hold209 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[5]),
    .clkout(net555));
 b15cbf034ar1n64x5 hold210 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[1]),
    .clkout(net556));
 b15cbf034ar1n64x5 hold211 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[6]),
    .clkout(net557));
 b15cbf034ar1n64x5 hold212 (.clk(u_tlul_adapter_sram_u_reqfifo_gen_normal_fifo_storage_rdata[2]),
    .clkout(net558));
 b15zdnd11an1n64x5 FILLER_0_8 ();
 b15zdnd11an1n64x5 FILLER_0_72 ();
 b15zdnd11an1n64x5 FILLER_0_136 ();
 b15zdnd11an1n64x5 FILLER_0_200 ();
 b15zdnd11an1n64x5 FILLER_0_264 ();
 b15zdnd11an1n64x5 FILLER_0_328 ();
 b15zdnd11an1n64x5 FILLER_0_392 ();
 b15zdnd11an1n64x5 FILLER_0_456 ();
 b15zdnd11an1n64x5 FILLER_0_520 ();
 b15zdnd11an1n64x5 FILLER_0_584 ();
 b15zdnd11an1n04x5 FILLER_0_648 ();
 b15zdnd00an1n02x5 FILLER_0_652 ();
 b15zdnd00an1n01x5 FILLER_0_654 ();
 b15zdnd11an1n04x5 FILLER_0_659 ();
 b15zdnd11an1n04x5 FILLER_0_670 ();
 b15zdnd00an1n02x5 FILLER_0_716 ();
 b15zdnd00an1n02x5 FILLER_0_726 ();
 b15zdnd11an1n64x5 FILLER_0_770 ();
 b15zdnd11an1n08x5 FILLER_0_834 ();
 b15zdnd00an1n02x5 FILLER_0_842 ();
 b15zdnd00an1n01x5 FILLER_0_844 ();
 b15zdnd11an1n04x5 FILLER_0_849 ();
 b15zdnd11an1n08x5 FILLER_0_857 ();
 b15zdnd00an1n02x5 FILLER_0_865 ();
 b15zdnd00an1n01x5 FILLER_0_867 ();
 b15zdnd11an1n04x5 FILLER_0_910 ();
 b15zdnd11an1n08x5 FILLER_0_918 ();
 b15zdnd00an1n02x5 FILLER_0_926 ();
 b15zdnd11an1n04x5 FILLER_0_932 ();
 b15zdnd11an1n08x5 FILLER_0_940 ();
 b15zdnd00an1n02x5 FILLER_0_948 ();
 b15zdnd00an1n01x5 FILLER_0_950 ();
 b15zdnd11an1n04x5 FILLER_0_955 ();
 b15zdnd11an1n04x5 FILLER_0_976 ();
 b15zdnd11an1n04x5 FILLER_0_1022 ();
 b15zdnd11an1n64x5 FILLER_0_1030 ();
 b15zdnd11an1n32x5 FILLER_0_1094 ();
 b15zdnd11an1n04x5 FILLER_0_1126 ();
 b15zdnd00an1n02x5 FILLER_0_1130 ();
 b15zdnd00an1n01x5 FILLER_0_1132 ();
 b15zdnd11an1n16x5 FILLER_0_1137 ();
 b15zdnd11an1n08x5 FILLER_0_1153 ();
 b15zdnd00an1n02x5 FILLER_0_1161 ();
 b15zdnd11an1n04x5 FILLER_0_1167 ();
 b15zdnd11an1n04x5 FILLER_0_1213 ();
 b15zdnd11an1n04x5 FILLER_0_1221 ();
 b15zdnd11an1n04x5 FILLER_0_1229 ();
 b15zdnd00an1n02x5 FILLER_0_1233 ();
 b15zdnd11an1n04x5 FILLER_0_1277 ();
 b15zdnd11an1n04x5 FILLER_0_1323 ();
 b15zdnd11an1n08x5 FILLER_0_1331 ();
 b15zdnd00an1n02x5 FILLER_0_1339 ();
 b15zdnd11an1n32x5 FILLER_0_1345 ();
 b15zdnd11an1n04x5 FILLER_0_1382 ();
 b15zdnd11an1n04x5 FILLER_0_1391 ();
 b15zdnd11an1n04x5 FILLER_0_1399 ();
 b15zdnd11an1n04x5 FILLER_0_1407 ();
 b15zdnd11an1n04x5 FILLER_0_1415 ();
 b15zdnd11an1n04x5 FILLER_0_1424 ();
 b15zdnd00an1n02x5 FILLER_0_1433 ();
 b15zdnd00an1n01x5 FILLER_0_1435 ();
 b15zdnd11an1n64x5 FILLER_0_1444 ();
 b15zdnd11an1n64x5 FILLER_0_1508 ();
 b15zdnd00an1n02x5 FILLER_0_1572 ();
 b15zdnd11an1n04x5 FILLER_0_1580 ();
 b15zdnd11an1n04x5 FILLER_0_1590 ();
 b15zdnd11an1n08x5 FILLER_0_1600 ();
 b15zdnd00an1n01x5 FILLER_0_1608 ();
 b15zdnd11an1n08x5 FILLER_0_1615 ();
 b15zdnd00an1n02x5 FILLER_0_1623 ();
 b15zdnd00an1n01x5 FILLER_0_1625 ();
 b15zdnd11an1n04x5 FILLER_0_1632 ();
 b15zdnd00an1n01x5 FILLER_0_1636 ();
 b15zdnd11an1n64x5 FILLER_0_1642 ();
 b15zdnd11an1n64x5 FILLER_0_1706 ();
 b15zdnd11an1n64x5 FILLER_0_1770 ();
 b15zdnd11an1n64x5 FILLER_0_1834 ();
 b15zdnd11an1n64x5 FILLER_0_1898 ();
 b15zdnd11an1n64x5 FILLER_0_1962 ();
 b15zdnd11an1n64x5 FILLER_0_2026 ();
 b15zdnd11an1n64x5 FILLER_0_2090 ();
 b15zdnd11an1n64x5 FILLER_0_2162 ();
 b15zdnd11an1n32x5 FILLER_0_2226 ();
 b15zdnd11an1n16x5 FILLER_0_2258 ();
 b15zdnd00an1n02x5 FILLER_0_2274 ();
 b15zdnd11an1n64x5 FILLER_1_0 ();
 b15zdnd11an1n64x5 FILLER_1_64 ();
 b15zdnd11an1n64x5 FILLER_1_128 ();
 b15zdnd11an1n64x5 FILLER_1_192 ();
 b15zdnd11an1n64x5 FILLER_1_256 ();
 b15zdnd11an1n64x5 FILLER_1_320 ();
 b15zdnd11an1n64x5 FILLER_1_384 ();
 b15zdnd11an1n64x5 FILLER_1_448 ();
 b15zdnd11an1n64x5 FILLER_1_512 ();
 b15zdnd11an1n64x5 FILLER_1_576 ();
 b15zdnd11an1n16x5 FILLER_1_640 ();
 b15zdnd00an1n02x5 FILLER_1_656 ();
 b15zdnd11an1n04x5 FILLER_1_700 ();
 b15zdnd11an1n04x5 FILLER_1_746 ();
 b15zdnd11an1n64x5 FILLER_1_761 ();
 b15zdnd11an1n16x5 FILLER_1_825 ();
 b15zdnd11an1n08x5 FILLER_1_841 ();
 b15zdnd11an1n04x5 FILLER_1_849 ();
 b15zdnd00an1n01x5 FILLER_1_853 ();
 b15zdnd11an1n64x5 FILLER_1_896 ();
 b15zdnd11an1n04x5 FILLER_1_960 ();
 b15zdnd11an1n04x5 FILLER_1_1006 ();
 b15zdnd11an1n64x5 FILLER_1_1030 ();
 b15zdnd11an1n64x5 FILLER_1_1094 ();
 b15zdnd11an1n16x5 FILLER_1_1158 ();
 b15zdnd11an1n08x5 FILLER_1_1174 ();
 b15zdnd00an1n01x5 FILLER_1_1182 ();
 b15zdnd11an1n04x5 FILLER_1_1187 ();
 b15zdnd11an1n04x5 FILLER_1_1195 ();
 b15zdnd11an1n04x5 FILLER_1_1203 ();
 b15zdnd11an1n16x5 FILLER_1_1211 ();
 b15zdnd00an1n02x5 FILLER_1_1227 ();
 b15zdnd00an1n01x5 FILLER_1_1229 ();
 b15zdnd11an1n08x5 FILLER_1_1234 ();
 b15zdnd00an1n02x5 FILLER_1_1242 ();
 b15zdnd00an1n01x5 FILLER_1_1244 ();
 b15zdnd11an1n16x5 FILLER_1_1287 ();
 b15zdnd11an1n04x5 FILLER_1_1303 ();
 b15zdnd11an1n64x5 FILLER_1_1312 ();
 b15zdnd11an1n04x5 FILLER_1_1376 ();
 b15zdnd00an1n02x5 FILLER_1_1380 ();
 b15zdnd00an1n01x5 FILLER_1_1382 ();
 b15zdnd11an1n04x5 FILLER_1_1388 ();
 b15zdnd00an1n01x5 FILLER_1_1392 ();
 b15zdnd11an1n04x5 FILLER_1_1398 ();
 b15zdnd11an1n64x5 FILLER_1_1406 ();
 b15zdnd11an1n64x5 FILLER_1_1470 ();
 b15zdnd11an1n64x5 FILLER_1_1534 ();
 b15zdnd11an1n64x5 FILLER_1_1598 ();
 b15zdnd11an1n64x5 FILLER_1_1662 ();
 b15zdnd11an1n64x5 FILLER_1_1726 ();
 b15zdnd11an1n64x5 FILLER_1_1790 ();
 b15zdnd11an1n64x5 FILLER_1_1854 ();
 b15zdnd11an1n64x5 FILLER_1_1918 ();
 b15zdnd11an1n64x5 FILLER_1_1982 ();
 b15zdnd11an1n64x5 FILLER_1_2046 ();
 b15zdnd11an1n64x5 FILLER_1_2110 ();
 b15zdnd11an1n64x5 FILLER_1_2174 ();
 b15zdnd11an1n32x5 FILLER_1_2238 ();
 b15zdnd11an1n08x5 FILLER_1_2270 ();
 b15zdnd11an1n04x5 FILLER_1_2278 ();
 b15zdnd00an1n02x5 FILLER_1_2282 ();
 b15zdnd11an1n64x5 FILLER_2_8 ();
 b15zdnd11an1n64x5 FILLER_2_72 ();
 b15zdnd11an1n64x5 FILLER_2_136 ();
 b15zdnd11an1n64x5 FILLER_2_200 ();
 b15zdnd11an1n64x5 FILLER_2_264 ();
 b15zdnd11an1n64x5 FILLER_2_328 ();
 b15zdnd11an1n64x5 FILLER_2_392 ();
 b15zdnd11an1n64x5 FILLER_2_456 ();
 b15zdnd11an1n64x5 FILLER_2_520 ();
 b15zdnd11an1n64x5 FILLER_2_584 ();
 b15zdnd00an1n02x5 FILLER_2_648 ();
 b15zdnd00an1n01x5 FILLER_2_650 ();
 b15zdnd11an1n04x5 FILLER_2_655 ();
 b15zdnd11an1n04x5 FILLER_2_701 ();
 b15zdnd00an1n02x5 FILLER_2_705 ();
 b15zdnd11an1n04x5 FILLER_2_714 ();
 b15zdnd00an1n02x5 FILLER_2_726 ();
 b15zdnd11an1n64x5 FILLER_2_732 ();
 b15zdnd11an1n64x5 FILLER_2_796 ();
 b15zdnd11an1n08x5 FILLER_2_860 ();
 b15zdnd11an1n04x5 FILLER_2_868 ();
 b15zdnd11an1n64x5 FILLER_2_883 ();
 b15zdnd11an1n16x5 FILLER_2_947 ();
 b15zdnd00an1n02x5 FILLER_2_963 ();
 b15zdnd00an1n01x5 FILLER_2_965 ();
 b15zdnd11an1n08x5 FILLER_2_986 ();
 b15zdnd00an1n02x5 FILLER_2_994 ();
 b15zdnd00an1n01x5 FILLER_2_996 ();
 b15zdnd11an1n16x5 FILLER_2_1017 ();
 b15zdnd00an1n02x5 FILLER_2_1033 ();
 b15zdnd00an1n01x5 FILLER_2_1035 ();
 b15zdnd11an1n64x5 FILLER_2_1053 ();
 b15zdnd11an1n64x5 FILLER_2_1117 ();
 b15zdnd11an1n32x5 FILLER_2_1181 ();
 b15zdnd11an1n16x5 FILLER_2_1213 ();
 b15zdnd00an1n02x5 FILLER_2_1229 ();
 b15zdnd00an1n01x5 FILLER_2_1231 ();
 b15zdnd11an1n04x5 FILLER_2_1236 ();
 b15zdnd00an1n02x5 FILLER_2_1240 ();
 b15zdnd00an1n01x5 FILLER_2_1242 ();
 b15zdnd11an1n04x5 FILLER_2_1247 ();
 b15zdnd11an1n04x5 FILLER_2_1255 ();
 b15zdnd11an1n64x5 FILLER_2_1263 ();
 b15zdnd11an1n64x5 FILLER_2_1327 ();
 b15zdnd11an1n04x5 FILLER_2_1391 ();
 b15zdnd00an1n01x5 FILLER_2_1395 ();
 b15zdnd11an1n04x5 FILLER_2_1400 ();
 b15zdnd11an1n64x5 FILLER_2_1408 ();
 b15zdnd11an1n64x5 FILLER_2_1472 ();
 b15zdnd11an1n32x5 FILLER_2_1536 ();
 b15zdnd11an1n16x5 FILLER_2_1568 ();
 b15zdnd11an1n08x5 FILLER_2_1584 ();
 b15zdnd11an1n64x5 FILLER_2_1598 ();
 b15zdnd11an1n64x5 FILLER_2_1662 ();
 b15zdnd11an1n64x5 FILLER_2_1726 ();
 b15zdnd11an1n64x5 FILLER_2_1790 ();
 b15zdnd11an1n64x5 FILLER_2_1854 ();
 b15zdnd11an1n64x5 FILLER_2_1918 ();
 b15zdnd11an1n64x5 FILLER_2_1982 ();
 b15zdnd11an1n64x5 FILLER_2_2046 ();
 b15zdnd11an1n32x5 FILLER_2_2110 ();
 b15zdnd11an1n08x5 FILLER_2_2142 ();
 b15zdnd11an1n04x5 FILLER_2_2150 ();
 b15zdnd11an1n64x5 FILLER_2_2162 ();
 b15zdnd11an1n32x5 FILLER_2_2226 ();
 b15zdnd11an1n16x5 FILLER_2_2258 ();
 b15zdnd00an1n02x5 FILLER_2_2274 ();
 b15zdnd11an1n64x5 FILLER_3_0 ();
 b15zdnd11an1n64x5 FILLER_3_64 ();
 b15zdnd11an1n64x5 FILLER_3_128 ();
 b15zdnd11an1n64x5 FILLER_3_192 ();
 b15zdnd11an1n64x5 FILLER_3_256 ();
 b15zdnd11an1n64x5 FILLER_3_320 ();
 b15zdnd11an1n64x5 FILLER_3_384 ();
 b15zdnd11an1n64x5 FILLER_3_448 ();
 b15zdnd11an1n64x5 FILLER_3_512 ();
 b15zdnd11an1n64x5 FILLER_3_576 ();
 b15zdnd11an1n32x5 FILLER_3_640 ();
 b15zdnd00an1n02x5 FILLER_3_672 ();
 b15zdnd00an1n01x5 FILLER_3_674 ();
 b15zdnd11an1n08x5 FILLER_3_682 ();
 b15zdnd11an1n08x5 FILLER_3_701 ();
 b15zdnd00an1n02x5 FILLER_3_709 ();
 b15zdnd00an1n01x5 FILLER_3_711 ();
 b15zdnd11an1n04x5 FILLER_3_719 ();
 b15zdnd11an1n64x5 FILLER_3_727 ();
 b15zdnd11an1n64x5 FILLER_3_791 ();
 b15zdnd11an1n64x5 FILLER_3_855 ();
 b15zdnd11an1n32x5 FILLER_3_919 ();
 b15zdnd11an1n16x5 FILLER_3_951 ();
 b15zdnd11an1n04x5 FILLER_3_967 ();
 b15zdnd00an1n02x5 FILLER_3_971 ();
 b15zdnd00an1n01x5 FILLER_3_973 ();
 b15zdnd11an1n32x5 FILLER_3_978 ();
 b15zdnd11an1n16x5 FILLER_3_1010 ();
 b15zdnd11an1n04x5 FILLER_3_1026 ();
 b15zdnd00an1n02x5 FILLER_3_1030 ();
 b15zdnd00an1n01x5 FILLER_3_1032 ();
 b15zdnd11an1n64x5 FILLER_3_1047 ();
 b15zdnd11an1n64x5 FILLER_3_1111 ();
 b15zdnd11an1n64x5 FILLER_3_1175 ();
 b15zdnd11an1n64x5 FILLER_3_1239 ();
 b15zdnd11an1n64x5 FILLER_3_1303 ();
 b15zdnd11an1n16x5 FILLER_3_1367 ();
 b15zdnd11an1n08x5 FILLER_3_1383 ();
 b15zdnd00an1n02x5 FILLER_3_1391 ();
 b15zdnd11an1n64x5 FILLER_3_1397 ();
 b15zdnd11an1n64x5 FILLER_3_1461 ();
 b15zdnd11an1n64x5 FILLER_3_1525 ();
 b15zdnd11an1n64x5 FILLER_3_1589 ();
 b15zdnd11an1n64x5 FILLER_3_1653 ();
 b15zdnd11an1n64x5 FILLER_3_1717 ();
 b15zdnd11an1n64x5 FILLER_3_1781 ();
 b15zdnd11an1n64x5 FILLER_3_1845 ();
 b15zdnd11an1n64x5 FILLER_3_1909 ();
 b15zdnd11an1n64x5 FILLER_3_1973 ();
 b15zdnd11an1n64x5 FILLER_3_2037 ();
 b15zdnd11an1n64x5 FILLER_3_2101 ();
 b15zdnd11an1n64x5 FILLER_3_2165 ();
 b15zdnd11an1n32x5 FILLER_3_2229 ();
 b15zdnd11an1n16x5 FILLER_3_2261 ();
 b15zdnd11an1n04x5 FILLER_3_2277 ();
 b15zdnd00an1n02x5 FILLER_3_2281 ();
 b15zdnd00an1n01x5 FILLER_3_2283 ();
 b15zdnd11an1n64x5 FILLER_4_8 ();
 b15zdnd11an1n64x5 FILLER_4_72 ();
 b15zdnd11an1n64x5 FILLER_4_136 ();
 b15zdnd11an1n64x5 FILLER_4_200 ();
 b15zdnd11an1n64x5 FILLER_4_264 ();
 b15zdnd11an1n64x5 FILLER_4_328 ();
 b15zdnd11an1n64x5 FILLER_4_392 ();
 b15zdnd11an1n64x5 FILLER_4_456 ();
 b15zdnd11an1n64x5 FILLER_4_520 ();
 b15zdnd11an1n64x5 FILLER_4_584 ();
 b15zdnd11an1n32x5 FILLER_4_648 ();
 b15zdnd11an1n04x5 FILLER_4_680 ();
 b15zdnd00an1n01x5 FILLER_4_684 ();
 b15zdnd11an1n08x5 FILLER_4_689 ();
 b15zdnd11an1n04x5 FILLER_4_697 ();
 b15zdnd00an1n01x5 FILLER_4_701 ();
 b15zdnd11an1n08x5 FILLER_4_709 ();
 b15zdnd00an1n01x5 FILLER_4_717 ();
 b15zdnd11an1n64x5 FILLER_4_726 ();
 b15zdnd11an1n64x5 FILLER_4_790 ();
 b15zdnd11an1n64x5 FILLER_4_854 ();
 b15zdnd11an1n64x5 FILLER_4_918 ();
 b15zdnd11an1n64x5 FILLER_4_982 ();
 b15zdnd11an1n64x5 FILLER_4_1046 ();
 b15zdnd11an1n64x5 FILLER_4_1110 ();
 b15zdnd11an1n64x5 FILLER_4_1174 ();
 b15zdnd11an1n64x5 FILLER_4_1238 ();
 b15zdnd11an1n64x5 FILLER_4_1302 ();
 b15zdnd11an1n64x5 FILLER_4_1366 ();
 b15zdnd11an1n32x5 FILLER_4_1430 ();
 b15zdnd11an1n16x5 FILLER_4_1462 ();
 b15zdnd11an1n08x5 FILLER_4_2265 ();
 b15zdnd00an1n02x5 FILLER_4_2273 ();
 b15zdnd00an1n01x5 FILLER_4_2275 ();
 b15zdnd11an1n64x5 FILLER_5_0 ();
 b15zdnd11an1n64x5 FILLER_5_64 ();
 b15zdnd11an1n64x5 FILLER_5_128 ();
 b15zdnd11an1n64x5 FILLER_5_192 ();
 b15zdnd11an1n64x5 FILLER_5_256 ();
 b15zdnd11an1n64x5 FILLER_5_320 ();
 b15zdnd11an1n64x5 FILLER_5_384 ();
 b15zdnd11an1n64x5 FILLER_5_448 ();
 b15zdnd11an1n64x5 FILLER_5_512 ();
 b15zdnd11an1n64x5 FILLER_5_576 ();
 b15zdnd11an1n64x5 FILLER_5_640 ();
 b15zdnd11an1n64x5 FILLER_5_704 ();
 b15zdnd11an1n64x5 FILLER_5_768 ();
 b15zdnd11an1n64x5 FILLER_5_832 ();
 b15zdnd11an1n64x5 FILLER_5_896 ();
 b15zdnd11an1n64x5 FILLER_5_960 ();
 b15zdnd11an1n64x5 FILLER_5_1024 ();
 b15zdnd11an1n64x5 FILLER_5_1088 ();
 b15zdnd11an1n64x5 FILLER_5_1152 ();
 b15zdnd11an1n64x5 FILLER_5_1216 ();
 b15zdnd11an1n64x5 FILLER_5_1280 ();
 b15zdnd11an1n64x5 FILLER_5_1344 ();
 b15zdnd11an1n64x5 FILLER_5_1408 ();
 b15zdnd11an1n08x5 FILLER_5_1472 ();
 b15zdnd11an1n04x5 FILLER_5_1480 ();
 b15zdnd00an1n02x5 FILLER_5_1484 ();
 b15zdnd11an1n16x5 FILLER_5_2257 ();
 b15zdnd11an1n08x5 FILLER_5_2273 ();
 b15zdnd00an1n02x5 FILLER_5_2281 ();
 b15zdnd00an1n01x5 FILLER_5_2283 ();
 b15zdnd11an1n64x5 FILLER_6_8 ();
 b15zdnd11an1n64x5 FILLER_6_72 ();
 b15zdnd11an1n64x5 FILLER_6_136 ();
 b15zdnd11an1n64x5 FILLER_6_200 ();
 b15zdnd11an1n64x5 FILLER_6_264 ();
 b15zdnd11an1n64x5 FILLER_6_328 ();
 b15zdnd11an1n64x5 FILLER_6_392 ();
 b15zdnd11an1n64x5 FILLER_6_456 ();
 b15zdnd11an1n64x5 FILLER_6_520 ();
 b15zdnd11an1n64x5 FILLER_6_584 ();
 b15zdnd11an1n64x5 FILLER_6_648 ();
 b15zdnd11an1n04x5 FILLER_6_712 ();
 b15zdnd00an1n02x5 FILLER_6_716 ();
 b15zdnd11an1n64x5 FILLER_6_726 ();
 b15zdnd11an1n64x5 FILLER_6_790 ();
 b15zdnd11an1n64x5 FILLER_6_854 ();
 b15zdnd11an1n64x5 FILLER_6_918 ();
 b15zdnd11an1n64x5 FILLER_6_982 ();
 b15zdnd11an1n64x5 FILLER_6_1046 ();
 b15zdnd11an1n64x5 FILLER_6_1110 ();
 b15zdnd11an1n64x5 FILLER_6_1174 ();
 b15zdnd11an1n64x5 FILLER_6_1238 ();
 b15zdnd11an1n64x5 FILLER_6_1302 ();
 b15zdnd11an1n64x5 FILLER_6_1366 ();
 b15zdnd11an1n32x5 FILLER_6_1430 ();
 b15zdnd11an1n16x5 FILLER_6_1462 ();
 b15zdnd11an1n08x5 FILLER_6_2265 ();
 b15zdnd00an1n02x5 FILLER_6_2273 ();
 b15zdnd00an1n01x5 FILLER_6_2275 ();
 b15zdnd11an1n64x5 FILLER_7_0 ();
 b15zdnd11an1n64x5 FILLER_7_64 ();
 b15zdnd11an1n64x5 FILLER_7_128 ();
 b15zdnd11an1n64x5 FILLER_7_192 ();
 b15zdnd11an1n64x5 FILLER_7_256 ();
 b15zdnd11an1n64x5 FILLER_7_320 ();
 b15zdnd11an1n64x5 FILLER_7_384 ();
 b15zdnd11an1n64x5 FILLER_7_448 ();
 b15zdnd11an1n64x5 FILLER_7_512 ();
 b15zdnd11an1n64x5 FILLER_7_576 ();
 b15zdnd11an1n64x5 FILLER_7_640 ();
 b15zdnd11an1n64x5 FILLER_7_704 ();
 b15zdnd11an1n64x5 FILLER_7_768 ();
 b15zdnd11an1n64x5 FILLER_7_832 ();
 b15zdnd11an1n16x5 FILLER_7_896 ();
 b15zdnd11an1n04x5 FILLER_7_912 ();
 b15zdnd11an1n64x5 FILLER_7_958 ();
 b15zdnd11an1n64x5 FILLER_7_1022 ();
 b15zdnd11an1n32x5 FILLER_7_1086 ();
 b15zdnd00an1n02x5 FILLER_7_1118 ();
 b15zdnd11an1n64x5 FILLER_7_1162 ();
 b15zdnd11an1n64x5 FILLER_7_1226 ();
 b15zdnd11an1n64x5 FILLER_7_1290 ();
 b15zdnd11an1n64x5 FILLER_7_1354 ();
 b15zdnd11an1n64x5 FILLER_7_1418 ();
 b15zdnd11an1n04x5 FILLER_7_1482 ();
 b15zdnd11an1n16x5 FILLER_7_2257 ();
 b15zdnd11an1n08x5 FILLER_7_2273 ();
 b15zdnd00an1n02x5 FILLER_7_2281 ();
 b15zdnd00an1n01x5 FILLER_7_2283 ();
 b15zdnd11an1n64x5 FILLER_8_8 ();
 b15zdnd11an1n64x5 FILLER_8_72 ();
 b15zdnd11an1n64x5 FILLER_8_136 ();
 b15zdnd11an1n64x5 FILLER_8_200 ();
 b15zdnd11an1n64x5 FILLER_8_264 ();
 b15zdnd11an1n64x5 FILLER_8_328 ();
 b15zdnd11an1n64x5 FILLER_8_392 ();
 b15zdnd11an1n64x5 FILLER_8_456 ();
 b15zdnd11an1n64x5 FILLER_8_520 ();
 b15zdnd11an1n64x5 FILLER_8_584 ();
 b15zdnd11an1n64x5 FILLER_8_648 ();
 b15zdnd11an1n04x5 FILLER_8_712 ();
 b15zdnd00an1n02x5 FILLER_8_716 ();
 b15zdnd11an1n64x5 FILLER_8_726 ();
 b15zdnd11an1n08x5 FILLER_8_790 ();
 b15zdnd00an1n02x5 FILLER_8_798 ();
 b15zdnd00an1n01x5 FILLER_8_800 ();
 b15zdnd11an1n16x5 FILLER_8_843 ();
 b15zdnd11an1n08x5 FILLER_8_859 ();
 b15zdnd11an1n16x5 FILLER_8_909 ();
 b15zdnd11an1n04x5 FILLER_8_925 ();
 b15zdnd00an1n01x5 FILLER_8_929 ();
 b15zdnd11an1n64x5 FILLER_8_972 ();
 b15zdnd11an1n64x5 FILLER_8_1036 ();
 b15zdnd11an1n32x5 FILLER_8_1100 ();
 b15zdnd11an1n08x5 FILLER_8_1132 ();
 b15zdnd11an1n04x5 FILLER_8_1140 ();
 b15zdnd00an1n02x5 FILLER_8_1144 ();
 b15zdnd11an1n16x5 FILLER_8_1188 ();
 b15zdnd00an1n02x5 FILLER_8_1204 ();
 b15zdnd00an1n01x5 FILLER_8_1206 ();
 b15zdnd11an1n64x5 FILLER_8_1249 ();
 b15zdnd11an1n64x5 FILLER_8_1313 ();
 b15zdnd11an1n64x5 FILLER_8_1377 ();
 b15zdnd11an1n32x5 FILLER_8_1441 ();
 b15zdnd11an1n04x5 FILLER_8_1473 ();
 b15zdnd00an1n01x5 FILLER_8_1477 ();
 b15zdnd11an1n08x5 FILLER_8_2265 ();
 b15zdnd00an1n02x5 FILLER_8_2273 ();
 b15zdnd00an1n01x5 FILLER_8_2275 ();
 b15zdnd11an1n64x5 FILLER_9_0 ();
 b15zdnd11an1n64x5 FILLER_9_64 ();
 b15zdnd11an1n64x5 FILLER_9_128 ();
 b15zdnd11an1n64x5 FILLER_9_192 ();
 b15zdnd11an1n64x5 FILLER_9_256 ();
 b15zdnd11an1n64x5 FILLER_9_320 ();
 b15zdnd11an1n64x5 FILLER_9_384 ();
 b15zdnd11an1n64x5 FILLER_9_448 ();
 b15zdnd11an1n64x5 FILLER_9_512 ();
 b15zdnd11an1n64x5 FILLER_9_576 ();
 b15zdnd11an1n64x5 FILLER_9_640 ();
 b15zdnd11an1n64x5 FILLER_9_704 ();
 b15zdnd11an1n64x5 FILLER_9_768 ();
 b15zdnd00an1n01x5 FILLER_9_832 ();
 b15zdnd11an1n08x5 FILLER_9_875 ();
 b15zdnd11an1n04x5 FILLER_9_883 ();
 b15zdnd11an1n16x5 FILLER_9_929 ();
 b15zdnd11an1n04x5 FILLER_9_987 ();
 b15zdnd00an1n01x5 FILLER_9_991 ();
 b15zdnd11an1n16x5 FILLER_9_1034 ();
 b15zdnd11an1n08x5 FILLER_9_1050 ();
 b15zdnd00an1n02x5 FILLER_9_1058 ();
 b15zdnd00an1n01x5 FILLER_9_1060 ();
 b15zdnd11an1n32x5 FILLER_9_1103 ();
 b15zdnd11an1n04x5 FILLER_9_1135 ();
 b15zdnd00an1n02x5 FILLER_9_1139 ();
 b15zdnd11an1n16x5 FILLER_9_1183 ();
 b15zdnd11an1n64x5 FILLER_9_1241 ();
 b15zdnd11an1n64x5 FILLER_9_1305 ();
 b15zdnd11an1n64x5 FILLER_9_1369 ();
 b15zdnd11an1n32x5 FILLER_9_1433 ();
 b15zdnd11an1n16x5 FILLER_9_1465 ();
 b15zdnd11an1n04x5 FILLER_9_1481 ();
 b15zdnd00an1n01x5 FILLER_9_1485 ();
 b15zdnd11an1n16x5 FILLER_9_2257 ();
 b15zdnd11an1n08x5 FILLER_9_2273 ();
 b15zdnd00an1n02x5 FILLER_9_2281 ();
 b15zdnd00an1n01x5 FILLER_9_2283 ();
 b15zdnd11an1n64x5 FILLER_10_8 ();
 b15zdnd11an1n64x5 FILLER_10_72 ();
 b15zdnd11an1n64x5 FILLER_10_136 ();
 b15zdnd11an1n64x5 FILLER_10_200 ();
 b15zdnd11an1n64x5 FILLER_10_264 ();
 b15zdnd11an1n64x5 FILLER_10_328 ();
 b15zdnd11an1n64x5 FILLER_10_392 ();
 b15zdnd11an1n64x5 FILLER_10_456 ();
 b15zdnd11an1n64x5 FILLER_10_520 ();
 b15zdnd11an1n64x5 FILLER_10_584 ();
 b15zdnd11an1n64x5 FILLER_10_648 ();
 b15zdnd11an1n04x5 FILLER_10_712 ();
 b15zdnd00an1n02x5 FILLER_10_716 ();
 b15zdnd11an1n64x5 FILLER_10_726 ();
 b15zdnd11an1n64x5 FILLER_10_790 ();
 b15zdnd11an1n32x5 FILLER_10_854 ();
 b15zdnd11an1n16x5 FILLER_10_886 ();
 b15zdnd11an1n08x5 FILLER_10_902 ();
 b15zdnd00an1n01x5 FILLER_10_910 ();
 b15zdnd11an1n32x5 FILLER_10_953 ();
 b15zdnd11an1n08x5 FILLER_10_985 ();
 b15zdnd00an1n01x5 FILLER_10_993 ();
 b15zdnd11an1n32x5 FILLER_10_1036 ();
 b15zdnd11an1n16x5 FILLER_10_1068 ();
 b15zdnd11an1n04x5 FILLER_10_1126 ();
 b15zdnd11an1n16x5 FILLER_10_1172 ();
 b15zdnd11an1n08x5 FILLER_10_1188 ();
 b15zdnd00an1n01x5 FILLER_10_1196 ();
 b15zdnd11an1n04x5 FILLER_10_1239 ();
 b15zdnd11an1n64x5 FILLER_10_1285 ();
 b15zdnd11an1n64x5 FILLER_10_1349 ();
 b15zdnd11an1n64x5 FILLER_10_1413 ();
 b15zdnd00an1n01x5 FILLER_10_1477 ();
 b15zdnd11an1n08x5 FILLER_10_2265 ();
 b15zdnd00an1n02x5 FILLER_10_2273 ();
 b15zdnd00an1n01x5 FILLER_10_2275 ();
 b15zdnd11an1n64x5 FILLER_11_0 ();
 b15zdnd11an1n64x5 FILLER_11_64 ();
 b15zdnd11an1n64x5 FILLER_11_128 ();
 b15zdnd11an1n64x5 FILLER_11_192 ();
 b15zdnd11an1n64x5 FILLER_11_256 ();
 b15zdnd11an1n64x5 FILLER_11_320 ();
 b15zdnd11an1n64x5 FILLER_11_384 ();
 b15zdnd11an1n64x5 FILLER_11_448 ();
 b15zdnd11an1n64x5 FILLER_11_512 ();
 b15zdnd11an1n64x5 FILLER_11_576 ();
 b15zdnd11an1n64x5 FILLER_11_640 ();
 b15zdnd11an1n64x5 FILLER_11_704 ();
 b15zdnd11an1n64x5 FILLER_11_768 ();
 b15zdnd11an1n64x5 FILLER_11_832 ();
 b15zdnd11an1n64x5 FILLER_11_896 ();
 b15zdnd11an1n64x5 FILLER_11_960 ();
 b15zdnd11an1n64x5 FILLER_11_1024 ();
 b15zdnd11an1n64x5 FILLER_11_1088 ();
 b15zdnd11an1n64x5 FILLER_11_1152 ();
 b15zdnd11an1n64x5 FILLER_11_1216 ();
 b15zdnd11an1n64x5 FILLER_11_1280 ();
 b15zdnd11an1n64x5 FILLER_11_1344 ();
 b15zdnd11an1n64x5 FILLER_11_1408 ();
 b15zdnd11an1n08x5 FILLER_11_1472 ();
 b15zdnd11an1n04x5 FILLER_11_1480 ();
 b15zdnd00an1n02x5 FILLER_11_1484 ();
 b15zdnd11an1n16x5 FILLER_11_2257 ();
 b15zdnd11an1n08x5 FILLER_11_2273 ();
 b15zdnd00an1n02x5 FILLER_11_2281 ();
 b15zdnd00an1n01x5 FILLER_11_2283 ();
 b15zdnd11an1n64x5 FILLER_12_8 ();
 b15zdnd11an1n64x5 FILLER_12_72 ();
 b15zdnd11an1n64x5 FILLER_12_136 ();
 b15zdnd11an1n64x5 FILLER_12_200 ();
 b15zdnd11an1n64x5 FILLER_12_264 ();
 b15zdnd11an1n64x5 FILLER_12_328 ();
 b15zdnd11an1n64x5 FILLER_12_392 ();
 b15zdnd11an1n64x5 FILLER_12_456 ();
 b15zdnd11an1n64x5 FILLER_12_520 ();
 b15zdnd11an1n64x5 FILLER_12_584 ();
 b15zdnd11an1n64x5 FILLER_12_648 ();
 b15zdnd11an1n04x5 FILLER_12_712 ();
 b15zdnd00an1n02x5 FILLER_12_716 ();
 b15zdnd11an1n64x5 FILLER_12_726 ();
 b15zdnd11an1n64x5 FILLER_12_790 ();
 b15zdnd11an1n64x5 FILLER_12_854 ();
 b15zdnd11an1n64x5 FILLER_12_918 ();
 b15zdnd11an1n64x5 FILLER_12_982 ();
 b15zdnd11an1n64x5 FILLER_12_1046 ();
 b15zdnd11an1n64x5 FILLER_12_1110 ();
 b15zdnd11an1n64x5 FILLER_12_1174 ();
 b15zdnd11an1n64x5 FILLER_12_1238 ();
 b15zdnd11an1n64x5 FILLER_12_1302 ();
 b15zdnd11an1n64x5 FILLER_12_1366 ();
 b15zdnd11an1n32x5 FILLER_12_1430 ();
 b15zdnd11an1n16x5 FILLER_12_1462 ();
 b15zdnd11an1n08x5 FILLER_12_2265 ();
 b15zdnd00an1n02x5 FILLER_12_2273 ();
 b15zdnd00an1n01x5 FILLER_12_2275 ();
 b15zdnd11an1n64x5 FILLER_13_0 ();
 b15zdnd11an1n64x5 FILLER_13_64 ();
 b15zdnd11an1n64x5 FILLER_13_128 ();
 b15zdnd11an1n64x5 FILLER_13_192 ();
 b15zdnd11an1n64x5 FILLER_13_256 ();
 b15zdnd11an1n64x5 FILLER_13_320 ();
 b15zdnd11an1n64x5 FILLER_13_384 ();
 b15zdnd11an1n64x5 FILLER_13_448 ();
 b15zdnd11an1n64x5 FILLER_13_512 ();
 b15zdnd11an1n64x5 FILLER_13_576 ();
 b15zdnd11an1n64x5 FILLER_13_640 ();
 b15zdnd11an1n64x5 FILLER_13_704 ();
 b15zdnd11an1n64x5 FILLER_13_768 ();
 b15zdnd11an1n64x5 FILLER_13_832 ();
 b15zdnd11an1n64x5 FILLER_13_896 ();
 b15zdnd11an1n64x5 FILLER_13_960 ();
 b15zdnd11an1n64x5 FILLER_13_1024 ();
 b15zdnd11an1n64x5 FILLER_13_1088 ();
 b15zdnd11an1n64x5 FILLER_13_1152 ();
 b15zdnd11an1n64x5 FILLER_13_1216 ();
 b15zdnd11an1n64x5 FILLER_13_1280 ();
 b15zdnd11an1n64x5 FILLER_13_1344 ();
 b15zdnd11an1n64x5 FILLER_13_1408 ();
 b15zdnd11an1n08x5 FILLER_13_1472 ();
 b15zdnd11an1n04x5 FILLER_13_1480 ();
 b15zdnd00an1n02x5 FILLER_13_1484 ();
 b15zdnd11an1n16x5 FILLER_13_2257 ();
 b15zdnd11an1n08x5 FILLER_13_2273 ();
 b15zdnd00an1n02x5 FILLER_13_2281 ();
 b15zdnd00an1n01x5 FILLER_13_2283 ();
 b15zdnd11an1n64x5 FILLER_14_8 ();
 b15zdnd11an1n64x5 FILLER_14_72 ();
 b15zdnd11an1n64x5 FILLER_14_136 ();
 b15zdnd11an1n64x5 FILLER_14_200 ();
 b15zdnd11an1n64x5 FILLER_14_264 ();
 b15zdnd11an1n64x5 FILLER_14_328 ();
 b15zdnd11an1n64x5 FILLER_14_392 ();
 b15zdnd11an1n64x5 FILLER_14_456 ();
 b15zdnd11an1n64x5 FILLER_14_520 ();
 b15zdnd11an1n64x5 FILLER_14_584 ();
 b15zdnd11an1n64x5 FILLER_14_648 ();
 b15zdnd11an1n04x5 FILLER_14_712 ();
 b15zdnd00an1n02x5 FILLER_14_716 ();
 b15zdnd11an1n64x5 FILLER_14_726 ();
 b15zdnd11an1n64x5 FILLER_14_790 ();
 b15zdnd11an1n64x5 FILLER_14_854 ();
 b15zdnd11an1n64x5 FILLER_14_918 ();
 b15zdnd11an1n64x5 FILLER_14_982 ();
 b15zdnd11an1n64x5 FILLER_14_1046 ();
 b15zdnd11an1n64x5 FILLER_14_1110 ();
 b15zdnd11an1n64x5 FILLER_14_1174 ();
 b15zdnd11an1n64x5 FILLER_14_1238 ();
 b15zdnd11an1n64x5 FILLER_14_1302 ();
 b15zdnd11an1n64x5 FILLER_14_1366 ();
 b15zdnd11an1n32x5 FILLER_14_1430 ();
 b15zdnd11an1n16x5 FILLER_14_1462 ();
 b15zdnd11an1n08x5 FILLER_14_2265 ();
 b15zdnd00an1n02x5 FILLER_14_2273 ();
 b15zdnd00an1n01x5 FILLER_14_2275 ();
 b15zdnd11an1n64x5 FILLER_15_0 ();
 b15zdnd11an1n64x5 FILLER_15_64 ();
 b15zdnd11an1n64x5 FILLER_15_128 ();
 b15zdnd11an1n64x5 FILLER_15_192 ();
 b15zdnd11an1n64x5 FILLER_15_256 ();
 b15zdnd11an1n64x5 FILLER_15_320 ();
 b15zdnd11an1n64x5 FILLER_15_384 ();
 b15zdnd11an1n64x5 FILLER_15_448 ();
 b15zdnd11an1n64x5 FILLER_15_512 ();
 b15zdnd11an1n64x5 FILLER_15_576 ();
 b15zdnd11an1n08x5 FILLER_15_640 ();
 b15zdnd11an1n04x5 FILLER_15_648 ();
 b15zdnd00an1n02x5 FILLER_15_652 ();
 b15zdnd00an1n01x5 FILLER_15_654 ();
 b15zdnd11an1n08x5 FILLER_15_658 ();
 b15zdnd11an1n04x5 FILLER_15_666 ();
 b15zdnd00an1n02x5 FILLER_15_670 ();
 b15zdnd00an1n01x5 FILLER_15_672 ();
 b15zdnd11an1n04x5 FILLER_15_676 ();
 b15zdnd11an1n04x5 FILLER_15_683 ();
 b15zdnd11an1n08x5 FILLER_15_690 ();
 b15zdnd00an1n02x5 FILLER_15_698 ();
 b15zdnd00an1n01x5 FILLER_15_700 ();
 b15zdnd11an1n04x5 FILLER_15_704 ();
 b15zdnd00an1n01x5 FILLER_15_708 ();
 b15zdnd11an1n64x5 FILLER_15_712 ();
 b15zdnd11an1n64x5 FILLER_15_776 ();
 b15zdnd11an1n64x5 FILLER_15_840 ();
 b15zdnd11an1n64x5 FILLER_15_904 ();
 b15zdnd11an1n64x5 FILLER_15_968 ();
 b15zdnd11an1n64x5 FILLER_15_1032 ();
 b15zdnd11an1n64x5 FILLER_15_1096 ();
 b15zdnd11an1n32x5 FILLER_15_1160 ();
 b15zdnd11an1n16x5 FILLER_15_1192 ();
 b15zdnd00an1n02x5 FILLER_15_1208 ();
 b15zdnd00an1n01x5 FILLER_15_1210 ();
 b15zdnd11an1n08x5 FILLER_15_1227 ();
 b15zdnd11an1n04x5 FILLER_15_1235 ();
 b15zdnd00an1n02x5 FILLER_15_1239 ();
 b15zdnd11an1n64x5 FILLER_15_1257 ();
 b15zdnd11an1n64x5 FILLER_15_1321 ();
 b15zdnd11an1n04x5 FILLER_15_1385 ();
 b15zdnd11an1n08x5 FILLER_15_1397 ();
 b15zdnd00an1n02x5 FILLER_15_1405 ();
 b15zdnd11an1n64x5 FILLER_15_1415 ();
 b15zdnd11an1n04x5 FILLER_15_1479 ();
 b15zdnd00an1n02x5 FILLER_15_1483 ();
 b15zdnd00an1n01x5 FILLER_15_1485 ();
 b15zdnd11an1n16x5 FILLER_15_2257 ();
 b15zdnd11an1n08x5 FILLER_15_2273 ();
 b15zdnd00an1n02x5 FILLER_15_2281 ();
 b15zdnd00an1n01x5 FILLER_15_2283 ();
 b15zdnd11an1n64x5 FILLER_16_8 ();
 b15zdnd11an1n64x5 FILLER_16_72 ();
 b15zdnd11an1n64x5 FILLER_16_136 ();
 b15zdnd11an1n64x5 FILLER_16_200 ();
 b15zdnd11an1n64x5 FILLER_16_264 ();
 b15zdnd11an1n64x5 FILLER_16_328 ();
 b15zdnd11an1n64x5 FILLER_16_392 ();
 b15zdnd11an1n64x5 FILLER_16_456 ();
 b15zdnd11an1n64x5 FILLER_16_520 ();
 b15zdnd11an1n32x5 FILLER_16_584 ();
 b15zdnd11an1n16x5 FILLER_16_616 ();
 b15zdnd00an1n02x5 FILLER_16_632 ();
 b15zdnd00an1n01x5 FILLER_16_634 ();
 b15zdnd11an1n08x5 FILLER_16_638 ();
 b15zdnd00an1n02x5 FILLER_16_646 ();
 b15zdnd11an1n04x5 FILLER_16_651 ();
 b15zdnd11an1n04x5 FILLER_16_658 ();
 b15zdnd11an1n04x5 FILLER_16_665 ();
 b15zdnd00an1n01x5 FILLER_16_669 ();
 b15zdnd11an1n04x5 FILLER_16_673 ();
 b15zdnd00an1n02x5 FILLER_16_677 ();
 b15zdnd11an1n04x5 FILLER_16_682 ();
 b15zdnd00an1n01x5 FILLER_16_686 ();
 b15zdnd11an1n04x5 FILLER_16_690 ();
 b15zdnd11an1n04x5 FILLER_16_697 ();
 b15zdnd00an1n01x5 FILLER_16_701 ();
 b15zdnd11an1n04x5 FILLER_16_705 ();
 b15zdnd00an1n01x5 FILLER_16_709 ();
 b15zdnd11an1n04x5 FILLER_16_713 ();
 b15zdnd00an1n01x5 FILLER_16_717 ();
 b15zdnd11an1n16x5 FILLER_16_726 ();
 b15zdnd00an1n02x5 FILLER_16_742 ();
 b15zdnd00an1n01x5 FILLER_16_744 ();
 b15zdnd11an1n64x5 FILLER_16_749 ();
 b15zdnd11an1n32x5 FILLER_16_813 ();
 b15zdnd11an1n16x5 FILLER_16_845 ();
 b15zdnd11an1n08x5 FILLER_16_861 ();
 b15zdnd11an1n04x5 FILLER_16_869 ();
 b15zdnd00an1n01x5 FILLER_16_873 ();
 b15zdnd11an1n08x5 FILLER_16_878 ();
 b15zdnd11an1n04x5 FILLER_16_886 ();
 b15zdnd11an1n08x5 FILLER_16_898 ();
 b15zdnd11an1n04x5 FILLER_16_906 ();
 b15zdnd00an1n02x5 FILLER_16_910 ();
 b15zdnd00an1n01x5 FILLER_16_912 ();
 b15zdnd11an1n04x5 FILLER_16_917 ();
 b15zdnd11an1n64x5 FILLER_16_925 ();
 b15zdnd11an1n64x5 FILLER_16_989 ();
 b15zdnd11an1n32x5 FILLER_16_1053 ();
 b15zdnd11an1n04x5 FILLER_16_1085 ();
 b15zdnd11an1n64x5 FILLER_16_1093 ();
 b15zdnd11an1n64x5 FILLER_16_1157 ();
 b15zdnd11an1n64x5 FILLER_16_1221 ();
 b15zdnd11an1n64x5 FILLER_16_1285 ();
 b15zdnd11an1n32x5 FILLER_16_1349 ();
 b15zdnd11an1n08x5 FILLER_16_1381 ();
 b15zdnd00an1n02x5 FILLER_16_1389 ();
 b15zdnd11an1n04x5 FILLER_16_1399 ();
 b15zdnd00an1n02x5 FILLER_16_1403 ();
 b15zdnd00an1n01x5 FILLER_16_1405 ();
 b15zdnd11an1n64x5 FILLER_16_1414 ();
 b15zdnd11an1n08x5 FILLER_16_2265 ();
 b15zdnd00an1n02x5 FILLER_16_2273 ();
 b15zdnd00an1n01x5 FILLER_16_2275 ();
 b15zdnd11an1n64x5 FILLER_17_0 ();
 b15zdnd11an1n64x5 FILLER_17_64 ();
 b15zdnd11an1n64x5 FILLER_17_128 ();
 b15zdnd11an1n64x5 FILLER_17_192 ();
 b15zdnd11an1n64x5 FILLER_17_256 ();
 b15zdnd11an1n64x5 FILLER_17_320 ();
 b15zdnd11an1n64x5 FILLER_17_384 ();
 b15zdnd11an1n64x5 FILLER_17_448 ();
 b15zdnd11an1n64x5 FILLER_17_512 ();
 b15zdnd11an1n32x5 FILLER_17_576 ();
 b15zdnd11an1n16x5 FILLER_17_608 ();
 b15zdnd11an1n08x5 FILLER_17_624 ();
 b15zdnd11an1n04x5 FILLER_17_632 ();
 b15zdnd11an1n16x5 FILLER_17_639 ();
 b15zdnd11an1n08x5 FILLER_17_655 ();
 b15zdnd11an1n04x5 FILLER_17_666 ();
 b15zdnd11an1n04x5 FILLER_17_673 ();
 b15zdnd00an1n01x5 FILLER_17_677 ();
 b15zdnd11an1n04x5 FILLER_17_681 ();
 b15zdnd11an1n04x5 FILLER_17_688 ();
 b15zdnd11an1n08x5 FILLER_17_695 ();
 b15zdnd11an1n04x5 FILLER_17_703 ();
 b15zdnd00an1n02x5 FILLER_17_707 ();
 b15zdnd00an1n01x5 FILLER_17_709 ();
 b15zdnd11an1n16x5 FILLER_17_718 ();
 b15zdnd11an1n04x5 FILLER_17_734 ();
 b15zdnd00an1n02x5 FILLER_17_738 ();
 b15zdnd11an1n08x5 FILLER_17_782 ();
 b15zdnd11an1n04x5 FILLER_17_790 ();
 b15zdnd11an1n08x5 FILLER_17_805 ();
 b15zdnd11an1n04x5 FILLER_17_813 ();
 b15zdnd11an1n16x5 FILLER_17_821 ();
 b15zdnd11an1n08x5 FILLER_17_837 ();
 b15zdnd00an1n02x5 FILLER_17_845 ();
 b15zdnd11an1n04x5 FILLER_17_858 ();
 b15zdnd11an1n64x5 FILLER_17_866 ();
 b15zdnd11an1n64x5 FILLER_17_930 ();
 b15zdnd11an1n32x5 FILLER_17_994 ();
 b15zdnd11an1n16x5 FILLER_17_1026 ();
 b15zdnd00an1n01x5 FILLER_17_1042 ();
 b15zdnd11an1n08x5 FILLER_17_1049 ();
 b15zdnd00an1n01x5 FILLER_17_1057 ();
 b15zdnd11an1n04x5 FILLER_17_1066 ();
 b15zdnd11an1n64x5 FILLER_17_1078 ();
 b15zdnd11an1n64x5 FILLER_17_1142 ();
 b15zdnd00an1n01x5 FILLER_17_1206 ();
 b15zdnd11an1n08x5 FILLER_17_1223 ();
 b15zdnd11an1n04x5 FILLER_17_1231 ();
 b15zdnd00an1n02x5 FILLER_17_1235 ();
 b15zdnd00an1n01x5 FILLER_17_1237 ();
 b15zdnd11an1n64x5 FILLER_17_1254 ();
 b15zdnd11an1n64x5 FILLER_17_1318 ();
 b15zdnd11an1n08x5 FILLER_17_1382 ();
 b15zdnd11an1n04x5 FILLER_17_1390 ();
 b15zdnd00an1n02x5 FILLER_17_1394 ();
 b15zdnd00an1n01x5 FILLER_17_1396 ();
 b15zdnd11an1n04x5 FILLER_17_1405 ();
 b15zdnd11an1n64x5 FILLER_17_1419 ();
 b15zdnd00an1n02x5 FILLER_17_1483 ();
 b15zdnd00an1n01x5 FILLER_17_1485 ();
 b15zdnd11an1n16x5 FILLER_17_2257 ();
 b15zdnd11an1n08x5 FILLER_17_2273 ();
 b15zdnd00an1n02x5 FILLER_17_2281 ();
 b15zdnd00an1n01x5 FILLER_17_2283 ();
 b15zdnd11an1n64x5 FILLER_18_8 ();
 b15zdnd11an1n64x5 FILLER_18_72 ();
 b15zdnd11an1n64x5 FILLER_18_136 ();
 b15zdnd11an1n64x5 FILLER_18_200 ();
 b15zdnd11an1n64x5 FILLER_18_264 ();
 b15zdnd11an1n64x5 FILLER_18_328 ();
 b15zdnd11an1n64x5 FILLER_18_392 ();
 b15zdnd11an1n64x5 FILLER_18_456 ();
 b15zdnd11an1n64x5 FILLER_18_520 ();
 b15zdnd11an1n16x5 FILLER_18_584 ();
 b15zdnd11an1n04x5 FILLER_18_600 ();
 b15zdnd00an1n02x5 FILLER_18_604 ();
 b15zdnd11an1n04x5 FILLER_18_623 ();
 b15zdnd00an1n01x5 FILLER_18_627 ();
 b15zdnd11an1n16x5 FILLER_18_645 ();
 b15zdnd11an1n08x5 FILLER_18_661 ();
 b15zdnd11an1n04x5 FILLER_18_669 ();
 b15zdnd00an1n02x5 FILLER_18_673 ();
 b15zdnd00an1n01x5 FILLER_18_675 ();
 b15zdnd11an1n04x5 FILLER_18_679 ();
 b15zdnd00an1n01x5 FILLER_18_683 ();
 b15zdnd11an1n04x5 FILLER_18_687 ();
 b15zdnd11an1n16x5 FILLER_18_694 ();
 b15zdnd11an1n08x5 FILLER_18_710 ();
 b15zdnd11an1n32x5 FILLER_18_726 ();
 b15zdnd11an1n04x5 FILLER_18_758 ();
 b15zdnd00an1n02x5 FILLER_18_762 ();
 b15zdnd00an1n01x5 FILLER_18_764 ();
 b15zdnd11an1n32x5 FILLER_18_807 ();
 b15zdnd11an1n08x5 FILLER_18_839 ();
 b15zdnd00an1n02x5 FILLER_18_847 ();
 b15zdnd11an1n04x5 FILLER_18_857 ();
 b15zdnd11an1n64x5 FILLER_18_877 ();
 b15zdnd11an1n08x5 FILLER_18_941 ();
 b15zdnd00an1n01x5 FILLER_18_949 ();
 b15zdnd11an1n08x5 FILLER_18_958 ();
 b15zdnd11an1n16x5 FILLER_18_974 ();
 b15zdnd00an1n02x5 FILLER_18_990 ();
 b15zdnd00an1n01x5 FILLER_18_992 ();
 b15zdnd11an1n32x5 FILLER_18_1005 ();
 b15zdnd11an1n16x5 FILLER_18_1079 ();
 b15zdnd11an1n04x5 FILLER_18_1095 ();
 b15zdnd11an1n16x5 FILLER_18_1115 ();
 b15zdnd11an1n04x5 FILLER_18_1137 ();
 b15zdnd11an1n16x5 FILLER_18_1149 ();
 b15zdnd11an1n08x5 FILLER_18_1165 ();
 b15zdnd11an1n04x5 FILLER_18_1173 ();
 b15zdnd00an1n01x5 FILLER_18_1177 ();
 b15zdnd11an1n32x5 FILLER_18_1182 ();
 b15zdnd11an1n08x5 FILLER_18_1214 ();
 b15zdnd00an1n02x5 FILLER_18_1222 ();
 b15zdnd00an1n01x5 FILLER_18_1224 ();
 b15zdnd11an1n08x5 FILLER_18_1267 ();
 b15zdnd11an1n04x5 FILLER_18_1275 ();
 b15zdnd00an1n01x5 FILLER_18_1279 ();
 b15zdnd11an1n04x5 FILLER_18_1293 ();
 b15zdnd11an1n32x5 FILLER_18_1307 ();
 b15zdnd11an1n08x5 FILLER_18_1339 ();
 b15zdnd00an1n02x5 FILLER_18_1347 ();
 b15zdnd11an1n64x5 FILLER_18_1365 ();
 b15zdnd11an1n32x5 FILLER_18_1429 ();
 b15zdnd11an1n16x5 FILLER_18_1461 ();
 b15zdnd00an1n01x5 FILLER_18_1477 ();
 b15zdnd11an1n08x5 FILLER_18_2265 ();
 b15zdnd00an1n02x5 FILLER_18_2273 ();
 b15zdnd00an1n01x5 FILLER_18_2275 ();
 b15zdnd11an1n64x5 FILLER_19_0 ();
 b15zdnd11an1n64x5 FILLER_19_64 ();
 b15zdnd11an1n64x5 FILLER_19_128 ();
 b15zdnd11an1n64x5 FILLER_19_192 ();
 b15zdnd11an1n64x5 FILLER_19_256 ();
 b15zdnd11an1n64x5 FILLER_19_320 ();
 b15zdnd11an1n64x5 FILLER_19_384 ();
 b15zdnd11an1n64x5 FILLER_19_448 ();
 b15zdnd11an1n64x5 FILLER_19_512 ();
 b15zdnd11an1n64x5 FILLER_19_576 ();
 b15zdnd11an1n32x5 FILLER_19_640 ();
 b15zdnd11an1n08x5 FILLER_19_672 ();
 b15zdnd00an1n02x5 FILLER_19_680 ();
 b15zdnd11an1n64x5 FILLER_19_685 ();
 b15zdnd11an1n64x5 FILLER_19_749 ();
 b15zdnd11an1n64x5 FILLER_19_813 ();
 b15zdnd11an1n64x5 FILLER_19_877 ();
 b15zdnd11an1n32x5 FILLER_19_941 ();
 b15zdnd00an1n02x5 FILLER_19_973 ();
 b15zdnd11an1n64x5 FILLER_19_991 ();
 b15zdnd11an1n64x5 FILLER_19_1055 ();
 b15zdnd11an1n64x5 FILLER_19_1119 ();
 b15zdnd11an1n32x5 FILLER_19_1183 ();
 b15zdnd11an1n16x5 FILLER_19_1215 ();
 b15zdnd00an1n02x5 FILLER_19_1231 ();
 b15zdnd11an1n64x5 FILLER_19_1239 ();
 b15zdnd11an1n64x5 FILLER_19_1303 ();
 b15zdnd11an1n64x5 FILLER_19_1367 ();
 b15zdnd11an1n32x5 FILLER_19_1431 ();
 b15zdnd11an1n16x5 FILLER_19_1463 ();
 b15zdnd11an1n04x5 FILLER_19_1479 ();
 b15zdnd00an1n02x5 FILLER_19_1483 ();
 b15zdnd00an1n01x5 FILLER_19_1485 ();
 b15zdnd11an1n16x5 FILLER_19_2257 ();
 b15zdnd11an1n08x5 FILLER_19_2273 ();
 b15zdnd00an1n02x5 FILLER_19_2281 ();
 b15zdnd00an1n01x5 FILLER_19_2283 ();
 b15zdnd11an1n64x5 FILLER_20_8 ();
 b15zdnd11an1n64x5 FILLER_20_72 ();
 b15zdnd11an1n64x5 FILLER_20_136 ();
 b15zdnd11an1n64x5 FILLER_20_200 ();
 b15zdnd11an1n64x5 FILLER_20_264 ();
 b15zdnd11an1n64x5 FILLER_20_328 ();
 b15zdnd11an1n64x5 FILLER_20_392 ();
 b15zdnd11an1n64x5 FILLER_20_456 ();
 b15zdnd11an1n64x5 FILLER_20_520 ();
 b15zdnd11an1n64x5 FILLER_20_584 ();
 b15zdnd11an1n64x5 FILLER_20_648 ();
 b15zdnd11an1n04x5 FILLER_20_712 ();
 b15zdnd00an1n02x5 FILLER_20_716 ();
 b15zdnd11an1n64x5 FILLER_20_726 ();
 b15zdnd11an1n64x5 FILLER_20_790 ();
 b15zdnd11an1n64x5 FILLER_20_854 ();
 b15zdnd11an1n32x5 FILLER_20_918 ();
 b15zdnd11an1n16x5 FILLER_20_950 ();
 b15zdnd00an1n02x5 FILLER_20_966 ();
 b15zdnd11an1n16x5 FILLER_20_1010 ();
 b15zdnd11an1n04x5 FILLER_20_1026 ();
 b15zdnd00an1n02x5 FILLER_20_1030 ();
 b15zdnd11an1n64x5 FILLER_20_1074 ();
 b15zdnd11an1n64x5 FILLER_20_1138 ();
 b15zdnd11an1n64x5 FILLER_20_1202 ();
 b15zdnd11an1n64x5 FILLER_20_1266 ();
 b15zdnd11an1n64x5 FILLER_20_1330 ();
 b15zdnd11an1n04x5 FILLER_20_1394 ();
 b15zdnd00an1n02x5 FILLER_20_1398 ();
 b15zdnd00an1n01x5 FILLER_20_1400 ();
 b15zdnd11an1n64x5 FILLER_20_1409 ();
 b15zdnd11an1n04x5 FILLER_20_1473 ();
 b15zdnd00an1n01x5 FILLER_20_1477 ();
 b15zdnd11an1n08x5 FILLER_20_2265 ();
 b15zdnd00an1n02x5 FILLER_20_2273 ();
 b15zdnd00an1n01x5 FILLER_20_2275 ();
 b15zdnd11an1n64x5 FILLER_21_0 ();
 b15zdnd11an1n64x5 FILLER_21_64 ();
 b15zdnd11an1n64x5 FILLER_21_128 ();
 b15zdnd11an1n64x5 FILLER_21_192 ();
 b15zdnd11an1n64x5 FILLER_21_256 ();
 b15zdnd11an1n64x5 FILLER_21_320 ();
 b15zdnd11an1n64x5 FILLER_21_384 ();
 b15zdnd11an1n64x5 FILLER_21_448 ();
 b15zdnd11an1n64x5 FILLER_21_512 ();
 b15zdnd11an1n64x5 FILLER_21_576 ();
 b15zdnd11an1n64x5 FILLER_21_640 ();
 b15zdnd11an1n64x5 FILLER_21_704 ();
 b15zdnd11an1n64x5 FILLER_21_768 ();
 b15zdnd11an1n64x5 FILLER_21_832 ();
 b15zdnd11an1n32x5 FILLER_21_896 ();
 b15zdnd11an1n16x5 FILLER_21_928 ();
 b15zdnd11an1n08x5 FILLER_21_944 ();
 b15zdnd11an1n04x5 FILLER_21_952 ();
 b15zdnd11an1n64x5 FILLER_21_970 ();
 b15zdnd11an1n64x5 FILLER_21_1034 ();
 b15zdnd11an1n64x5 FILLER_21_1098 ();
 b15zdnd11an1n64x5 FILLER_21_1162 ();
 b15zdnd11an1n32x5 FILLER_21_1226 ();
 b15zdnd00an1n01x5 FILLER_21_1258 ();
 b15zdnd11an1n64x5 FILLER_21_1275 ();
 b15zdnd11an1n64x5 FILLER_21_1339 ();
 b15zdnd11an1n64x5 FILLER_21_1403 ();
 b15zdnd11an1n16x5 FILLER_21_1467 ();
 b15zdnd00an1n02x5 FILLER_21_1483 ();
 b15zdnd00an1n01x5 FILLER_21_1485 ();
 b15zdnd11an1n16x5 FILLER_21_2257 ();
 b15zdnd11an1n08x5 FILLER_21_2273 ();
 b15zdnd00an1n02x5 FILLER_21_2281 ();
 b15zdnd00an1n01x5 FILLER_21_2283 ();
 b15zdnd11an1n64x5 FILLER_22_8 ();
 b15zdnd11an1n64x5 FILLER_22_72 ();
 b15zdnd11an1n64x5 FILLER_22_136 ();
 b15zdnd11an1n64x5 FILLER_22_200 ();
 b15zdnd11an1n64x5 FILLER_22_264 ();
 b15zdnd11an1n64x5 FILLER_22_328 ();
 b15zdnd11an1n64x5 FILLER_22_392 ();
 b15zdnd11an1n64x5 FILLER_22_456 ();
 b15zdnd11an1n64x5 FILLER_22_520 ();
 b15zdnd11an1n64x5 FILLER_22_584 ();
 b15zdnd11an1n64x5 FILLER_22_648 ();
 b15zdnd11an1n04x5 FILLER_22_712 ();
 b15zdnd00an1n02x5 FILLER_22_716 ();
 b15zdnd11an1n64x5 FILLER_22_726 ();
 b15zdnd11an1n64x5 FILLER_22_790 ();
 b15zdnd11an1n64x5 FILLER_22_854 ();
 b15zdnd11an1n64x5 FILLER_22_918 ();
 b15zdnd11an1n08x5 FILLER_22_982 ();
 b15zdnd11an1n04x5 FILLER_22_990 ();
 b15zdnd00an1n01x5 FILLER_22_994 ();
 b15zdnd11an1n64x5 FILLER_22_1009 ();
 b15zdnd11an1n64x5 FILLER_22_1073 ();
 b15zdnd11an1n64x5 FILLER_22_1137 ();
 b15zdnd11an1n64x5 FILLER_22_1201 ();
 b15zdnd11an1n64x5 FILLER_22_1265 ();
 b15zdnd11an1n16x5 FILLER_22_1329 ();
 b15zdnd11an1n08x5 FILLER_22_1345 ();
 b15zdnd00an1n02x5 FILLER_22_1353 ();
 b15zdnd11an1n64x5 FILLER_22_1371 ();
 b15zdnd11an1n32x5 FILLER_22_1435 ();
 b15zdnd11an1n08x5 FILLER_22_1467 ();
 b15zdnd00an1n02x5 FILLER_22_1475 ();
 b15zdnd00an1n01x5 FILLER_22_1477 ();
 b15zdnd11an1n08x5 FILLER_22_2265 ();
 b15zdnd00an1n02x5 FILLER_22_2273 ();
 b15zdnd00an1n01x5 FILLER_22_2275 ();
 b15zdnd11an1n64x5 FILLER_23_0 ();
 b15zdnd11an1n64x5 FILLER_23_64 ();
 b15zdnd11an1n64x5 FILLER_23_128 ();
 b15zdnd11an1n64x5 FILLER_23_192 ();
 b15zdnd11an1n64x5 FILLER_23_256 ();
 b15zdnd11an1n64x5 FILLER_23_320 ();
 b15zdnd11an1n64x5 FILLER_23_384 ();
 b15zdnd11an1n64x5 FILLER_23_448 ();
 b15zdnd11an1n64x5 FILLER_23_512 ();
 b15zdnd11an1n64x5 FILLER_23_576 ();
 b15zdnd11an1n64x5 FILLER_23_640 ();
 b15zdnd11an1n64x5 FILLER_23_704 ();
 b15zdnd11an1n64x5 FILLER_23_768 ();
 b15zdnd11an1n64x5 FILLER_23_832 ();
 b15zdnd11an1n64x5 FILLER_23_896 ();
 b15zdnd11an1n64x5 FILLER_23_960 ();
 b15zdnd11an1n64x5 FILLER_23_1024 ();
 b15zdnd11an1n64x5 FILLER_23_1088 ();
 b15zdnd11an1n64x5 FILLER_23_1152 ();
 b15zdnd11an1n64x5 FILLER_23_1216 ();
 b15zdnd11an1n64x5 FILLER_23_1280 ();
 b15zdnd11an1n64x5 FILLER_23_1344 ();
 b15zdnd11an1n64x5 FILLER_23_1408 ();
 b15zdnd11an1n08x5 FILLER_23_1472 ();
 b15zdnd11an1n04x5 FILLER_23_1480 ();
 b15zdnd00an1n02x5 FILLER_23_1484 ();
 b15zdnd11an1n16x5 FILLER_23_2257 ();
 b15zdnd11an1n08x5 FILLER_23_2273 ();
 b15zdnd00an1n02x5 FILLER_23_2281 ();
 b15zdnd00an1n01x5 FILLER_23_2283 ();
 b15zdnd11an1n64x5 FILLER_24_8 ();
 b15zdnd11an1n64x5 FILLER_24_72 ();
 b15zdnd11an1n64x5 FILLER_24_136 ();
 b15zdnd11an1n64x5 FILLER_24_200 ();
 b15zdnd11an1n64x5 FILLER_24_264 ();
 b15zdnd11an1n64x5 FILLER_24_328 ();
 b15zdnd11an1n64x5 FILLER_24_392 ();
 b15zdnd11an1n64x5 FILLER_24_456 ();
 b15zdnd11an1n64x5 FILLER_24_520 ();
 b15zdnd11an1n16x5 FILLER_24_584 ();
 b15zdnd11an1n64x5 FILLER_24_642 ();
 b15zdnd11an1n08x5 FILLER_24_706 ();
 b15zdnd11an1n04x5 FILLER_24_714 ();
 b15zdnd11an1n64x5 FILLER_24_726 ();
 b15zdnd11an1n64x5 FILLER_24_790 ();
 b15zdnd11an1n32x5 FILLER_24_854 ();
 b15zdnd11an1n16x5 FILLER_24_886 ();
 b15zdnd11an1n64x5 FILLER_24_918 ();
 b15zdnd11an1n64x5 FILLER_24_982 ();
 b15zdnd11an1n64x5 FILLER_24_1046 ();
 b15zdnd11an1n64x5 FILLER_24_1110 ();
 b15zdnd11an1n64x5 FILLER_24_1174 ();
 b15zdnd11an1n64x5 FILLER_24_1238 ();
 b15zdnd11an1n64x5 FILLER_24_1302 ();
 b15zdnd11an1n64x5 FILLER_24_1366 ();
 b15zdnd11an1n32x5 FILLER_24_1430 ();
 b15zdnd11an1n16x5 FILLER_24_1462 ();
 b15zdnd11an1n08x5 FILLER_24_2265 ();
 b15zdnd00an1n02x5 FILLER_24_2273 ();
 b15zdnd00an1n01x5 FILLER_24_2275 ();
 b15zdnd11an1n64x5 FILLER_25_0 ();
 b15zdnd11an1n64x5 FILLER_25_64 ();
 b15zdnd11an1n64x5 FILLER_25_128 ();
 b15zdnd11an1n64x5 FILLER_25_192 ();
 b15zdnd11an1n64x5 FILLER_25_256 ();
 b15zdnd11an1n64x5 FILLER_25_320 ();
 b15zdnd11an1n64x5 FILLER_25_384 ();
 b15zdnd11an1n64x5 FILLER_25_448 ();
 b15zdnd11an1n64x5 FILLER_25_512 ();
 b15zdnd11an1n32x5 FILLER_25_576 ();
 b15zdnd11an1n08x5 FILLER_25_608 ();
 b15zdnd11an1n04x5 FILLER_25_616 ();
 b15zdnd00an1n01x5 FILLER_25_620 ();
 b15zdnd11an1n64x5 FILLER_25_663 ();
 b15zdnd11an1n64x5 FILLER_25_727 ();
 b15zdnd11an1n64x5 FILLER_25_791 ();
 b15zdnd11an1n64x5 FILLER_25_855 ();
 b15zdnd11an1n64x5 FILLER_25_919 ();
 b15zdnd11an1n64x5 FILLER_25_983 ();
 b15zdnd11an1n64x5 FILLER_25_1047 ();
 b15zdnd11an1n64x5 FILLER_25_1111 ();
 b15zdnd11an1n64x5 FILLER_25_1175 ();
 b15zdnd11an1n64x5 FILLER_25_1239 ();
 b15zdnd11an1n64x5 FILLER_25_1303 ();
 b15zdnd11an1n64x5 FILLER_25_1367 ();
 b15zdnd11an1n32x5 FILLER_25_1431 ();
 b15zdnd11an1n16x5 FILLER_25_1463 ();
 b15zdnd11an1n04x5 FILLER_25_1479 ();
 b15zdnd00an1n02x5 FILLER_25_1483 ();
 b15zdnd00an1n01x5 FILLER_25_1485 ();
 b15zdnd11an1n16x5 FILLER_25_2257 ();
 b15zdnd11an1n08x5 FILLER_25_2273 ();
 b15zdnd00an1n02x5 FILLER_25_2281 ();
 b15zdnd00an1n01x5 FILLER_25_2283 ();
 b15zdnd11an1n64x5 FILLER_26_8 ();
 b15zdnd11an1n64x5 FILLER_26_72 ();
 b15zdnd11an1n64x5 FILLER_26_136 ();
 b15zdnd11an1n64x5 FILLER_26_200 ();
 b15zdnd11an1n64x5 FILLER_26_264 ();
 b15zdnd11an1n64x5 FILLER_26_328 ();
 b15zdnd11an1n64x5 FILLER_26_392 ();
 b15zdnd11an1n64x5 FILLER_26_456 ();
 b15zdnd11an1n64x5 FILLER_26_520 ();
 b15zdnd11an1n16x5 FILLER_26_584 ();
 b15zdnd11an1n04x5 FILLER_26_600 ();
 b15zdnd00an1n01x5 FILLER_26_604 ();
 b15zdnd11an1n08x5 FILLER_26_647 ();
 b15zdnd11an1n04x5 FILLER_26_655 ();
 b15zdnd11an1n16x5 FILLER_26_701 ();
 b15zdnd00an1n01x5 FILLER_26_717 ();
 b15zdnd11an1n64x5 FILLER_26_726 ();
 b15zdnd11an1n64x5 FILLER_26_790 ();
 b15zdnd11an1n64x5 FILLER_26_854 ();
 b15zdnd11an1n64x5 FILLER_26_918 ();
 b15zdnd11an1n64x5 FILLER_26_982 ();
 b15zdnd11an1n32x5 FILLER_26_1046 ();
 b15zdnd11an1n08x5 FILLER_26_1078 ();
 b15zdnd11an1n04x5 FILLER_26_1086 ();
 b15zdnd00an1n02x5 FILLER_26_1090 ();
 b15zdnd11an1n64x5 FILLER_26_1134 ();
 b15zdnd11an1n64x5 FILLER_26_1198 ();
 b15zdnd11an1n64x5 FILLER_26_1262 ();
 b15zdnd11an1n64x5 FILLER_26_1326 ();
 b15zdnd11an1n64x5 FILLER_26_1390 ();
 b15zdnd11an1n16x5 FILLER_26_1454 ();
 b15zdnd11an1n08x5 FILLER_26_1470 ();
 b15zdnd11an1n08x5 FILLER_26_2265 ();
 b15zdnd00an1n02x5 FILLER_26_2273 ();
 b15zdnd00an1n01x5 FILLER_26_2275 ();
 b15zdnd11an1n64x5 FILLER_27_0 ();
 b15zdnd11an1n64x5 FILLER_27_64 ();
 b15zdnd11an1n64x5 FILLER_27_128 ();
 b15zdnd11an1n64x5 FILLER_27_192 ();
 b15zdnd11an1n64x5 FILLER_27_256 ();
 b15zdnd11an1n64x5 FILLER_27_320 ();
 b15zdnd11an1n64x5 FILLER_27_384 ();
 b15zdnd11an1n64x5 FILLER_27_448 ();
 b15zdnd11an1n64x5 FILLER_27_512 ();
 b15zdnd11an1n64x5 FILLER_27_576 ();
 b15zdnd11an1n16x5 FILLER_27_640 ();
 b15zdnd00an1n01x5 FILLER_27_656 ();
 b15zdnd11an1n64x5 FILLER_27_699 ();
 b15zdnd11an1n64x5 FILLER_27_763 ();
 b15zdnd11an1n64x5 FILLER_27_827 ();
 b15zdnd11an1n64x5 FILLER_27_891 ();
 b15zdnd11an1n64x5 FILLER_27_955 ();
 b15zdnd11an1n64x5 FILLER_27_1019 ();
 b15zdnd11an1n32x5 FILLER_27_1083 ();
 b15zdnd11an1n16x5 FILLER_27_1115 ();
 b15zdnd00an1n02x5 FILLER_27_1131 ();
 b15zdnd00an1n01x5 FILLER_27_1133 ();
 b15zdnd11an1n64x5 FILLER_27_1176 ();
 b15zdnd11an1n64x5 FILLER_27_1240 ();
 b15zdnd11an1n64x5 FILLER_27_1304 ();
 b15zdnd11an1n64x5 FILLER_27_1368 ();
 b15zdnd11an1n32x5 FILLER_27_1432 ();
 b15zdnd11an1n16x5 FILLER_27_1464 ();
 b15zdnd11an1n04x5 FILLER_27_1480 ();
 b15zdnd00an1n02x5 FILLER_27_1484 ();
 b15zdnd11an1n16x5 FILLER_27_2257 ();
 b15zdnd11an1n08x5 FILLER_27_2273 ();
 b15zdnd00an1n02x5 FILLER_27_2281 ();
 b15zdnd00an1n01x5 FILLER_27_2283 ();
 b15zdnd11an1n64x5 FILLER_28_8 ();
 b15zdnd11an1n64x5 FILLER_28_72 ();
 b15zdnd11an1n64x5 FILLER_28_136 ();
 b15zdnd11an1n64x5 FILLER_28_200 ();
 b15zdnd11an1n64x5 FILLER_28_264 ();
 b15zdnd11an1n64x5 FILLER_28_328 ();
 b15zdnd11an1n64x5 FILLER_28_392 ();
 b15zdnd11an1n64x5 FILLER_28_456 ();
 b15zdnd11an1n64x5 FILLER_28_520 ();
 b15zdnd11an1n64x5 FILLER_28_584 ();
 b15zdnd11an1n64x5 FILLER_28_648 ();
 b15zdnd11an1n04x5 FILLER_28_712 ();
 b15zdnd00an1n02x5 FILLER_28_716 ();
 b15zdnd11an1n64x5 FILLER_28_726 ();
 b15zdnd11an1n64x5 FILLER_28_790 ();
 b15zdnd11an1n04x5 FILLER_28_854 ();
 b15zdnd00an1n02x5 FILLER_28_858 ();
 b15zdnd00an1n01x5 FILLER_28_860 ();
 b15zdnd11an1n64x5 FILLER_28_903 ();
 b15zdnd11an1n64x5 FILLER_28_967 ();
 b15zdnd11an1n64x5 FILLER_28_1031 ();
 b15zdnd11an1n64x5 FILLER_28_1095 ();
 b15zdnd11an1n64x5 FILLER_28_1159 ();
 b15zdnd11an1n64x5 FILLER_28_1223 ();
 b15zdnd11an1n64x5 FILLER_28_1287 ();
 b15zdnd11an1n64x5 FILLER_28_1351 ();
 b15zdnd11an1n32x5 FILLER_28_1415 ();
 b15zdnd11an1n16x5 FILLER_28_1447 ();
 b15zdnd11an1n08x5 FILLER_28_1463 ();
 b15zdnd11an1n04x5 FILLER_28_1471 ();
 b15zdnd00an1n02x5 FILLER_28_1475 ();
 b15zdnd00an1n01x5 FILLER_28_1477 ();
 b15zdnd11an1n08x5 FILLER_28_2265 ();
 b15zdnd00an1n02x5 FILLER_28_2273 ();
 b15zdnd00an1n01x5 FILLER_28_2275 ();
 b15zdnd11an1n64x5 FILLER_29_0 ();
 b15zdnd11an1n64x5 FILLER_29_64 ();
 b15zdnd11an1n64x5 FILLER_29_128 ();
 b15zdnd11an1n64x5 FILLER_29_192 ();
 b15zdnd11an1n64x5 FILLER_29_256 ();
 b15zdnd11an1n64x5 FILLER_29_320 ();
 b15zdnd11an1n64x5 FILLER_29_384 ();
 b15zdnd11an1n64x5 FILLER_29_448 ();
 b15zdnd11an1n64x5 FILLER_29_512 ();
 b15zdnd11an1n64x5 FILLER_29_576 ();
 b15zdnd11an1n64x5 FILLER_29_640 ();
 b15zdnd11an1n64x5 FILLER_29_704 ();
 b15zdnd11an1n32x5 FILLER_29_768 ();
 b15zdnd11an1n08x5 FILLER_29_800 ();
 b15zdnd00an1n02x5 FILLER_29_808 ();
 b15zdnd11an1n32x5 FILLER_29_852 ();
 b15zdnd11an1n08x5 FILLER_29_884 ();
 b15zdnd11an1n04x5 FILLER_29_892 ();
 b15zdnd00an1n02x5 FILLER_29_896 ();
 b15zdnd00an1n01x5 FILLER_29_898 ();
 b15zdnd11an1n64x5 FILLER_29_941 ();
 b15zdnd11an1n32x5 FILLER_29_1005 ();
 b15zdnd11an1n64x5 FILLER_29_1079 ();
 b15zdnd11an1n64x5 FILLER_29_1143 ();
 b15zdnd11an1n16x5 FILLER_29_1207 ();
 b15zdnd11an1n08x5 FILLER_29_1223 ();
 b15zdnd11an1n04x5 FILLER_29_1231 ();
 b15zdnd00an1n01x5 FILLER_29_1235 ();
 b15zdnd11an1n64x5 FILLER_29_1278 ();
 b15zdnd11an1n64x5 FILLER_29_1342 ();
 b15zdnd11an1n64x5 FILLER_29_1406 ();
 b15zdnd11an1n16x5 FILLER_29_1470 ();
 b15zdnd11an1n16x5 FILLER_29_2257 ();
 b15zdnd11an1n08x5 FILLER_29_2273 ();
 b15zdnd00an1n02x5 FILLER_29_2281 ();
 b15zdnd00an1n01x5 FILLER_29_2283 ();
 b15zdnd11an1n64x5 FILLER_30_8 ();
 b15zdnd11an1n64x5 FILLER_30_72 ();
 b15zdnd11an1n64x5 FILLER_30_136 ();
 b15zdnd11an1n64x5 FILLER_30_200 ();
 b15zdnd11an1n64x5 FILLER_30_264 ();
 b15zdnd11an1n64x5 FILLER_30_328 ();
 b15zdnd11an1n64x5 FILLER_30_392 ();
 b15zdnd11an1n64x5 FILLER_30_456 ();
 b15zdnd11an1n64x5 FILLER_30_520 ();
 b15zdnd11an1n64x5 FILLER_30_584 ();
 b15zdnd11an1n64x5 FILLER_30_648 ();
 b15zdnd11an1n04x5 FILLER_30_712 ();
 b15zdnd00an1n02x5 FILLER_30_716 ();
 b15zdnd11an1n64x5 FILLER_30_726 ();
 b15zdnd11an1n64x5 FILLER_30_790 ();
 b15zdnd11an1n64x5 FILLER_30_854 ();
 b15zdnd11an1n64x5 FILLER_30_918 ();
 b15zdnd11an1n64x5 FILLER_30_982 ();
 b15zdnd11an1n16x5 FILLER_30_1046 ();
 b15zdnd00an1n01x5 FILLER_30_1062 ();
 b15zdnd11an1n64x5 FILLER_30_1105 ();
 b15zdnd11an1n64x5 FILLER_30_1169 ();
 b15zdnd11an1n64x5 FILLER_30_1233 ();
 b15zdnd11an1n64x5 FILLER_30_1297 ();
 b15zdnd11an1n64x5 FILLER_30_1361 ();
 b15zdnd11an1n32x5 FILLER_30_1425 ();
 b15zdnd11an1n16x5 FILLER_30_1457 ();
 b15zdnd11an1n04x5 FILLER_30_1473 ();
 b15zdnd00an1n01x5 FILLER_30_1477 ();
 b15zdnd11an1n08x5 FILLER_30_2265 ();
 b15zdnd00an1n02x5 FILLER_30_2273 ();
 b15zdnd00an1n01x5 FILLER_30_2275 ();
 b15zdnd11an1n64x5 FILLER_31_0 ();
 b15zdnd11an1n64x5 FILLER_31_64 ();
 b15zdnd11an1n64x5 FILLER_31_128 ();
 b15zdnd11an1n64x5 FILLER_31_192 ();
 b15zdnd11an1n64x5 FILLER_31_256 ();
 b15zdnd11an1n64x5 FILLER_31_320 ();
 b15zdnd11an1n64x5 FILLER_31_384 ();
 b15zdnd11an1n64x5 FILLER_31_448 ();
 b15zdnd11an1n64x5 FILLER_31_512 ();
 b15zdnd11an1n64x5 FILLER_31_576 ();
 b15zdnd11an1n64x5 FILLER_31_640 ();
 b15zdnd11an1n64x5 FILLER_31_704 ();
 b15zdnd11an1n32x5 FILLER_31_768 ();
 b15zdnd00an1n02x5 FILLER_31_800 ();
 b15zdnd11an1n64x5 FILLER_31_844 ();
 b15zdnd11an1n64x5 FILLER_31_908 ();
 b15zdnd11an1n64x5 FILLER_31_972 ();
 b15zdnd11an1n64x5 FILLER_31_1036 ();
 b15zdnd11an1n64x5 FILLER_31_1100 ();
 b15zdnd11an1n64x5 FILLER_31_1164 ();
 b15zdnd11an1n64x5 FILLER_31_1228 ();
 b15zdnd11an1n64x5 FILLER_31_1292 ();
 b15zdnd11an1n64x5 FILLER_31_1356 ();
 b15zdnd11an1n64x5 FILLER_31_1420 ();
 b15zdnd00an1n02x5 FILLER_31_1484 ();
 b15zdnd11an1n16x5 FILLER_31_2257 ();
 b15zdnd11an1n08x5 FILLER_31_2273 ();
 b15zdnd00an1n02x5 FILLER_31_2281 ();
 b15zdnd00an1n01x5 FILLER_31_2283 ();
 b15zdnd11an1n64x5 FILLER_32_8 ();
 b15zdnd11an1n64x5 FILLER_32_72 ();
 b15zdnd11an1n64x5 FILLER_32_136 ();
 b15zdnd11an1n64x5 FILLER_32_200 ();
 b15zdnd11an1n64x5 FILLER_32_264 ();
 b15zdnd11an1n64x5 FILLER_32_328 ();
 b15zdnd11an1n64x5 FILLER_32_392 ();
 b15zdnd11an1n64x5 FILLER_32_456 ();
 b15zdnd11an1n64x5 FILLER_32_520 ();
 b15zdnd11an1n64x5 FILLER_32_584 ();
 b15zdnd11an1n64x5 FILLER_32_648 ();
 b15zdnd11an1n04x5 FILLER_32_712 ();
 b15zdnd00an1n02x5 FILLER_32_716 ();
 b15zdnd11an1n16x5 FILLER_32_726 ();
 b15zdnd11an1n04x5 FILLER_32_742 ();
 b15zdnd00an1n02x5 FILLER_32_746 ();
 b15zdnd00an1n01x5 FILLER_32_748 ();
 b15zdnd11an1n16x5 FILLER_32_791 ();
 b15zdnd11an1n04x5 FILLER_32_807 ();
 b15zdnd11an1n64x5 FILLER_32_853 ();
 b15zdnd11an1n64x5 FILLER_32_917 ();
 b15zdnd11an1n32x5 FILLER_32_981 ();
 b15zdnd11an1n16x5 FILLER_32_1013 ();
 b15zdnd11an1n08x5 FILLER_32_1029 ();
 b15zdnd11an1n04x5 FILLER_32_1037 ();
 b15zdnd11an1n64x5 FILLER_32_1058 ();
 b15zdnd11an1n08x5 FILLER_32_1122 ();
 b15zdnd00an1n02x5 FILLER_32_1130 ();
 b15zdnd00an1n01x5 FILLER_32_1132 ();
 b15zdnd11an1n64x5 FILLER_32_1175 ();
 b15zdnd11an1n32x5 FILLER_32_1239 ();
 b15zdnd11an1n08x5 FILLER_32_1271 ();
 b15zdnd11an1n04x5 FILLER_32_1279 ();
 b15zdnd11an1n64x5 FILLER_32_1293 ();
 b15zdnd11an1n64x5 FILLER_32_1357 ();
 b15zdnd11an1n32x5 FILLER_32_1421 ();
 b15zdnd11an1n16x5 FILLER_32_1453 ();
 b15zdnd11an1n08x5 FILLER_32_1469 ();
 b15zdnd00an1n01x5 FILLER_32_1477 ();
 b15zdnd11an1n08x5 FILLER_32_2265 ();
 b15zdnd00an1n02x5 FILLER_32_2273 ();
 b15zdnd00an1n01x5 FILLER_32_2275 ();
 b15zdnd11an1n64x5 FILLER_33_0 ();
 b15zdnd11an1n64x5 FILLER_33_64 ();
 b15zdnd11an1n64x5 FILLER_33_128 ();
 b15zdnd11an1n64x5 FILLER_33_192 ();
 b15zdnd11an1n64x5 FILLER_33_256 ();
 b15zdnd11an1n64x5 FILLER_33_320 ();
 b15zdnd11an1n64x5 FILLER_33_384 ();
 b15zdnd11an1n64x5 FILLER_33_448 ();
 b15zdnd11an1n64x5 FILLER_33_512 ();
 b15zdnd11an1n64x5 FILLER_33_576 ();
 b15zdnd11an1n64x5 FILLER_33_640 ();
 b15zdnd11an1n32x5 FILLER_33_704 ();
 b15zdnd11an1n08x5 FILLER_33_736 ();
 b15zdnd11an1n04x5 FILLER_33_744 ();
 b15zdnd00an1n02x5 FILLER_33_748 ();
 b15zdnd00an1n01x5 FILLER_33_750 ();
 b15zdnd11an1n64x5 FILLER_33_793 ();
 b15zdnd11an1n64x5 FILLER_33_857 ();
 b15zdnd11an1n64x5 FILLER_33_921 ();
 b15zdnd11an1n64x5 FILLER_33_985 ();
 b15zdnd11an1n64x5 FILLER_33_1049 ();
 b15zdnd11an1n64x5 FILLER_33_1113 ();
 b15zdnd11an1n64x5 FILLER_33_1177 ();
 b15zdnd11an1n64x5 FILLER_33_1241 ();
 b15zdnd11an1n64x5 FILLER_33_1305 ();
 b15zdnd11an1n64x5 FILLER_33_1369 ();
 b15zdnd11an1n32x5 FILLER_33_1433 ();
 b15zdnd11an1n16x5 FILLER_33_1465 ();
 b15zdnd11an1n04x5 FILLER_33_1481 ();
 b15zdnd00an1n01x5 FILLER_33_1485 ();
 b15zdnd11an1n16x5 FILLER_33_2257 ();
 b15zdnd11an1n08x5 FILLER_33_2273 ();
 b15zdnd00an1n02x5 FILLER_33_2281 ();
 b15zdnd00an1n01x5 FILLER_33_2283 ();
 b15zdnd11an1n64x5 FILLER_34_8 ();
 b15zdnd11an1n64x5 FILLER_34_72 ();
 b15zdnd11an1n64x5 FILLER_34_136 ();
 b15zdnd11an1n64x5 FILLER_34_200 ();
 b15zdnd11an1n64x5 FILLER_34_264 ();
 b15zdnd11an1n64x5 FILLER_34_328 ();
 b15zdnd11an1n64x5 FILLER_34_392 ();
 b15zdnd11an1n64x5 FILLER_34_456 ();
 b15zdnd11an1n64x5 FILLER_34_520 ();
 b15zdnd11an1n64x5 FILLER_34_584 ();
 b15zdnd11an1n64x5 FILLER_34_648 ();
 b15zdnd11an1n04x5 FILLER_34_712 ();
 b15zdnd00an1n02x5 FILLER_34_716 ();
 b15zdnd00an1n02x5 FILLER_34_726 ();
 b15zdnd11an1n64x5 FILLER_34_770 ();
 b15zdnd11an1n64x5 FILLER_34_834 ();
 b15zdnd11an1n64x5 FILLER_34_898 ();
 b15zdnd11an1n64x5 FILLER_34_962 ();
 b15zdnd11an1n64x5 FILLER_34_1026 ();
 b15zdnd11an1n64x5 FILLER_34_1090 ();
 b15zdnd11an1n32x5 FILLER_34_1154 ();
 b15zdnd11an1n16x5 FILLER_34_1186 ();
 b15zdnd11an1n08x5 FILLER_34_1202 ();
 b15zdnd11an1n04x5 FILLER_34_1210 ();
 b15zdnd00an1n01x5 FILLER_34_1214 ();
 b15zdnd11an1n64x5 FILLER_34_1221 ();
 b15zdnd11an1n64x5 FILLER_34_1285 ();
 b15zdnd11an1n64x5 FILLER_34_1349 ();
 b15zdnd11an1n64x5 FILLER_34_1413 ();
 b15zdnd00an1n01x5 FILLER_34_1477 ();
 b15zdnd11an1n08x5 FILLER_34_2265 ();
 b15zdnd00an1n02x5 FILLER_34_2273 ();
 b15zdnd00an1n01x5 FILLER_34_2275 ();
 b15zdnd11an1n64x5 FILLER_35_0 ();
 b15zdnd11an1n64x5 FILLER_35_64 ();
 b15zdnd11an1n64x5 FILLER_35_128 ();
 b15zdnd11an1n64x5 FILLER_35_192 ();
 b15zdnd11an1n64x5 FILLER_35_256 ();
 b15zdnd11an1n64x5 FILLER_35_320 ();
 b15zdnd11an1n64x5 FILLER_35_384 ();
 b15zdnd11an1n64x5 FILLER_35_448 ();
 b15zdnd11an1n64x5 FILLER_35_512 ();
 b15zdnd11an1n64x5 FILLER_35_576 ();
 b15zdnd11an1n64x5 FILLER_35_640 ();
 b15zdnd11an1n64x5 FILLER_35_704 ();
 b15zdnd11an1n64x5 FILLER_35_768 ();
 b15zdnd11an1n64x5 FILLER_35_832 ();
 b15zdnd11an1n64x5 FILLER_35_896 ();
 b15zdnd11an1n64x5 FILLER_35_960 ();
 b15zdnd11an1n64x5 FILLER_35_1024 ();
 b15zdnd11an1n64x5 FILLER_35_1088 ();
 b15zdnd11an1n64x5 FILLER_35_1152 ();
 b15zdnd11an1n64x5 FILLER_35_1216 ();
 b15zdnd11an1n64x5 FILLER_35_1280 ();
 b15zdnd11an1n64x5 FILLER_35_1344 ();
 b15zdnd11an1n64x5 FILLER_35_1408 ();
 b15zdnd11an1n08x5 FILLER_35_1472 ();
 b15zdnd11an1n04x5 FILLER_35_1480 ();
 b15zdnd00an1n02x5 FILLER_35_1484 ();
 b15zdnd11an1n16x5 FILLER_35_2257 ();
 b15zdnd11an1n08x5 FILLER_35_2273 ();
 b15zdnd00an1n02x5 FILLER_35_2281 ();
 b15zdnd00an1n01x5 FILLER_35_2283 ();
 b15zdnd11an1n64x5 FILLER_36_8 ();
 b15zdnd11an1n64x5 FILLER_36_72 ();
 b15zdnd11an1n64x5 FILLER_36_136 ();
 b15zdnd11an1n64x5 FILLER_36_200 ();
 b15zdnd11an1n64x5 FILLER_36_264 ();
 b15zdnd11an1n64x5 FILLER_36_328 ();
 b15zdnd11an1n64x5 FILLER_36_392 ();
 b15zdnd11an1n64x5 FILLER_36_456 ();
 b15zdnd11an1n64x5 FILLER_36_520 ();
 b15zdnd11an1n64x5 FILLER_36_584 ();
 b15zdnd11an1n16x5 FILLER_36_648 ();
 b15zdnd11an1n08x5 FILLER_36_706 ();
 b15zdnd11an1n04x5 FILLER_36_714 ();
 b15zdnd11an1n64x5 FILLER_36_726 ();
 b15zdnd11an1n64x5 FILLER_36_790 ();
 b15zdnd11an1n64x5 FILLER_36_854 ();
 b15zdnd11an1n64x5 FILLER_36_918 ();
 b15zdnd11an1n64x5 FILLER_36_982 ();
 b15zdnd11an1n32x5 FILLER_36_1046 ();
 b15zdnd00an1n02x5 FILLER_36_1078 ();
 b15zdnd00an1n01x5 FILLER_36_1080 ();
 b15zdnd11an1n64x5 FILLER_36_1095 ();
 b15zdnd11an1n64x5 FILLER_36_1159 ();
 b15zdnd11an1n64x5 FILLER_36_1223 ();
 b15zdnd11an1n32x5 FILLER_36_1287 ();
 b15zdnd11an1n08x5 FILLER_36_1319 ();
 b15zdnd11an1n04x5 FILLER_36_1327 ();
 b15zdnd00an1n02x5 FILLER_36_1331 ();
 b15zdnd00an1n01x5 FILLER_36_1333 ();
 b15zdnd11an1n64x5 FILLER_36_1350 ();
 b15zdnd11an1n64x5 FILLER_36_1414 ();
 b15zdnd11an1n08x5 FILLER_36_2265 ();
 b15zdnd00an1n02x5 FILLER_36_2273 ();
 b15zdnd00an1n01x5 FILLER_36_2275 ();
 b15zdnd11an1n64x5 FILLER_37_0 ();
 b15zdnd11an1n64x5 FILLER_37_64 ();
 b15zdnd11an1n64x5 FILLER_37_128 ();
 b15zdnd11an1n64x5 FILLER_37_192 ();
 b15zdnd11an1n64x5 FILLER_37_256 ();
 b15zdnd11an1n64x5 FILLER_37_320 ();
 b15zdnd11an1n64x5 FILLER_37_384 ();
 b15zdnd11an1n64x5 FILLER_37_448 ();
 b15zdnd11an1n64x5 FILLER_37_512 ();
 b15zdnd11an1n64x5 FILLER_37_576 ();
 b15zdnd11an1n64x5 FILLER_37_640 ();
 b15zdnd11an1n64x5 FILLER_37_704 ();
 b15zdnd11an1n64x5 FILLER_37_768 ();
 b15zdnd11an1n64x5 FILLER_37_832 ();
 b15zdnd11an1n64x5 FILLER_37_896 ();
 b15zdnd11an1n64x5 FILLER_37_960 ();
 b15zdnd11an1n64x5 FILLER_37_1024 ();
 b15zdnd11an1n64x5 FILLER_37_1088 ();
 b15zdnd11an1n64x5 FILLER_37_1152 ();
 b15zdnd11an1n08x5 FILLER_37_1216 ();
 b15zdnd11an1n04x5 FILLER_37_1224 ();
 b15zdnd00an1n02x5 FILLER_37_1228 ();
 b15zdnd11an1n64x5 FILLER_37_1244 ();
 b15zdnd11an1n64x5 FILLER_37_1308 ();
 b15zdnd11an1n64x5 FILLER_37_1372 ();
 b15zdnd11an1n32x5 FILLER_37_1436 ();
 b15zdnd11an1n16x5 FILLER_37_1468 ();
 b15zdnd00an1n02x5 FILLER_37_1484 ();
 b15zdnd11an1n16x5 FILLER_37_2257 ();
 b15zdnd11an1n08x5 FILLER_37_2273 ();
 b15zdnd00an1n02x5 FILLER_37_2281 ();
 b15zdnd00an1n01x5 FILLER_37_2283 ();
 b15zdnd11an1n64x5 FILLER_38_8 ();
 b15zdnd11an1n64x5 FILLER_38_72 ();
 b15zdnd11an1n64x5 FILLER_38_136 ();
 b15zdnd11an1n64x5 FILLER_38_200 ();
 b15zdnd11an1n64x5 FILLER_38_264 ();
 b15zdnd11an1n64x5 FILLER_38_328 ();
 b15zdnd11an1n64x5 FILLER_38_392 ();
 b15zdnd11an1n64x5 FILLER_38_456 ();
 b15zdnd11an1n64x5 FILLER_38_520 ();
 b15zdnd11an1n64x5 FILLER_38_584 ();
 b15zdnd11an1n64x5 FILLER_38_648 ();
 b15zdnd11an1n04x5 FILLER_38_712 ();
 b15zdnd00an1n02x5 FILLER_38_716 ();
 b15zdnd11an1n64x5 FILLER_38_726 ();
 b15zdnd11an1n64x5 FILLER_38_790 ();
 b15zdnd11an1n64x5 FILLER_38_854 ();
 b15zdnd11an1n64x5 FILLER_38_918 ();
 b15zdnd11an1n64x5 FILLER_38_982 ();
 b15zdnd11an1n64x5 FILLER_38_1046 ();
 b15zdnd11an1n64x5 FILLER_38_1110 ();
 b15zdnd11an1n64x5 FILLER_38_1174 ();
 b15zdnd11an1n32x5 FILLER_38_1238 ();
 b15zdnd11an1n16x5 FILLER_38_1270 ();
 b15zdnd00an1n02x5 FILLER_38_1286 ();
 b15zdnd11an1n32x5 FILLER_38_1304 ();
 b15zdnd11an1n64x5 FILLER_38_1346 ();
 b15zdnd11an1n64x5 FILLER_38_1410 ();
 b15zdnd11an1n04x5 FILLER_38_1474 ();
 b15zdnd11an1n08x5 FILLER_38_2265 ();
 b15zdnd00an1n02x5 FILLER_38_2273 ();
 b15zdnd00an1n01x5 FILLER_38_2275 ();
 b15zdnd11an1n64x5 FILLER_39_0 ();
 b15zdnd11an1n64x5 FILLER_39_64 ();
 b15zdnd11an1n64x5 FILLER_39_128 ();
 b15zdnd11an1n64x5 FILLER_39_192 ();
 b15zdnd11an1n64x5 FILLER_39_256 ();
 b15zdnd11an1n64x5 FILLER_39_320 ();
 b15zdnd11an1n64x5 FILLER_39_384 ();
 b15zdnd11an1n64x5 FILLER_39_448 ();
 b15zdnd11an1n64x5 FILLER_39_512 ();
 b15zdnd11an1n64x5 FILLER_39_576 ();
 b15zdnd11an1n64x5 FILLER_39_640 ();
 b15zdnd11an1n64x5 FILLER_39_704 ();
 b15zdnd11an1n64x5 FILLER_39_768 ();
 b15zdnd00an1n02x5 FILLER_39_832 ();
 b15zdnd00an1n01x5 FILLER_39_834 ();
 b15zdnd11an1n64x5 FILLER_39_852 ();
 b15zdnd11an1n64x5 FILLER_39_916 ();
 b15zdnd11an1n64x5 FILLER_39_980 ();
 b15zdnd11an1n64x5 FILLER_39_1044 ();
 b15zdnd11an1n64x5 FILLER_39_1108 ();
 b15zdnd11an1n64x5 FILLER_39_1172 ();
 b15zdnd11an1n64x5 FILLER_39_1236 ();
 b15zdnd11an1n64x5 FILLER_39_1300 ();
 b15zdnd11an1n64x5 FILLER_39_1364 ();
 b15zdnd11an1n32x5 FILLER_39_1428 ();
 b15zdnd11an1n16x5 FILLER_39_1460 ();
 b15zdnd11an1n08x5 FILLER_39_1476 ();
 b15zdnd00an1n02x5 FILLER_39_1484 ();
 b15zdnd11an1n16x5 FILLER_39_2257 ();
 b15zdnd11an1n08x5 FILLER_39_2273 ();
 b15zdnd00an1n02x5 FILLER_39_2281 ();
 b15zdnd00an1n01x5 FILLER_39_2283 ();
 b15zdnd11an1n64x5 FILLER_40_8 ();
 b15zdnd11an1n64x5 FILLER_40_72 ();
 b15zdnd11an1n64x5 FILLER_40_136 ();
 b15zdnd11an1n64x5 FILLER_40_200 ();
 b15zdnd11an1n64x5 FILLER_40_264 ();
 b15zdnd11an1n64x5 FILLER_40_328 ();
 b15zdnd11an1n64x5 FILLER_40_392 ();
 b15zdnd11an1n64x5 FILLER_40_456 ();
 b15zdnd11an1n64x5 FILLER_40_520 ();
 b15zdnd11an1n64x5 FILLER_40_584 ();
 b15zdnd11an1n64x5 FILLER_40_648 ();
 b15zdnd11an1n04x5 FILLER_40_712 ();
 b15zdnd00an1n02x5 FILLER_40_716 ();
 b15zdnd11an1n64x5 FILLER_40_726 ();
 b15zdnd11an1n64x5 FILLER_40_790 ();
 b15zdnd11an1n64x5 FILLER_40_854 ();
 b15zdnd11an1n32x5 FILLER_40_918 ();
 b15zdnd11an1n08x5 FILLER_40_950 ();
 b15zdnd00an1n02x5 FILLER_40_958 ();
 b15zdnd11an1n64x5 FILLER_40_970 ();
 b15zdnd11an1n64x5 FILLER_40_1034 ();
 b15zdnd11an1n64x5 FILLER_40_1098 ();
 b15zdnd11an1n64x5 FILLER_40_1162 ();
 b15zdnd11an1n64x5 FILLER_40_1226 ();
 b15zdnd11an1n32x5 FILLER_40_1290 ();
 b15zdnd11an1n04x5 FILLER_40_1322 ();
 b15zdnd00an1n02x5 FILLER_40_1326 ();
 b15zdnd11an1n32x5 FILLER_40_1341 ();
 b15zdnd11an1n16x5 FILLER_40_1373 ();
 b15zdnd11an1n04x5 FILLER_40_1389 ();
 b15zdnd00an1n02x5 FILLER_40_1393 ();
 b15zdnd11an1n64x5 FILLER_40_1403 ();
 b15zdnd11an1n08x5 FILLER_40_1467 ();
 b15zdnd00an1n02x5 FILLER_40_1475 ();
 b15zdnd00an1n01x5 FILLER_40_1477 ();
 b15zdnd11an1n08x5 FILLER_40_2265 ();
 b15zdnd00an1n02x5 FILLER_40_2273 ();
 b15zdnd00an1n01x5 FILLER_40_2275 ();
 b15zdnd11an1n64x5 FILLER_41_0 ();
 b15zdnd11an1n64x5 FILLER_41_64 ();
 b15zdnd11an1n64x5 FILLER_41_128 ();
 b15zdnd11an1n64x5 FILLER_41_192 ();
 b15zdnd11an1n64x5 FILLER_41_256 ();
 b15zdnd11an1n64x5 FILLER_41_320 ();
 b15zdnd11an1n64x5 FILLER_41_384 ();
 b15zdnd11an1n64x5 FILLER_41_448 ();
 b15zdnd11an1n64x5 FILLER_41_512 ();
 b15zdnd11an1n64x5 FILLER_41_576 ();
 b15zdnd11an1n64x5 FILLER_41_640 ();
 b15zdnd11an1n64x5 FILLER_41_704 ();
 b15zdnd11an1n16x5 FILLER_41_768 ();
 b15zdnd11an1n04x5 FILLER_41_784 ();
 b15zdnd00an1n02x5 FILLER_41_788 ();
 b15zdnd11an1n32x5 FILLER_41_807 ();
 b15zdnd11an1n04x5 FILLER_41_839 ();
 b15zdnd00an1n02x5 FILLER_41_843 ();
 b15zdnd11an1n64x5 FILLER_41_865 ();
 b15zdnd11an1n64x5 FILLER_41_929 ();
 b15zdnd11an1n08x5 FILLER_41_993 ();
 b15zdnd00an1n01x5 FILLER_41_1001 ();
 b15zdnd11an1n08x5 FILLER_41_1014 ();
 b15zdnd11an1n04x5 FILLER_41_1036 ();
 b15zdnd11an1n64x5 FILLER_41_1056 ();
 b15zdnd11an1n64x5 FILLER_41_1120 ();
 b15zdnd11an1n32x5 FILLER_41_1184 ();
 b15zdnd11an1n16x5 FILLER_41_1216 ();
 b15zdnd11an1n08x5 FILLER_41_1232 ();
 b15zdnd11an1n04x5 FILLER_41_1240 ();
 b15zdnd11an1n04x5 FILLER_41_1254 ();
 b15zdnd11an1n32x5 FILLER_41_1270 ();
 b15zdnd11an1n16x5 FILLER_41_1302 ();
 b15zdnd11an1n08x5 FILLER_41_1318 ();
 b15zdnd11an1n04x5 FILLER_41_1326 ();
 b15zdnd00an1n01x5 FILLER_41_1330 ();
 b15zdnd11an1n64x5 FILLER_41_1341 ();
 b15zdnd11an1n64x5 FILLER_41_1405 ();
 b15zdnd11an1n16x5 FILLER_41_1469 ();
 b15zdnd00an1n01x5 FILLER_41_1485 ();
 b15zdnd11an1n16x5 FILLER_41_2257 ();
 b15zdnd11an1n08x5 FILLER_41_2273 ();
 b15zdnd00an1n02x5 FILLER_41_2281 ();
 b15zdnd00an1n01x5 FILLER_41_2283 ();
 b15zdnd11an1n64x5 FILLER_42_8 ();
 b15zdnd11an1n64x5 FILLER_42_72 ();
 b15zdnd11an1n64x5 FILLER_42_136 ();
 b15zdnd11an1n64x5 FILLER_42_200 ();
 b15zdnd11an1n64x5 FILLER_42_264 ();
 b15zdnd11an1n64x5 FILLER_42_328 ();
 b15zdnd11an1n64x5 FILLER_42_392 ();
 b15zdnd11an1n64x5 FILLER_42_456 ();
 b15zdnd11an1n64x5 FILLER_42_520 ();
 b15zdnd11an1n64x5 FILLER_42_584 ();
 b15zdnd11an1n64x5 FILLER_42_648 ();
 b15zdnd11an1n04x5 FILLER_42_712 ();
 b15zdnd00an1n02x5 FILLER_42_716 ();
 b15zdnd11an1n08x5 FILLER_42_726 ();
 b15zdnd11an1n64x5 FILLER_42_751 ();
 b15zdnd11an1n64x5 FILLER_42_815 ();
 b15zdnd11an1n64x5 FILLER_42_879 ();
 b15zdnd11an1n64x5 FILLER_42_955 ();
 b15zdnd11an1n64x5 FILLER_42_1019 ();
 b15zdnd11an1n32x5 FILLER_42_1083 ();
 b15zdnd11an1n16x5 FILLER_42_1115 ();
 b15zdnd11an1n08x5 FILLER_42_1131 ();
 b15zdnd11an1n04x5 FILLER_42_1139 ();
 b15zdnd11an1n64x5 FILLER_42_1185 ();
 b15zdnd11an1n64x5 FILLER_42_1249 ();
 b15zdnd11an1n64x5 FILLER_42_1313 ();
 b15zdnd11an1n64x5 FILLER_42_1377 ();
 b15zdnd11an1n32x5 FILLER_42_1441 ();
 b15zdnd11an1n04x5 FILLER_42_1473 ();
 b15zdnd00an1n01x5 FILLER_42_1477 ();
 b15zdnd11an1n08x5 FILLER_42_2265 ();
 b15zdnd00an1n02x5 FILLER_42_2273 ();
 b15zdnd00an1n01x5 FILLER_42_2275 ();
 b15zdnd11an1n64x5 FILLER_43_0 ();
 b15zdnd11an1n64x5 FILLER_43_64 ();
 b15zdnd11an1n64x5 FILLER_43_128 ();
 b15zdnd11an1n64x5 FILLER_43_192 ();
 b15zdnd11an1n64x5 FILLER_43_256 ();
 b15zdnd11an1n64x5 FILLER_43_320 ();
 b15zdnd11an1n64x5 FILLER_43_384 ();
 b15zdnd11an1n64x5 FILLER_43_448 ();
 b15zdnd11an1n64x5 FILLER_43_512 ();
 b15zdnd11an1n64x5 FILLER_43_576 ();
 b15zdnd11an1n32x5 FILLER_43_640 ();
 b15zdnd11an1n16x5 FILLER_43_672 ();
 b15zdnd00an1n02x5 FILLER_43_688 ();
 b15zdnd00an1n01x5 FILLER_43_690 ();
 b15zdnd11an1n32x5 FILLER_43_703 ();
 b15zdnd11an1n08x5 FILLER_43_735 ();
 b15zdnd00an1n02x5 FILLER_43_743 ();
 b15zdnd11an1n64x5 FILLER_43_765 ();
 b15zdnd11an1n64x5 FILLER_43_829 ();
 b15zdnd11an1n64x5 FILLER_43_893 ();
 b15zdnd11an1n64x5 FILLER_43_957 ();
 b15zdnd11an1n64x5 FILLER_43_1021 ();
 b15zdnd11an1n64x5 FILLER_43_1085 ();
 b15zdnd11an1n16x5 FILLER_43_1149 ();
 b15zdnd11an1n08x5 FILLER_43_1165 ();
 b15zdnd11an1n04x5 FILLER_43_1173 ();
 b15zdnd00an1n02x5 FILLER_43_1177 ();
 b15zdnd11an1n64x5 FILLER_43_1195 ();
 b15zdnd11an1n64x5 FILLER_43_1259 ();
 b15zdnd11an1n64x5 FILLER_43_1323 ();
 b15zdnd11an1n64x5 FILLER_43_1387 ();
 b15zdnd11an1n32x5 FILLER_43_1451 ();
 b15zdnd00an1n02x5 FILLER_43_1483 ();
 b15zdnd00an1n01x5 FILLER_43_1485 ();
 b15zdnd11an1n16x5 FILLER_43_2257 ();
 b15zdnd11an1n08x5 FILLER_43_2273 ();
 b15zdnd00an1n02x5 FILLER_43_2281 ();
 b15zdnd00an1n01x5 FILLER_43_2283 ();
 b15zdnd11an1n64x5 FILLER_44_8 ();
 b15zdnd11an1n64x5 FILLER_44_72 ();
 b15zdnd11an1n64x5 FILLER_44_136 ();
 b15zdnd11an1n64x5 FILLER_44_200 ();
 b15zdnd11an1n64x5 FILLER_44_264 ();
 b15zdnd11an1n64x5 FILLER_44_328 ();
 b15zdnd11an1n64x5 FILLER_44_392 ();
 b15zdnd11an1n64x5 FILLER_44_456 ();
 b15zdnd11an1n64x5 FILLER_44_520 ();
 b15zdnd11an1n64x5 FILLER_44_584 ();
 b15zdnd11an1n64x5 FILLER_44_648 ();
 b15zdnd11an1n04x5 FILLER_44_712 ();
 b15zdnd00an1n02x5 FILLER_44_716 ();
 b15zdnd11an1n64x5 FILLER_44_726 ();
 b15zdnd11an1n64x5 FILLER_44_790 ();
 b15zdnd11an1n64x5 FILLER_44_854 ();
 b15zdnd11an1n64x5 FILLER_44_918 ();
 b15zdnd11an1n32x5 FILLER_44_982 ();
 b15zdnd11an1n08x5 FILLER_44_1014 ();
 b15zdnd11an1n04x5 FILLER_44_1022 ();
 b15zdnd00an1n02x5 FILLER_44_1026 ();
 b15zdnd11an1n64x5 FILLER_44_1042 ();
 b15zdnd11an1n64x5 FILLER_44_1106 ();
 b15zdnd11an1n64x5 FILLER_44_1170 ();
 b15zdnd11an1n16x5 FILLER_44_1234 ();
 b15zdnd11an1n04x5 FILLER_44_1250 ();
 b15zdnd00an1n01x5 FILLER_44_1254 ();
 b15zdnd11an1n64x5 FILLER_44_1268 ();
 b15zdnd11an1n64x5 FILLER_44_1332 ();
 b15zdnd11an1n64x5 FILLER_44_1396 ();
 b15zdnd11an1n16x5 FILLER_44_1460 ();
 b15zdnd00an1n02x5 FILLER_44_1476 ();
 b15zdnd11an1n08x5 FILLER_44_2265 ();
 b15zdnd00an1n02x5 FILLER_44_2273 ();
 b15zdnd00an1n01x5 FILLER_44_2275 ();
 b15zdnd11an1n64x5 FILLER_45_0 ();
 b15zdnd11an1n64x5 FILLER_45_64 ();
 b15zdnd11an1n64x5 FILLER_45_128 ();
 b15zdnd11an1n64x5 FILLER_45_192 ();
 b15zdnd11an1n64x5 FILLER_45_256 ();
 b15zdnd11an1n64x5 FILLER_45_320 ();
 b15zdnd11an1n64x5 FILLER_45_384 ();
 b15zdnd11an1n64x5 FILLER_45_448 ();
 b15zdnd11an1n64x5 FILLER_45_512 ();
 b15zdnd11an1n64x5 FILLER_45_576 ();
 b15zdnd11an1n32x5 FILLER_45_640 ();
 b15zdnd11an1n16x5 FILLER_45_672 ();
 b15zdnd11an1n16x5 FILLER_45_712 ();
 b15zdnd00an1n02x5 FILLER_45_728 ();
 b15zdnd11an1n64x5 FILLER_45_742 ();
 b15zdnd00an1n01x5 FILLER_45_806 ();
 b15zdnd11an1n32x5 FILLER_45_827 ();
 b15zdnd11an1n16x5 FILLER_45_859 ();
 b15zdnd11an1n64x5 FILLER_45_891 ();
 b15zdnd11an1n64x5 FILLER_45_955 ();
 b15zdnd11an1n64x5 FILLER_45_1019 ();
 b15zdnd11an1n64x5 FILLER_45_1083 ();
 b15zdnd11an1n64x5 FILLER_45_1147 ();
 b15zdnd11an1n64x5 FILLER_45_1211 ();
 b15zdnd11an1n64x5 FILLER_45_1275 ();
 b15zdnd11an1n64x5 FILLER_45_1339 ();
 b15zdnd11an1n64x5 FILLER_45_1403 ();
 b15zdnd11an1n16x5 FILLER_45_1467 ();
 b15zdnd00an1n02x5 FILLER_45_1483 ();
 b15zdnd00an1n01x5 FILLER_45_1485 ();
 b15zdnd11an1n16x5 FILLER_45_2257 ();
 b15zdnd11an1n08x5 FILLER_45_2273 ();
 b15zdnd00an1n02x5 FILLER_45_2281 ();
 b15zdnd00an1n01x5 FILLER_45_2283 ();
 b15zdnd11an1n64x5 FILLER_46_8 ();
 b15zdnd11an1n64x5 FILLER_46_72 ();
 b15zdnd11an1n64x5 FILLER_46_136 ();
 b15zdnd11an1n64x5 FILLER_46_200 ();
 b15zdnd11an1n64x5 FILLER_46_264 ();
 b15zdnd11an1n64x5 FILLER_46_328 ();
 b15zdnd11an1n64x5 FILLER_46_392 ();
 b15zdnd11an1n64x5 FILLER_46_456 ();
 b15zdnd11an1n64x5 FILLER_46_520 ();
 b15zdnd11an1n64x5 FILLER_46_584 ();
 b15zdnd11an1n64x5 FILLER_46_648 ();
 b15zdnd11an1n04x5 FILLER_46_712 ();
 b15zdnd00an1n02x5 FILLER_46_716 ();
 b15zdnd11an1n16x5 FILLER_46_726 ();
 b15zdnd11an1n64x5 FILLER_46_754 ();
 b15zdnd11an1n64x5 FILLER_46_818 ();
 b15zdnd11an1n64x5 FILLER_46_882 ();
 b15zdnd11an1n64x5 FILLER_46_946 ();
 b15zdnd11an1n64x5 FILLER_46_1010 ();
 b15zdnd11an1n32x5 FILLER_46_1074 ();
 b15zdnd11an1n08x5 FILLER_46_1106 ();
 b15zdnd11an1n64x5 FILLER_46_1128 ();
 b15zdnd11an1n64x5 FILLER_46_1192 ();
 b15zdnd11an1n64x5 FILLER_46_1256 ();
 b15zdnd11an1n64x5 FILLER_46_1320 ();
 b15zdnd11an1n64x5 FILLER_46_1384 ();
 b15zdnd11an1n16x5 FILLER_46_1448 ();
 b15zdnd11an1n08x5 FILLER_46_1464 ();
 b15zdnd11an1n04x5 FILLER_46_1472 ();
 b15zdnd00an1n02x5 FILLER_46_1476 ();
 b15zdnd11an1n08x5 FILLER_46_2265 ();
 b15zdnd00an1n02x5 FILLER_46_2273 ();
 b15zdnd00an1n01x5 FILLER_46_2275 ();
 b15zdnd11an1n64x5 FILLER_47_0 ();
 b15zdnd11an1n64x5 FILLER_47_64 ();
 b15zdnd11an1n64x5 FILLER_47_128 ();
 b15zdnd11an1n64x5 FILLER_47_192 ();
 b15zdnd11an1n64x5 FILLER_47_256 ();
 b15zdnd11an1n64x5 FILLER_47_320 ();
 b15zdnd11an1n64x5 FILLER_47_384 ();
 b15zdnd11an1n32x5 FILLER_47_448 ();
 b15zdnd11an1n16x5 FILLER_47_480 ();
 b15zdnd11an1n08x5 FILLER_47_496 ();
 b15zdnd00an1n02x5 FILLER_47_504 ();
 b15zdnd00an1n01x5 FILLER_47_506 ();
 b15zdnd11an1n64x5 FILLER_47_517 ();
 b15zdnd11an1n64x5 FILLER_47_581 ();
 b15zdnd11an1n32x5 FILLER_47_645 ();
 b15zdnd11an1n04x5 FILLER_47_697 ();
 b15zdnd11an1n64x5 FILLER_47_721 ();
 b15zdnd11an1n64x5 FILLER_47_785 ();
 b15zdnd11an1n64x5 FILLER_47_849 ();
 b15zdnd11an1n64x5 FILLER_47_913 ();
 b15zdnd11an1n64x5 FILLER_47_977 ();
 b15zdnd11an1n64x5 FILLER_47_1041 ();
 b15zdnd11an1n64x5 FILLER_47_1105 ();
 b15zdnd11an1n64x5 FILLER_47_1169 ();
 b15zdnd11an1n64x5 FILLER_47_1233 ();
 b15zdnd11an1n64x5 FILLER_47_1297 ();
 b15zdnd11an1n64x5 FILLER_47_1361 ();
 b15zdnd11an1n32x5 FILLER_47_1425 ();
 b15zdnd11an1n16x5 FILLER_47_1457 ();
 b15zdnd11an1n08x5 FILLER_47_1473 ();
 b15zdnd11an1n04x5 FILLER_47_1481 ();
 b15zdnd00an1n01x5 FILLER_47_1485 ();
 b15zdnd11an1n16x5 FILLER_47_2257 ();
 b15zdnd11an1n08x5 FILLER_47_2273 ();
 b15zdnd00an1n02x5 FILLER_47_2281 ();
 b15zdnd00an1n01x5 FILLER_47_2283 ();
 b15zdnd11an1n64x5 FILLER_48_8 ();
 b15zdnd11an1n64x5 FILLER_48_72 ();
 b15zdnd11an1n64x5 FILLER_48_136 ();
 b15zdnd11an1n64x5 FILLER_48_200 ();
 b15zdnd11an1n64x5 FILLER_48_264 ();
 b15zdnd11an1n64x5 FILLER_48_328 ();
 b15zdnd11an1n16x5 FILLER_48_392 ();
 b15zdnd00an1n02x5 FILLER_48_408 ();
 b15zdnd11an1n64x5 FILLER_48_413 ();
 b15zdnd11an1n16x5 FILLER_48_477 ();
 b15zdnd00an1n02x5 FILLER_48_493 ();
 b15zdnd11an1n16x5 FILLER_48_505 ();
 b15zdnd11an1n08x5 FILLER_48_521 ();
 b15zdnd11an1n04x5 FILLER_48_529 ();
 b15zdnd11an1n64x5 FILLER_48_545 ();
 b15zdnd11an1n64x5 FILLER_48_609 ();
 b15zdnd11an1n32x5 FILLER_48_673 ();
 b15zdnd11an1n08x5 FILLER_48_705 ();
 b15zdnd11an1n04x5 FILLER_48_713 ();
 b15zdnd00an1n01x5 FILLER_48_717 ();
 b15zdnd11an1n64x5 FILLER_48_726 ();
 b15zdnd11an1n64x5 FILLER_48_790 ();
 b15zdnd11an1n64x5 FILLER_48_854 ();
 b15zdnd11an1n64x5 FILLER_48_918 ();
 b15zdnd11an1n64x5 FILLER_48_982 ();
 b15zdnd11an1n64x5 FILLER_48_1046 ();
 b15zdnd11an1n64x5 FILLER_48_1110 ();
 b15zdnd11an1n64x5 FILLER_48_1174 ();
 b15zdnd11an1n64x5 FILLER_48_1238 ();
 b15zdnd11an1n64x5 FILLER_48_1302 ();
 b15zdnd11an1n64x5 FILLER_48_1366 ();
 b15zdnd11an1n16x5 FILLER_48_1430 ();
 b15zdnd11an1n08x5 FILLER_48_1446 ();
 b15zdnd00an1n02x5 FILLER_48_1454 ();
 b15zdnd00an1n01x5 FILLER_48_1456 ();
 b15zdnd11an1n04x5 FILLER_48_1473 ();
 b15zdnd00an1n01x5 FILLER_48_1477 ();
 b15zdnd11an1n08x5 FILLER_48_2265 ();
 b15zdnd00an1n02x5 FILLER_48_2273 ();
 b15zdnd00an1n01x5 FILLER_48_2275 ();
 b15zdnd11an1n64x5 FILLER_49_0 ();
 b15zdnd11an1n64x5 FILLER_49_64 ();
 b15zdnd11an1n64x5 FILLER_49_128 ();
 b15zdnd11an1n64x5 FILLER_49_192 ();
 b15zdnd11an1n64x5 FILLER_49_256 ();
 b15zdnd11an1n64x5 FILLER_49_320 ();
 b15zdnd11an1n64x5 FILLER_49_384 ();
 b15zdnd11an1n64x5 FILLER_49_448 ();
 b15zdnd11an1n64x5 FILLER_49_512 ();
 b15zdnd11an1n64x5 FILLER_49_576 ();
 b15zdnd11an1n32x5 FILLER_49_640 ();
 b15zdnd11an1n16x5 FILLER_49_672 ();
 b15zdnd11an1n08x5 FILLER_49_688 ();
 b15zdnd11an1n04x5 FILLER_49_696 ();
 b15zdnd11an1n64x5 FILLER_49_717 ();
 b15zdnd11an1n64x5 FILLER_49_781 ();
 b15zdnd11an1n64x5 FILLER_49_845 ();
 b15zdnd11an1n64x5 FILLER_49_909 ();
 b15zdnd11an1n64x5 FILLER_49_973 ();
 b15zdnd11an1n64x5 FILLER_49_1037 ();
 b15zdnd11an1n64x5 FILLER_49_1101 ();
 b15zdnd11an1n64x5 FILLER_49_1165 ();
 b15zdnd11an1n64x5 FILLER_49_1229 ();
 b15zdnd11an1n64x5 FILLER_49_1293 ();
 b15zdnd11an1n64x5 FILLER_49_1357 ();
 b15zdnd11an1n32x5 FILLER_49_1421 ();
 b15zdnd11an1n04x5 FILLER_49_1453 ();
 b15zdnd00an1n02x5 FILLER_49_1457 ();
 b15zdnd00an1n01x5 FILLER_49_1459 ();
 b15zdnd11an1n08x5 FILLER_49_1474 ();
 b15zdnd11an1n04x5 FILLER_49_1482 ();
 b15zdnd11an1n16x5 FILLER_49_2257 ();
 b15zdnd11an1n08x5 FILLER_49_2273 ();
 b15zdnd00an1n02x5 FILLER_49_2281 ();
 b15zdnd00an1n01x5 FILLER_49_2283 ();
 b15zdnd11an1n64x5 FILLER_50_8 ();
 b15zdnd11an1n64x5 FILLER_50_72 ();
 b15zdnd11an1n64x5 FILLER_50_136 ();
 b15zdnd11an1n64x5 FILLER_50_200 ();
 b15zdnd11an1n64x5 FILLER_50_264 ();
 b15zdnd11an1n64x5 FILLER_50_328 ();
 b15zdnd11an1n64x5 FILLER_50_392 ();
 b15zdnd11an1n64x5 FILLER_50_456 ();
 b15zdnd11an1n64x5 FILLER_50_520 ();
 b15zdnd11an1n64x5 FILLER_50_584 ();
 b15zdnd11an1n04x5 FILLER_50_648 ();
 b15zdnd00an1n01x5 FILLER_50_652 ();
 b15zdnd11an1n08x5 FILLER_50_663 ();
 b15zdnd00an1n02x5 FILLER_50_671 ();
 b15zdnd00an1n01x5 FILLER_50_673 ();
 b15zdnd00an1n02x5 FILLER_50_716 ();
 b15zdnd11an1n64x5 FILLER_50_726 ();
 b15zdnd11an1n64x5 FILLER_50_790 ();
 b15zdnd11an1n64x5 FILLER_50_854 ();
 b15zdnd11an1n64x5 FILLER_50_918 ();
 b15zdnd11an1n16x5 FILLER_50_982 ();
 b15zdnd11an1n04x5 FILLER_50_998 ();
 b15zdnd11an1n08x5 FILLER_50_1044 ();
 b15zdnd11an1n04x5 FILLER_50_1052 ();
 b15zdnd00an1n02x5 FILLER_50_1056 ();
 b15zdnd00an1n01x5 FILLER_50_1058 ();
 b15zdnd11an1n64x5 FILLER_50_1076 ();
 b15zdnd11an1n64x5 FILLER_50_1140 ();
 b15zdnd11an1n64x5 FILLER_50_1204 ();
 b15zdnd11an1n64x5 FILLER_50_1268 ();
 b15zdnd11an1n64x5 FILLER_50_1332 ();
 b15zdnd11an1n64x5 FILLER_50_1396 ();
 b15zdnd11an1n16x5 FILLER_50_1460 ();
 b15zdnd00an1n02x5 FILLER_50_1476 ();
 b15zdnd11an1n08x5 FILLER_50_2265 ();
 b15zdnd00an1n02x5 FILLER_50_2273 ();
 b15zdnd00an1n01x5 FILLER_50_2275 ();
 b15zdnd11an1n64x5 FILLER_51_0 ();
 b15zdnd11an1n64x5 FILLER_51_64 ();
 b15zdnd11an1n64x5 FILLER_51_128 ();
 b15zdnd11an1n64x5 FILLER_51_192 ();
 b15zdnd11an1n64x5 FILLER_51_256 ();
 b15zdnd11an1n64x5 FILLER_51_320 ();
 b15zdnd11an1n64x5 FILLER_51_384 ();
 b15zdnd11an1n64x5 FILLER_51_448 ();
 b15zdnd11an1n64x5 FILLER_51_512 ();
 b15zdnd11an1n64x5 FILLER_51_576 ();
 b15zdnd11an1n08x5 FILLER_51_640 ();
 b15zdnd00an1n02x5 FILLER_51_648 ();
 b15zdnd00an1n01x5 FILLER_51_650 ();
 b15zdnd11an1n16x5 FILLER_51_661 ();
 b15zdnd11an1n08x5 FILLER_51_677 ();
 b15zdnd11an1n64x5 FILLER_51_727 ();
 b15zdnd11an1n64x5 FILLER_51_791 ();
 b15zdnd11an1n64x5 FILLER_51_855 ();
 b15zdnd11an1n64x5 FILLER_51_919 ();
 b15zdnd11an1n16x5 FILLER_51_983 ();
 b15zdnd11an1n08x5 FILLER_51_999 ();
 b15zdnd00an1n02x5 FILLER_51_1007 ();
 b15zdnd11an1n64x5 FILLER_51_1051 ();
 b15zdnd11an1n64x5 FILLER_51_1115 ();
 b15zdnd11an1n64x5 FILLER_51_1179 ();
 b15zdnd11an1n04x5 FILLER_51_1243 ();
 b15zdnd00an1n01x5 FILLER_51_1247 ();
 b15zdnd11an1n64x5 FILLER_51_1260 ();
 b15zdnd11an1n64x5 FILLER_51_1324 ();
 b15zdnd11an1n64x5 FILLER_51_1388 ();
 b15zdnd11an1n32x5 FILLER_51_1452 ();
 b15zdnd00an1n02x5 FILLER_51_1484 ();
 b15zdnd11an1n16x5 FILLER_51_2257 ();
 b15zdnd11an1n08x5 FILLER_51_2273 ();
 b15zdnd00an1n02x5 FILLER_51_2281 ();
 b15zdnd00an1n01x5 FILLER_51_2283 ();
 b15zdnd11an1n64x5 FILLER_52_8 ();
 b15zdnd11an1n64x5 FILLER_52_72 ();
 b15zdnd11an1n64x5 FILLER_52_136 ();
 b15zdnd11an1n64x5 FILLER_52_200 ();
 b15zdnd11an1n64x5 FILLER_52_264 ();
 b15zdnd11an1n64x5 FILLER_52_328 ();
 b15zdnd11an1n64x5 FILLER_52_392 ();
 b15zdnd11an1n64x5 FILLER_52_456 ();
 b15zdnd11an1n64x5 FILLER_52_520 ();
 b15zdnd11an1n64x5 FILLER_52_584 ();
 b15zdnd11an1n64x5 FILLER_52_648 ();
 b15zdnd11an1n04x5 FILLER_52_712 ();
 b15zdnd00an1n02x5 FILLER_52_716 ();
 b15zdnd11an1n64x5 FILLER_52_726 ();
 b15zdnd11an1n64x5 FILLER_52_790 ();
 b15zdnd11an1n64x5 FILLER_52_854 ();
 b15zdnd11an1n64x5 FILLER_52_918 ();
 b15zdnd11an1n64x5 FILLER_52_982 ();
 b15zdnd11an1n64x5 FILLER_52_1046 ();
 b15zdnd11an1n64x5 FILLER_52_1110 ();
 b15zdnd11an1n64x5 FILLER_52_1174 ();
 b15zdnd11an1n64x5 FILLER_52_1238 ();
 b15zdnd11an1n64x5 FILLER_52_1302 ();
 b15zdnd11an1n64x5 FILLER_52_1366 ();
 b15zdnd11an1n32x5 FILLER_52_1430 ();
 b15zdnd11an1n16x5 FILLER_52_1462 ();
 b15zdnd11an1n08x5 FILLER_52_2265 ();
 b15zdnd00an1n02x5 FILLER_52_2273 ();
 b15zdnd00an1n01x5 FILLER_52_2275 ();
 b15zdnd11an1n64x5 FILLER_53_0 ();
 b15zdnd11an1n64x5 FILLER_53_64 ();
 b15zdnd11an1n64x5 FILLER_53_128 ();
 b15zdnd11an1n64x5 FILLER_53_192 ();
 b15zdnd11an1n64x5 FILLER_53_256 ();
 b15zdnd11an1n64x5 FILLER_53_320 ();
 b15zdnd11an1n64x5 FILLER_53_384 ();
 b15zdnd11an1n64x5 FILLER_53_448 ();
 b15zdnd11an1n64x5 FILLER_53_512 ();
 b15zdnd11an1n64x5 FILLER_53_576 ();
 b15zdnd11an1n64x5 FILLER_53_640 ();
 b15zdnd11an1n64x5 FILLER_53_704 ();
 b15zdnd11an1n64x5 FILLER_53_768 ();
 b15zdnd11an1n64x5 FILLER_53_832 ();
 b15zdnd11an1n64x5 FILLER_53_896 ();
 b15zdnd11an1n64x5 FILLER_53_960 ();
 b15zdnd11an1n64x5 FILLER_53_1024 ();
 b15zdnd11an1n64x5 FILLER_53_1088 ();
 b15zdnd11an1n64x5 FILLER_53_1152 ();
 b15zdnd11an1n64x5 FILLER_53_1216 ();
 b15zdnd11an1n64x5 FILLER_53_1280 ();
 b15zdnd11an1n64x5 FILLER_53_1344 ();
 b15zdnd11an1n64x5 FILLER_53_1408 ();
 b15zdnd11an1n08x5 FILLER_53_1472 ();
 b15zdnd11an1n04x5 FILLER_53_1480 ();
 b15zdnd00an1n02x5 FILLER_53_1484 ();
 b15zdnd11an1n16x5 FILLER_53_2257 ();
 b15zdnd11an1n08x5 FILLER_53_2273 ();
 b15zdnd00an1n02x5 FILLER_53_2281 ();
 b15zdnd00an1n01x5 FILLER_53_2283 ();
 b15zdnd11an1n64x5 FILLER_54_8 ();
 b15zdnd11an1n64x5 FILLER_54_72 ();
 b15zdnd11an1n64x5 FILLER_54_136 ();
 b15zdnd11an1n64x5 FILLER_54_200 ();
 b15zdnd11an1n64x5 FILLER_54_264 ();
 b15zdnd11an1n64x5 FILLER_54_328 ();
 b15zdnd11an1n64x5 FILLER_54_392 ();
 b15zdnd11an1n64x5 FILLER_54_456 ();
 b15zdnd11an1n64x5 FILLER_54_520 ();
 b15zdnd11an1n16x5 FILLER_54_584 ();
 b15zdnd11an1n08x5 FILLER_54_600 ();
 b15zdnd11an1n64x5 FILLER_54_628 ();
 b15zdnd11an1n16x5 FILLER_54_692 ();
 b15zdnd11an1n08x5 FILLER_54_708 ();
 b15zdnd00an1n02x5 FILLER_54_716 ();
 b15zdnd11an1n64x5 FILLER_54_726 ();
 b15zdnd11an1n64x5 FILLER_54_790 ();
 b15zdnd11an1n64x5 FILLER_54_854 ();
 b15zdnd11an1n64x5 FILLER_54_918 ();
 b15zdnd11an1n64x5 FILLER_54_982 ();
 b15zdnd11an1n64x5 FILLER_54_1046 ();
 b15zdnd11an1n64x5 FILLER_54_1110 ();
 b15zdnd11an1n64x5 FILLER_54_1174 ();
 b15zdnd11an1n64x5 FILLER_54_1238 ();
 b15zdnd11an1n64x5 FILLER_54_1302 ();
 b15zdnd11an1n64x5 FILLER_54_1366 ();
 b15zdnd11an1n32x5 FILLER_54_1430 ();
 b15zdnd11an1n16x5 FILLER_54_1462 ();
 b15zdnd11an1n08x5 FILLER_54_2265 ();
 b15zdnd00an1n02x5 FILLER_54_2273 ();
 b15zdnd00an1n01x5 FILLER_54_2275 ();
 b15zdnd11an1n64x5 FILLER_55_0 ();
 b15zdnd11an1n64x5 FILLER_55_64 ();
 b15zdnd11an1n64x5 FILLER_55_128 ();
 b15zdnd11an1n64x5 FILLER_55_192 ();
 b15zdnd11an1n64x5 FILLER_55_256 ();
 b15zdnd11an1n64x5 FILLER_55_320 ();
 b15zdnd11an1n64x5 FILLER_55_384 ();
 b15zdnd11an1n64x5 FILLER_55_448 ();
 b15zdnd11an1n64x5 FILLER_55_512 ();
 b15zdnd11an1n64x5 FILLER_55_576 ();
 b15zdnd11an1n64x5 FILLER_55_640 ();
 b15zdnd11an1n64x5 FILLER_55_704 ();
 b15zdnd11an1n64x5 FILLER_55_768 ();
 b15zdnd11an1n64x5 FILLER_55_832 ();
 b15zdnd11an1n64x5 FILLER_55_896 ();
 b15zdnd11an1n64x5 FILLER_55_960 ();
 b15zdnd11an1n16x5 FILLER_55_1024 ();
 b15zdnd11an1n08x5 FILLER_55_1040 ();
 b15zdnd11an1n64x5 FILLER_55_1090 ();
 b15zdnd11an1n64x5 FILLER_55_1154 ();
 b15zdnd11an1n64x5 FILLER_55_1218 ();
 b15zdnd11an1n64x5 FILLER_55_1282 ();
 b15zdnd11an1n64x5 FILLER_55_1346 ();
 b15zdnd11an1n64x5 FILLER_55_1410 ();
 b15zdnd11an1n08x5 FILLER_55_1474 ();
 b15zdnd11an1n04x5 FILLER_55_1482 ();
 b15zdnd11an1n16x5 FILLER_55_2257 ();
 b15zdnd11an1n08x5 FILLER_55_2273 ();
 b15zdnd00an1n02x5 FILLER_55_2281 ();
 b15zdnd00an1n01x5 FILLER_55_2283 ();
 b15zdnd11an1n64x5 FILLER_56_8 ();
 b15zdnd11an1n64x5 FILLER_56_72 ();
 b15zdnd11an1n64x5 FILLER_56_136 ();
 b15zdnd11an1n64x5 FILLER_56_200 ();
 b15zdnd11an1n64x5 FILLER_56_264 ();
 b15zdnd11an1n64x5 FILLER_56_328 ();
 b15zdnd11an1n64x5 FILLER_56_392 ();
 b15zdnd11an1n64x5 FILLER_56_456 ();
 b15zdnd11an1n64x5 FILLER_56_520 ();
 b15zdnd11an1n64x5 FILLER_56_584 ();
 b15zdnd11an1n64x5 FILLER_56_648 ();
 b15zdnd11an1n04x5 FILLER_56_712 ();
 b15zdnd00an1n02x5 FILLER_56_716 ();
 b15zdnd11an1n64x5 FILLER_56_726 ();
 b15zdnd11an1n64x5 FILLER_56_790 ();
 b15zdnd11an1n64x5 FILLER_56_854 ();
 b15zdnd11an1n64x5 FILLER_56_918 ();
 b15zdnd11an1n64x5 FILLER_56_982 ();
 b15zdnd11an1n64x5 FILLER_56_1046 ();
 b15zdnd11an1n64x5 FILLER_56_1110 ();
 b15zdnd11an1n64x5 FILLER_56_1174 ();
 b15zdnd11an1n64x5 FILLER_56_1238 ();
 b15zdnd11an1n64x5 FILLER_56_1302 ();
 b15zdnd11an1n64x5 FILLER_56_1366 ();
 b15zdnd11an1n32x5 FILLER_56_1430 ();
 b15zdnd11an1n16x5 FILLER_56_1462 ();
 b15zdnd11an1n08x5 FILLER_56_2265 ();
 b15zdnd00an1n02x5 FILLER_56_2273 ();
 b15zdnd00an1n01x5 FILLER_56_2275 ();
 b15zdnd11an1n64x5 FILLER_57_0 ();
 b15zdnd11an1n64x5 FILLER_57_64 ();
 b15zdnd11an1n64x5 FILLER_57_128 ();
 b15zdnd11an1n64x5 FILLER_57_192 ();
 b15zdnd11an1n64x5 FILLER_57_256 ();
 b15zdnd11an1n64x5 FILLER_57_320 ();
 b15zdnd11an1n64x5 FILLER_57_384 ();
 b15zdnd11an1n64x5 FILLER_57_448 ();
 b15zdnd11an1n64x5 FILLER_57_512 ();
 b15zdnd11an1n64x5 FILLER_57_576 ();
 b15zdnd11an1n64x5 FILLER_57_640 ();
 b15zdnd11an1n64x5 FILLER_57_704 ();
 b15zdnd11an1n64x5 FILLER_57_768 ();
 b15zdnd11an1n16x5 FILLER_57_832 ();
 b15zdnd00an1n01x5 FILLER_57_848 ();
 b15zdnd11an1n64x5 FILLER_57_891 ();
 b15zdnd11an1n64x5 FILLER_57_955 ();
 b15zdnd11an1n16x5 FILLER_57_1019 ();
 b15zdnd11an1n08x5 FILLER_57_1035 ();
 b15zdnd00an1n02x5 FILLER_57_1043 ();
 b15zdnd11an1n64x5 FILLER_57_1087 ();
 b15zdnd11an1n64x5 FILLER_57_1151 ();
 b15zdnd11an1n64x5 FILLER_57_1215 ();
 b15zdnd11an1n64x5 FILLER_57_1279 ();
 b15zdnd11an1n64x5 FILLER_57_1343 ();
 b15zdnd11an1n64x5 FILLER_57_1407 ();
 b15zdnd11an1n08x5 FILLER_57_1471 ();
 b15zdnd11an1n04x5 FILLER_57_1479 ();
 b15zdnd00an1n02x5 FILLER_57_1483 ();
 b15zdnd00an1n01x5 FILLER_57_1485 ();
 b15zdnd11an1n16x5 FILLER_57_2257 ();
 b15zdnd11an1n08x5 FILLER_57_2273 ();
 b15zdnd00an1n02x5 FILLER_57_2281 ();
 b15zdnd00an1n01x5 FILLER_57_2283 ();
 b15zdnd11an1n64x5 FILLER_58_8 ();
 b15zdnd11an1n64x5 FILLER_58_72 ();
 b15zdnd11an1n64x5 FILLER_58_136 ();
 b15zdnd11an1n64x5 FILLER_58_200 ();
 b15zdnd11an1n64x5 FILLER_58_264 ();
 b15zdnd11an1n64x5 FILLER_58_328 ();
 b15zdnd11an1n64x5 FILLER_58_392 ();
 b15zdnd11an1n64x5 FILLER_58_456 ();
 b15zdnd11an1n64x5 FILLER_58_520 ();
 b15zdnd11an1n64x5 FILLER_58_584 ();
 b15zdnd11an1n64x5 FILLER_58_648 ();
 b15zdnd11an1n04x5 FILLER_58_712 ();
 b15zdnd00an1n02x5 FILLER_58_716 ();
 b15zdnd11an1n64x5 FILLER_58_726 ();
 b15zdnd11an1n64x5 FILLER_58_790 ();
 b15zdnd11an1n64x5 FILLER_58_854 ();
 b15zdnd11an1n64x5 FILLER_58_918 ();
 b15zdnd11an1n64x5 FILLER_58_982 ();
 b15zdnd11an1n64x5 FILLER_58_1046 ();
 b15zdnd11an1n64x5 FILLER_58_1110 ();
 b15zdnd11an1n64x5 FILLER_58_1174 ();
 b15zdnd11an1n64x5 FILLER_58_1238 ();
 b15zdnd11an1n64x5 FILLER_58_1302 ();
 b15zdnd11an1n64x5 FILLER_58_1366 ();
 b15zdnd11an1n32x5 FILLER_58_1430 ();
 b15zdnd11an1n16x5 FILLER_58_1462 ();
 b15zdnd11an1n08x5 FILLER_58_2265 ();
 b15zdnd00an1n02x5 FILLER_58_2273 ();
 b15zdnd00an1n01x5 FILLER_58_2275 ();
 b15zdnd11an1n64x5 FILLER_59_0 ();
 b15zdnd11an1n64x5 FILLER_59_64 ();
 b15zdnd11an1n64x5 FILLER_59_128 ();
 b15zdnd11an1n64x5 FILLER_59_192 ();
 b15zdnd11an1n64x5 FILLER_59_256 ();
 b15zdnd11an1n64x5 FILLER_59_320 ();
 b15zdnd11an1n64x5 FILLER_59_384 ();
 b15zdnd11an1n64x5 FILLER_59_448 ();
 b15zdnd11an1n64x5 FILLER_59_512 ();
 b15zdnd11an1n64x5 FILLER_59_576 ();
 b15zdnd11an1n64x5 FILLER_59_640 ();
 b15zdnd11an1n64x5 FILLER_59_704 ();
 b15zdnd11an1n64x5 FILLER_59_768 ();
 b15zdnd11an1n64x5 FILLER_59_832 ();
 b15zdnd11an1n64x5 FILLER_59_896 ();
 b15zdnd11an1n64x5 FILLER_59_960 ();
 b15zdnd11an1n64x5 FILLER_59_1024 ();
 b15zdnd11an1n64x5 FILLER_59_1088 ();
 b15zdnd11an1n64x5 FILLER_59_1152 ();
 b15zdnd11an1n64x5 FILLER_59_1216 ();
 b15zdnd11an1n64x5 FILLER_59_1280 ();
 b15zdnd11an1n64x5 FILLER_59_1344 ();
 b15zdnd11an1n64x5 FILLER_59_1408 ();
 b15zdnd11an1n08x5 FILLER_59_1472 ();
 b15zdnd11an1n04x5 FILLER_59_1480 ();
 b15zdnd00an1n02x5 FILLER_59_1484 ();
 b15zdnd11an1n16x5 FILLER_59_2257 ();
 b15zdnd11an1n08x5 FILLER_59_2273 ();
 b15zdnd00an1n02x5 FILLER_59_2281 ();
 b15zdnd00an1n01x5 FILLER_59_2283 ();
 b15zdnd11an1n64x5 FILLER_60_8 ();
 b15zdnd11an1n64x5 FILLER_60_72 ();
 b15zdnd11an1n64x5 FILLER_60_136 ();
 b15zdnd11an1n64x5 FILLER_60_200 ();
 b15zdnd11an1n64x5 FILLER_60_264 ();
 b15zdnd11an1n64x5 FILLER_60_328 ();
 b15zdnd11an1n64x5 FILLER_60_392 ();
 b15zdnd11an1n64x5 FILLER_60_456 ();
 b15zdnd11an1n64x5 FILLER_60_520 ();
 b15zdnd11an1n64x5 FILLER_60_584 ();
 b15zdnd11an1n64x5 FILLER_60_648 ();
 b15zdnd11an1n04x5 FILLER_60_712 ();
 b15zdnd00an1n02x5 FILLER_60_716 ();
 b15zdnd11an1n64x5 FILLER_60_726 ();
 b15zdnd11an1n64x5 FILLER_60_790 ();
 b15zdnd11an1n64x5 FILLER_60_854 ();
 b15zdnd11an1n64x5 FILLER_60_918 ();
 b15zdnd11an1n32x5 FILLER_60_982 ();
 b15zdnd00an1n02x5 FILLER_60_1014 ();
 b15zdnd00an1n01x5 FILLER_60_1016 ();
 b15zdnd11an1n64x5 FILLER_60_1059 ();
 b15zdnd11an1n64x5 FILLER_60_1123 ();
 b15zdnd11an1n64x5 FILLER_60_1187 ();
 b15zdnd11an1n64x5 FILLER_60_1251 ();
 b15zdnd11an1n64x5 FILLER_60_1315 ();
 b15zdnd11an1n64x5 FILLER_60_1379 ();
 b15zdnd11an1n32x5 FILLER_60_1443 ();
 b15zdnd00an1n02x5 FILLER_60_1475 ();
 b15zdnd00an1n01x5 FILLER_60_1477 ();
 b15zdnd11an1n08x5 FILLER_60_2265 ();
 b15zdnd00an1n02x5 FILLER_60_2273 ();
 b15zdnd00an1n01x5 FILLER_60_2275 ();
 b15zdnd11an1n64x5 FILLER_61_0 ();
 b15zdnd11an1n64x5 FILLER_61_64 ();
 b15zdnd11an1n64x5 FILLER_61_128 ();
 b15zdnd11an1n64x5 FILLER_61_192 ();
 b15zdnd11an1n64x5 FILLER_61_256 ();
 b15zdnd11an1n64x5 FILLER_61_320 ();
 b15zdnd11an1n64x5 FILLER_61_384 ();
 b15zdnd11an1n64x5 FILLER_61_448 ();
 b15zdnd11an1n64x5 FILLER_61_512 ();
 b15zdnd11an1n64x5 FILLER_61_576 ();
 b15zdnd11an1n64x5 FILLER_61_640 ();
 b15zdnd11an1n64x5 FILLER_61_704 ();
 b15zdnd11an1n64x5 FILLER_61_768 ();
 b15zdnd11an1n64x5 FILLER_61_832 ();
 b15zdnd11an1n64x5 FILLER_61_896 ();
 b15zdnd11an1n32x5 FILLER_61_960 ();
 b15zdnd11an1n08x5 FILLER_61_992 ();
 b15zdnd00an1n02x5 FILLER_61_1000 ();
 b15zdnd11an1n64x5 FILLER_61_1044 ();
 b15zdnd11an1n64x5 FILLER_61_1108 ();
 b15zdnd11an1n64x5 FILLER_61_1172 ();
 b15zdnd11an1n64x5 FILLER_61_1236 ();
 b15zdnd11an1n64x5 FILLER_61_1300 ();
 b15zdnd11an1n64x5 FILLER_61_1364 ();
 b15zdnd11an1n32x5 FILLER_61_1428 ();
 b15zdnd11an1n16x5 FILLER_61_1460 ();
 b15zdnd11an1n08x5 FILLER_61_1476 ();
 b15zdnd00an1n02x5 FILLER_61_1484 ();
 b15zdnd11an1n16x5 FILLER_61_2257 ();
 b15zdnd11an1n08x5 FILLER_61_2273 ();
 b15zdnd00an1n02x5 FILLER_61_2281 ();
 b15zdnd00an1n01x5 FILLER_61_2283 ();
 b15zdnd11an1n64x5 FILLER_62_8 ();
 b15zdnd11an1n64x5 FILLER_62_72 ();
 b15zdnd11an1n64x5 FILLER_62_136 ();
 b15zdnd11an1n64x5 FILLER_62_200 ();
 b15zdnd11an1n64x5 FILLER_62_264 ();
 b15zdnd11an1n64x5 FILLER_62_328 ();
 b15zdnd11an1n64x5 FILLER_62_392 ();
 b15zdnd11an1n64x5 FILLER_62_456 ();
 b15zdnd11an1n64x5 FILLER_62_520 ();
 b15zdnd11an1n64x5 FILLER_62_584 ();
 b15zdnd11an1n64x5 FILLER_62_648 ();
 b15zdnd11an1n04x5 FILLER_62_712 ();
 b15zdnd00an1n02x5 FILLER_62_716 ();
 b15zdnd11an1n08x5 FILLER_62_726 ();
 b15zdnd11an1n04x5 FILLER_62_734 ();
 b15zdnd00an1n02x5 FILLER_62_738 ();
 b15zdnd11an1n64x5 FILLER_62_782 ();
 b15zdnd11an1n32x5 FILLER_62_846 ();
 b15zdnd11an1n16x5 FILLER_62_878 ();
 b15zdnd11an1n08x5 FILLER_62_894 ();
 b15zdnd00an1n02x5 FILLER_62_902 ();
 b15zdnd00an1n01x5 FILLER_62_904 ();
 b15zdnd11an1n64x5 FILLER_62_947 ();
 b15zdnd11an1n64x5 FILLER_62_1011 ();
 b15zdnd11an1n64x5 FILLER_62_1075 ();
 b15zdnd11an1n64x5 FILLER_62_1139 ();
 b15zdnd11an1n64x5 FILLER_62_1203 ();
 b15zdnd11an1n64x5 FILLER_62_1267 ();
 b15zdnd11an1n64x5 FILLER_62_1331 ();
 b15zdnd11an1n64x5 FILLER_62_1395 ();
 b15zdnd11an1n16x5 FILLER_62_1459 ();
 b15zdnd00an1n02x5 FILLER_62_1475 ();
 b15zdnd00an1n01x5 FILLER_62_1477 ();
 b15zdnd11an1n08x5 FILLER_62_2265 ();
 b15zdnd00an1n02x5 FILLER_62_2273 ();
 b15zdnd00an1n01x5 FILLER_62_2275 ();
 b15zdnd11an1n64x5 FILLER_63_0 ();
 b15zdnd11an1n64x5 FILLER_63_64 ();
 b15zdnd11an1n64x5 FILLER_63_128 ();
 b15zdnd11an1n64x5 FILLER_63_192 ();
 b15zdnd11an1n64x5 FILLER_63_256 ();
 b15zdnd11an1n64x5 FILLER_63_320 ();
 b15zdnd11an1n64x5 FILLER_63_384 ();
 b15zdnd11an1n64x5 FILLER_63_448 ();
 b15zdnd11an1n64x5 FILLER_63_512 ();
 b15zdnd11an1n64x5 FILLER_63_576 ();
 b15zdnd11an1n64x5 FILLER_63_640 ();
 b15zdnd11an1n32x5 FILLER_63_704 ();
 b15zdnd11an1n08x5 FILLER_63_736 ();
 b15zdnd11an1n04x5 FILLER_63_744 ();
 b15zdnd00an1n01x5 FILLER_63_748 ();
 b15zdnd11an1n64x5 FILLER_63_791 ();
 b15zdnd11an1n64x5 FILLER_63_855 ();
 b15zdnd11an1n64x5 FILLER_63_919 ();
 b15zdnd11an1n64x5 FILLER_63_983 ();
 b15zdnd11an1n08x5 FILLER_63_1047 ();
 b15zdnd11an1n64x5 FILLER_63_1097 ();
 b15zdnd11an1n64x5 FILLER_63_1161 ();
 b15zdnd11an1n64x5 FILLER_63_1225 ();
 b15zdnd11an1n64x5 FILLER_63_1289 ();
 b15zdnd11an1n64x5 FILLER_63_1353 ();
 b15zdnd11an1n64x5 FILLER_63_1417 ();
 b15zdnd11an1n04x5 FILLER_63_1481 ();
 b15zdnd00an1n01x5 FILLER_63_1485 ();
 b15zdnd11an1n16x5 FILLER_63_2257 ();
 b15zdnd11an1n08x5 FILLER_63_2273 ();
 b15zdnd00an1n02x5 FILLER_63_2281 ();
 b15zdnd00an1n01x5 FILLER_63_2283 ();
 b15zdnd11an1n64x5 FILLER_64_8 ();
 b15zdnd11an1n64x5 FILLER_64_72 ();
 b15zdnd11an1n64x5 FILLER_64_136 ();
 b15zdnd11an1n64x5 FILLER_64_200 ();
 b15zdnd11an1n64x5 FILLER_64_264 ();
 b15zdnd11an1n64x5 FILLER_64_328 ();
 b15zdnd11an1n64x5 FILLER_64_392 ();
 b15zdnd11an1n64x5 FILLER_64_456 ();
 b15zdnd11an1n64x5 FILLER_64_520 ();
 b15zdnd11an1n64x5 FILLER_64_584 ();
 b15zdnd11an1n64x5 FILLER_64_648 ();
 b15zdnd11an1n04x5 FILLER_64_712 ();
 b15zdnd00an1n02x5 FILLER_64_716 ();
 b15zdnd11an1n08x5 FILLER_64_726 ();
 b15zdnd11an1n04x5 FILLER_64_734 ();
 b15zdnd00an1n02x5 FILLER_64_738 ();
 b15zdnd11an1n64x5 FILLER_64_782 ();
 b15zdnd11an1n64x5 FILLER_64_846 ();
 b15zdnd11an1n64x5 FILLER_64_910 ();
 b15zdnd11an1n64x5 FILLER_64_974 ();
 b15zdnd11an1n64x5 FILLER_64_1038 ();
 b15zdnd11an1n64x5 FILLER_64_1102 ();
 b15zdnd11an1n64x5 FILLER_64_1166 ();
 b15zdnd11an1n64x5 FILLER_64_1230 ();
 b15zdnd11an1n64x5 FILLER_64_1294 ();
 b15zdnd11an1n64x5 FILLER_64_1358 ();
 b15zdnd11an1n32x5 FILLER_64_1422 ();
 b15zdnd11an1n16x5 FILLER_64_1454 ();
 b15zdnd11an1n08x5 FILLER_64_1470 ();
 b15zdnd11an1n08x5 FILLER_64_2265 ();
 b15zdnd00an1n02x5 FILLER_64_2273 ();
 b15zdnd00an1n01x5 FILLER_64_2275 ();
 b15zdnd11an1n64x5 FILLER_65_0 ();
 b15zdnd11an1n64x5 FILLER_65_64 ();
 b15zdnd11an1n64x5 FILLER_65_128 ();
 b15zdnd11an1n64x5 FILLER_65_192 ();
 b15zdnd11an1n64x5 FILLER_65_256 ();
 b15zdnd11an1n64x5 FILLER_65_320 ();
 b15zdnd11an1n16x5 FILLER_65_384 ();
 b15zdnd11an1n04x5 FILLER_65_400 ();
 b15zdnd00an1n02x5 FILLER_65_404 ();
 b15zdnd11an1n08x5 FILLER_65_419 ();
 b15zdnd11an1n04x5 FILLER_65_427 ();
 b15zdnd00an1n02x5 FILLER_65_431 ();
 b15zdnd00an1n01x5 FILLER_65_433 ();
 b15zdnd11an1n64x5 FILLER_65_457 ();
 b15zdnd11an1n64x5 FILLER_65_521 ();
 b15zdnd11an1n64x5 FILLER_65_585 ();
 b15zdnd11an1n64x5 FILLER_65_649 ();
 b15zdnd11an1n64x5 FILLER_65_713 ();
 b15zdnd11an1n64x5 FILLER_65_777 ();
 b15zdnd11an1n64x5 FILLER_65_841 ();
 b15zdnd11an1n64x5 FILLER_65_905 ();
 b15zdnd11an1n64x5 FILLER_65_969 ();
 b15zdnd11an1n64x5 FILLER_65_1033 ();
 b15zdnd11an1n64x5 FILLER_65_1097 ();
 b15zdnd11an1n64x5 FILLER_65_1161 ();
 b15zdnd11an1n64x5 FILLER_65_1225 ();
 b15zdnd11an1n64x5 FILLER_65_1289 ();
 b15zdnd11an1n64x5 FILLER_65_1353 ();
 b15zdnd11an1n64x5 FILLER_65_1417 ();
 b15zdnd11an1n04x5 FILLER_65_1481 ();
 b15zdnd00an1n01x5 FILLER_65_1485 ();
 b15zdnd11an1n16x5 FILLER_65_2257 ();
 b15zdnd11an1n08x5 FILLER_65_2273 ();
 b15zdnd00an1n02x5 FILLER_65_2281 ();
 b15zdnd00an1n01x5 FILLER_65_2283 ();
 b15zdnd11an1n64x5 FILLER_66_8 ();
 b15zdnd11an1n64x5 FILLER_66_72 ();
 b15zdnd11an1n64x5 FILLER_66_136 ();
 b15zdnd11an1n64x5 FILLER_66_200 ();
 b15zdnd11an1n64x5 FILLER_66_264 ();
 b15zdnd11an1n64x5 FILLER_66_328 ();
 b15zdnd11an1n64x5 FILLER_66_392 ();
 b15zdnd11an1n64x5 FILLER_66_456 ();
 b15zdnd11an1n64x5 FILLER_66_520 ();
 b15zdnd11an1n64x5 FILLER_66_584 ();
 b15zdnd11an1n64x5 FILLER_66_648 ();
 b15zdnd11an1n04x5 FILLER_66_712 ();
 b15zdnd00an1n02x5 FILLER_66_716 ();
 b15zdnd11an1n64x5 FILLER_66_726 ();
 b15zdnd11an1n64x5 FILLER_66_790 ();
 b15zdnd11an1n64x5 FILLER_66_854 ();
 b15zdnd11an1n64x5 FILLER_66_918 ();
 b15zdnd11an1n64x5 FILLER_66_982 ();
 b15zdnd11an1n64x5 FILLER_66_1046 ();
 b15zdnd11an1n64x5 FILLER_66_1110 ();
 b15zdnd11an1n64x5 FILLER_66_1174 ();
 b15zdnd11an1n64x5 FILLER_66_1238 ();
 b15zdnd11an1n64x5 FILLER_66_1302 ();
 b15zdnd11an1n64x5 FILLER_66_1366 ();
 b15zdnd11an1n32x5 FILLER_66_1430 ();
 b15zdnd11an1n16x5 FILLER_66_1462 ();
 b15zdnd11an1n08x5 FILLER_66_2265 ();
 b15zdnd00an1n02x5 FILLER_66_2273 ();
 b15zdnd00an1n01x5 FILLER_66_2275 ();
 b15zdnd11an1n64x5 FILLER_67_0 ();
 b15zdnd11an1n64x5 FILLER_67_64 ();
 b15zdnd11an1n64x5 FILLER_67_128 ();
 b15zdnd11an1n64x5 FILLER_67_192 ();
 b15zdnd11an1n64x5 FILLER_67_256 ();
 b15zdnd11an1n64x5 FILLER_67_320 ();
 b15zdnd11an1n64x5 FILLER_67_384 ();
 b15zdnd11an1n04x5 FILLER_67_448 ();
 b15zdnd00an1n01x5 FILLER_67_452 ();
 b15zdnd11an1n64x5 FILLER_67_476 ();
 b15zdnd11an1n64x5 FILLER_67_540 ();
 b15zdnd11an1n64x5 FILLER_67_604 ();
 b15zdnd11an1n32x5 FILLER_67_668 ();
 b15zdnd11an1n08x5 FILLER_67_700 ();
 b15zdnd00an1n02x5 FILLER_67_708 ();
 b15zdnd00an1n01x5 FILLER_67_710 ();
 b15zdnd11an1n64x5 FILLER_67_753 ();
 b15zdnd11an1n64x5 FILLER_67_817 ();
 b15zdnd11an1n64x5 FILLER_67_881 ();
 b15zdnd11an1n64x5 FILLER_67_945 ();
 b15zdnd11an1n64x5 FILLER_67_1009 ();
 b15zdnd11an1n64x5 FILLER_67_1073 ();
 b15zdnd11an1n64x5 FILLER_67_1137 ();
 b15zdnd11an1n64x5 FILLER_67_1201 ();
 b15zdnd11an1n64x5 FILLER_67_1265 ();
 b15zdnd11an1n64x5 FILLER_67_1329 ();
 b15zdnd11an1n64x5 FILLER_67_1393 ();
 b15zdnd11an1n16x5 FILLER_67_1457 ();
 b15zdnd11an1n08x5 FILLER_67_1473 ();
 b15zdnd11an1n04x5 FILLER_67_1481 ();
 b15zdnd00an1n01x5 FILLER_67_1485 ();
 b15zdnd11an1n16x5 FILLER_67_2257 ();
 b15zdnd11an1n08x5 FILLER_67_2273 ();
 b15zdnd00an1n02x5 FILLER_67_2281 ();
 b15zdnd00an1n01x5 FILLER_67_2283 ();
 b15zdnd11an1n64x5 FILLER_68_8 ();
 b15zdnd11an1n64x5 FILLER_68_72 ();
 b15zdnd11an1n64x5 FILLER_68_136 ();
 b15zdnd11an1n64x5 FILLER_68_200 ();
 b15zdnd11an1n64x5 FILLER_68_264 ();
 b15zdnd11an1n64x5 FILLER_68_328 ();
 b15zdnd11an1n32x5 FILLER_68_392 ();
 b15zdnd00an1n01x5 FILLER_68_424 ();
 b15zdnd11an1n64x5 FILLER_68_431 ();
 b15zdnd11an1n64x5 FILLER_68_495 ();
 b15zdnd11an1n64x5 FILLER_68_559 ();
 b15zdnd11an1n64x5 FILLER_68_623 ();
 b15zdnd11an1n16x5 FILLER_68_687 ();
 b15zdnd11an1n08x5 FILLER_68_703 ();
 b15zdnd11an1n04x5 FILLER_68_711 ();
 b15zdnd00an1n02x5 FILLER_68_715 ();
 b15zdnd00an1n01x5 FILLER_68_717 ();
 b15zdnd11an1n64x5 FILLER_68_726 ();
 b15zdnd11an1n64x5 FILLER_68_790 ();
 b15zdnd11an1n64x5 FILLER_68_854 ();
 b15zdnd11an1n64x5 FILLER_68_918 ();
 b15zdnd11an1n64x5 FILLER_68_982 ();
 b15zdnd11an1n64x5 FILLER_68_1046 ();
 b15zdnd11an1n64x5 FILLER_68_1110 ();
 b15zdnd11an1n64x5 FILLER_68_1174 ();
 b15zdnd11an1n64x5 FILLER_68_1238 ();
 b15zdnd11an1n64x5 FILLER_68_1302 ();
 b15zdnd11an1n64x5 FILLER_68_1366 ();
 b15zdnd11an1n32x5 FILLER_68_1430 ();
 b15zdnd11an1n16x5 FILLER_68_1462 ();
 b15zdnd11an1n08x5 FILLER_68_2265 ();
 b15zdnd00an1n02x5 FILLER_68_2273 ();
 b15zdnd00an1n01x5 FILLER_68_2275 ();
 b15zdnd11an1n64x5 FILLER_69_0 ();
 b15zdnd11an1n64x5 FILLER_69_64 ();
 b15zdnd11an1n64x5 FILLER_69_128 ();
 b15zdnd11an1n64x5 FILLER_69_192 ();
 b15zdnd11an1n64x5 FILLER_69_256 ();
 b15zdnd11an1n64x5 FILLER_69_320 ();
 b15zdnd11an1n64x5 FILLER_69_384 ();
 b15zdnd11an1n64x5 FILLER_69_448 ();
 b15zdnd11an1n64x5 FILLER_69_512 ();
 b15zdnd11an1n64x5 FILLER_69_576 ();
 b15zdnd11an1n64x5 FILLER_69_640 ();
 b15zdnd11an1n04x5 FILLER_69_704 ();
 b15zdnd11an1n64x5 FILLER_69_750 ();
 b15zdnd11an1n64x5 FILLER_69_814 ();
 b15zdnd11an1n64x5 FILLER_69_878 ();
 b15zdnd11an1n64x5 FILLER_69_942 ();
 b15zdnd11an1n64x5 FILLER_69_1006 ();
 b15zdnd11an1n64x5 FILLER_69_1070 ();
 b15zdnd11an1n64x5 FILLER_69_1134 ();
 b15zdnd11an1n64x5 FILLER_69_1198 ();
 b15zdnd11an1n64x5 FILLER_69_1262 ();
 b15zdnd11an1n64x5 FILLER_69_1326 ();
 b15zdnd11an1n64x5 FILLER_69_1390 ();
 b15zdnd11an1n32x5 FILLER_69_1454 ();
 b15zdnd11an1n16x5 FILLER_69_2257 ();
 b15zdnd11an1n08x5 FILLER_69_2273 ();
 b15zdnd00an1n02x5 FILLER_69_2281 ();
 b15zdnd00an1n01x5 FILLER_69_2283 ();
 b15zdnd11an1n64x5 FILLER_70_8 ();
 b15zdnd11an1n64x5 FILLER_70_72 ();
 b15zdnd11an1n64x5 FILLER_70_136 ();
 b15zdnd11an1n64x5 FILLER_70_200 ();
 b15zdnd11an1n64x5 FILLER_70_264 ();
 b15zdnd11an1n64x5 FILLER_70_328 ();
 b15zdnd11an1n64x5 FILLER_70_392 ();
 b15zdnd11an1n64x5 FILLER_70_456 ();
 b15zdnd11an1n64x5 FILLER_70_520 ();
 b15zdnd11an1n64x5 FILLER_70_584 ();
 b15zdnd11an1n64x5 FILLER_70_648 ();
 b15zdnd11an1n04x5 FILLER_70_712 ();
 b15zdnd00an1n02x5 FILLER_70_716 ();
 b15zdnd11an1n64x5 FILLER_70_726 ();
 b15zdnd11an1n64x5 FILLER_70_790 ();
 b15zdnd11an1n64x5 FILLER_70_854 ();
 b15zdnd11an1n64x5 FILLER_70_918 ();
 b15zdnd11an1n64x5 FILLER_70_982 ();
 b15zdnd11an1n64x5 FILLER_70_1046 ();
 b15zdnd11an1n64x5 FILLER_70_1110 ();
 b15zdnd11an1n64x5 FILLER_70_1174 ();
 b15zdnd11an1n64x5 FILLER_70_1238 ();
 b15zdnd11an1n64x5 FILLER_70_1302 ();
 b15zdnd11an1n64x5 FILLER_70_1366 ();
 b15zdnd11an1n32x5 FILLER_70_1430 ();
 b15zdnd11an1n16x5 FILLER_70_1462 ();
 b15zdnd11an1n08x5 FILLER_70_2265 ();
 b15zdnd00an1n02x5 FILLER_70_2273 ();
 b15zdnd00an1n01x5 FILLER_70_2275 ();
 b15zdnd11an1n64x5 FILLER_71_0 ();
 b15zdnd11an1n64x5 FILLER_71_64 ();
 b15zdnd11an1n64x5 FILLER_71_128 ();
 b15zdnd11an1n64x5 FILLER_71_192 ();
 b15zdnd11an1n64x5 FILLER_71_256 ();
 b15zdnd11an1n64x5 FILLER_71_320 ();
 b15zdnd11an1n64x5 FILLER_71_384 ();
 b15zdnd11an1n64x5 FILLER_71_448 ();
 b15zdnd11an1n64x5 FILLER_71_512 ();
 b15zdnd11an1n64x5 FILLER_71_576 ();
 b15zdnd11an1n32x5 FILLER_71_640 ();
 b15zdnd11an1n08x5 FILLER_71_672 ();
 b15zdnd00an1n02x5 FILLER_71_680 ();
 b15zdnd00an1n01x5 FILLER_71_682 ();
 b15zdnd11an1n64x5 FILLER_71_725 ();
 b15zdnd11an1n64x5 FILLER_71_789 ();
 b15zdnd11an1n64x5 FILLER_71_853 ();
 b15zdnd11an1n64x5 FILLER_71_917 ();
 b15zdnd11an1n64x5 FILLER_71_981 ();
 b15zdnd11an1n64x5 FILLER_71_1045 ();
 b15zdnd11an1n64x5 FILLER_71_1109 ();
 b15zdnd11an1n64x5 FILLER_71_1173 ();
 b15zdnd11an1n64x5 FILLER_71_1237 ();
 b15zdnd11an1n64x5 FILLER_71_1301 ();
 b15zdnd11an1n64x5 FILLER_71_1365 ();
 b15zdnd11an1n32x5 FILLER_71_1429 ();
 b15zdnd11an1n16x5 FILLER_71_1461 ();
 b15zdnd11an1n08x5 FILLER_71_1477 ();
 b15zdnd00an1n01x5 FILLER_71_1485 ();
 b15zdnd11an1n16x5 FILLER_71_2257 ();
 b15zdnd11an1n08x5 FILLER_71_2273 ();
 b15zdnd00an1n02x5 FILLER_71_2281 ();
 b15zdnd00an1n01x5 FILLER_71_2283 ();
 b15zdnd11an1n64x5 FILLER_72_8 ();
 b15zdnd11an1n64x5 FILLER_72_72 ();
 b15zdnd11an1n64x5 FILLER_72_136 ();
 b15zdnd11an1n64x5 FILLER_72_200 ();
 b15zdnd11an1n64x5 FILLER_72_264 ();
 b15zdnd11an1n64x5 FILLER_72_328 ();
 b15zdnd11an1n08x5 FILLER_72_392 ();
 b15zdnd00an1n02x5 FILLER_72_400 ();
 b15zdnd00an1n01x5 FILLER_72_402 ();
 b15zdnd11an1n64x5 FILLER_72_408 ();
 b15zdnd11an1n64x5 FILLER_72_472 ();
 b15zdnd11an1n64x5 FILLER_72_536 ();
 b15zdnd11an1n64x5 FILLER_72_600 ();
 b15zdnd11an1n32x5 FILLER_72_664 ();
 b15zdnd11an1n16x5 FILLER_72_696 ();
 b15zdnd11an1n04x5 FILLER_72_712 ();
 b15zdnd00an1n02x5 FILLER_72_716 ();
 b15zdnd11an1n64x5 FILLER_72_726 ();
 b15zdnd11an1n64x5 FILLER_72_790 ();
 b15zdnd11an1n64x5 FILLER_72_854 ();
 b15zdnd11an1n64x5 FILLER_72_918 ();
 b15zdnd11an1n64x5 FILLER_72_982 ();
 b15zdnd11an1n64x5 FILLER_72_1046 ();
 b15zdnd11an1n64x5 FILLER_72_1110 ();
 b15zdnd11an1n64x5 FILLER_72_1174 ();
 b15zdnd11an1n64x5 FILLER_72_1238 ();
 b15zdnd11an1n64x5 FILLER_72_1302 ();
 b15zdnd11an1n64x5 FILLER_72_1366 ();
 b15zdnd11an1n32x5 FILLER_72_1430 ();
 b15zdnd11an1n16x5 FILLER_72_1462 ();
 b15zdnd11an1n08x5 FILLER_72_2265 ();
 b15zdnd00an1n02x5 FILLER_72_2273 ();
 b15zdnd00an1n01x5 FILLER_72_2275 ();
 b15zdnd11an1n64x5 FILLER_73_0 ();
 b15zdnd11an1n64x5 FILLER_73_64 ();
 b15zdnd11an1n64x5 FILLER_73_128 ();
 b15zdnd11an1n64x5 FILLER_73_192 ();
 b15zdnd11an1n64x5 FILLER_73_256 ();
 b15zdnd11an1n64x5 FILLER_73_320 ();
 b15zdnd11an1n64x5 FILLER_73_384 ();
 b15zdnd11an1n64x5 FILLER_73_448 ();
 b15zdnd11an1n64x5 FILLER_73_512 ();
 b15zdnd11an1n64x5 FILLER_73_576 ();
 b15zdnd11an1n64x5 FILLER_73_640 ();
 b15zdnd11an1n64x5 FILLER_73_704 ();
 b15zdnd11an1n64x5 FILLER_73_768 ();
 b15zdnd11an1n64x5 FILLER_73_832 ();
 b15zdnd11an1n64x5 FILLER_73_896 ();
 b15zdnd11an1n64x5 FILLER_73_960 ();
 b15zdnd11an1n64x5 FILLER_73_1024 ();
 b15zdnd11an1n64x5 FILLER_73_1088 ();
 b15zdnd11an1n64x5 FILLER_73_1152 ();
 b15zdnd11an1n64x5 FILLER_73_1216 ();
 b15zdnd11an1n64x5 FILLER_73_1280 ();
 b15zdnd11an1n64x5 FILLER_73_1344 ();
 b15zdnd11an1n64x5 FILLER_73_1408 ();
 b15zdnd11an1n08x5 FILLER_73_1472 ();
 b15zdnd11an1n04x5 FILLER_73_1480 ();
 b15zdnd00an1n02x5 FILLER_73_1484 ();
 b15zdnd11an1n16x5 FILLER_73_2257 ();
 b15zdnd11an1n08x5 FILLER_73_2273 ();
 b15zdnd00an1n02x5 FILLER_73_2281 ();
 b15zdnd00an1n01x5 FILLER_73_2283 ();
 b15zdnd11an1n64x5 FILLER_74_8 ();
 b15zdnd11an1n64x5 FILLER_74_72 ();
 b15zdnd11an1n64x5 FILLER_74_136 ();
 b15zdnd11an1n64x5 FILLER_74_200 ();
 b15zdnd11an1n64x5 FILLER_74_264 ();
 b15zdnd11an1n64x5 FILLER_74_328 ();
 b15zdnd11an1n64x5 FILLER_74_392 ();
 b15zdnd11an1n64x5 FILLER_74_456 ();
 b15zdnd11an1n64x5 FILLER_74_520 ();
 b15zdnd11an1n64x5 FILLER_74_584 ();
 b15zdnd11an1n64x5 FILLER_74_648 ();
 b15zdnd11an1n04x5 FILLER_74_712 ();
 b15zdnd00an1n02x5 FILLER_74_716 ();
 b15zdnd11an1n32x5 FILLER_74_726 ();
 b15zdnd11an1n16x5 FILLER_74_758 ();
 b15zdnd11an1n08x5 FILLER_74_774 ();
 b15zdnd11an1n64x5 FILLER_74_824 ();
 b15zdnd11an1n64x5 FILLER_74_888 ();
 b15zdnd11an1n64x5 FILLER_74_952 ();
 b15zdnd11an1n64x5 FILLER_74_1016 ();
 b15zdnd11an1n64x5 FILLER_74_1080 ();
 b15zdnd11an1n64x5 FILLER_74_1144 ();
 b15zdnd11an1n64x5 FILLER_74_1208 ();
 b15zdnd11an1n64x5 FILLER_74_1272 ();
 b15zdnd11an1n64x5 FILLER_74_1336 ();
 b15zdnd11an1n64x5 FILLER_74_1400 ();
 b15zdnd11an1n08x5 FILLER_74_1464 ();
 b15zdnd11an1n04x5 FILLER_74_1472 ();
 b15zdnd00an1n02x5 FILLER_74_1476 ();
 b15zdnd11an1n08x5 FILLER_74_2265 ();
 b15zdnd00an1n02x5 FILLER_74_2273 ();
 b15zdnd00an1n01x5 FILLER_74_2275 ();
 b15zdnd11an1n64x5 FILLER_75_0 ();
 b15zdnd11an1n64x5 FILLER_75_64 ();
 b15zdnd11an1n64x5 FILLER_75_128 ();
 b15zdnd11an1n64x5 FILLER_75_192 ();
 b15zdnd11an1n64x5 FILLER_75_256 ();
 b15zdnd11an1n64x5 FILLER_75_320 ();
 b15zdnd11an1n64x5 FILLER_75_384 ();
 b15zdnd11an1n64x5 FILLER_75_448 ();
 b15zdnd11an1n64x5 FILLER_75_512 ();
 b15zdnd11an1n64x5 FILLER_75_576 ();
 b15zdnd11an1n64x5 FILLER_75_640 ();
 b15zdnd11an1n64x5 FILLER_75_704 ();
 b15zdnd11an1n64x5 FILLER_75_768 ();
 b15zdnd11an1n64x5 FILLER_75_832 ();
 b15zdnd11an1n64x5 FILLER_75_896 ();
 b15zdnd11an1n64x5 FILLER_75_960 ();
 b15zdnd11an1n64x5 FILLER_75_1024 ();
 b15zdnd11an1n64x5 FILLER_75_1088 ();
 b15zdnd11an1n64x5 FILLER_75_1152 ();
 b15zdnd11an1n64x5 FILLER_75_1216 ();
 b15zdnd11an1n64x5 FILLER_75_1280 ();
 b15zdnd11an1n64x5 FILLER_75_1344 ();
 b15zdnd11an1n64x5 FILLER_75_1408 ();
 b15zdnd11an1n08x5 FILLER_75_1472 ();
 b15zdnd11an1n04x5 FILLER_75_1480 ();
 b15zdnd00an1n02x5 FILLER_75_1484 ();
 b15zdnd11an1n16x5 FILLER_75_2257 ();
 b15zdnd11an1n08x5 FILLER_75_2273 ();
 b15zdnd00an1n02x5 FILLER_75_2281 ();
 b15zdnd00an1n01x5 FILLER_75_2283 ();
 b15zdnd11an1n64x5 FILLER_76_8 ();
 b15zdnd11an1n64x5 FILLER_76_72 ();
 b15zdnd11an1n64x5 FILLER_76_136 ();
 b15zdnd11an1n64x5 FILLER_76_200 ();
 b15zdnd11an1n64x5 FILLER_76_264 ();
 b15zdnd11an1n64x5 FILLER_76_328 ();
 b15zdnd11an1n64x5 FILLER_76_392 ();
 b15zdnd11an1n64x5 FILLER_76_456 ();
 b15zdnd11an1n64x5 FILLER_76_520 ();
 b15zdnd11an1n64x5 FILLER_76_584 ();
 b15zdnd11an1n64x5 FILLER_76_648 ();
 b15zdnd11an1n04x5 FILLER_76_712 ();
 b15zdnd00an1n02x5 FILLER_76_716 ();
 b15zdnd11an1n64x5 FILLER_76_726 ();
 b15zdnd11an1n64x5 FILLER_76_790 ();
 b15zdnd11an1n64x5 FILLER_76_854 ();
 b15zdnd11an1n64x5 FILLER_76_918 ();
 b15zdnd11an1n08x5 FILLER_76_982 ();
 b15zdnd00an1n02x5 FILLER_76_990 ();
 b15zdnd11an1n64x5 FILLER_76_1036 ();
 b15zdnd11an1n64x5 FILLER_76_1100 ();
 b15zdnd11an1n64x5 FILLER_76_1164 ();
 b15zdnd11an1n64x5 FILLER_76_1228 ();
 b15zdnd11an1n64x5 FILLER_76_1292 ();
 b15zdnd11an1n64x5 FILLER_76_1356 ();
 b15zdnd11an1n32x5 FILLER_76_1420 ();
 b15zdnd11an1n16x5 FILLER_76_1452 ();
 b15zdnd11an1n08x5 FILLER_76_1468 ();
 b15zdnd00an1n02x5 FILLER_76_1476 ();
 b15zdnd11an1n08x5 FILLER_76_2265 ();
 b15zdnd00an1n02x5 FILLER_76_2273 ();
 b15zdnd00an1n01x5 FILLER_76_2275 ();
 b15zdnd11an1n64x5 FILLER_77_0 ();
 b15zdnd11an1n64x5 FILLER_77_64 ();
 b15zdnd11an1n64x5 FILLER_77_128 ();
 b15zdnd11an1n64x5 FILLER_77_192 ();
 b15zdnd11an1n64x5 FILLER_77_256 ();
 b15zdnd11an1n64x5 FILLER_77_320 ();
 b15zdnd11an1n64x5 FILLER_77_384 ();
 b15zdnd11an1n64x5 FILLER_77_448 ();
 b15zdnd11an1n64x5 FILLER_77_512 ();
 b15zdnd11an1n64x5 FILLER_77_576 ();
 b15zdnd11an1n64x5 FILLER_77_640 ();
 b15zdnd00an1n02x5 FILLER_77_704 ();
 b15zdnd11an1n64x5 FILLER_77_748 ();
 b15zdnd11an1n64x5 FILLER_77_812 ();
 b15zdnd11an1n64x5 FILLER_77_876 ();
 b15zdnd11an1n32x5 FILLER_77_940 ();
 b15zdnd11an1n08x5 FILLER_77_972 ();
 b15zdnd11an1n04x5 FILLER_77_980 ();
 b15zdnd00an1n02x5 FILLER_77_984 ();
 b15zdnd11an1n04x5 FILLER_77_989 ();
 b15zdnd00an1n02x5 FILLER_77_993 ();
 b15zdnd11an1n64x5 FILLER_77_998 ();
 b15zdnd11an1n64x5 FILLER_77_1062 ();
 b15zdnd11an1n64x5 FILLER_77_1126 ();
 b15zdnd11an1n64x5 FILLER_77_1190 ();
 b15zdnd11an1n64x5 FILLER_77_1254 ();
 b15zdnd11an1n64x5 FILLER_77_1318 ();
 b15zdnd11an1n64x5 FILLER_77_1382 ();
 b15zdnd11an1n32x5 FILLER_77_1446 ();
 b15zdnd11an1n08x5 FILLER_77_1478 ();
 b15zdnd11an1n16x5 FILLER_77_2257 ();
 b15zdnd11an1n08x5 FILLER_77_2273 ();
 b15zdnd00an1n02x5 FILLER_77_2281 ();
 b15zdnd00an1n01x5 FILLER_77_2283 ();
 b15zdnd11an1n64x5 FILLER_78_8 ();
 b15zdnd11an1n64x5 FILLER_78_72 ();
 b15zdnd11an1n64x5 FILLER_78_136 ();
 b15zdnd11an1n64x5 FILLER_78_200 ();
 b15zdnd11an1n64x5 FILLER_78_264 ();
 b15zdnd11an1n64x5 FILLER_78_328 ();
 b15zdnd11an1n64x5 FILLER_78_392 ();
 b15zdnd11an1n64x5 FILLER_78_456 ();
 b15zdnd11an1n64x5 FILLER_78_520 ();
 b15zdnd11an1n64x5 FILLER_78_584 ();
 b15zdnd11an1n64x5 FILLER_78_648 ();
 b15zdnd11an1n04x5 FILLER_78_712 ();
 b15zdnd00an1n02x5 FILLER_78_716 ();
 b15zdnd11an1n64x5 FILLER_78_726 ();
 b15zdnd11an1n64x5 FILLER_78_790 ();
 b15zdnd11an1n64x5 FILLER_78_854 ();
 b15zdnd11an1n64x5 FILLER_78_918 ();
 b15zdnd11an1n04x5 FILLER_78_982 ();
 b15zdnd00an1n02x5 FILLER_78_986 ();
 b15zdnd00an1n01x5 FILLER_78_988 ();
 b15zdnd11an1n04x5 FILLER_78_992 ();
 b15zdnd11an1n64x5 FILLER_78_1040 ();
 b15zdnd11an1n64x5 FILLER_78_1104 ();
 b15zdnd11an1n64x5 FILLER_78_1168 ();
 b15zdnd11an1n64x5 FILLER_78_1232 ();
 b15zdnd11an1n64x5 FILLER_78_1296 ();
 b15zdnd11an1n64x5 FILLER_78_1360 ();
 b15zdnd11an1n32x5 FILLER_78_1424 ();
 b15zdnd11an1n16x5 FILLER_78_1456 ();
 b15zdnd11an1n04x5 FILLER_78_1472 ();
 b15zdnd00an1n02x5 FILLER_78_1476 ();
 b15zdnd11an1n08x5 FILLER_78_2265 ();
 b15zdnd00an1n02x5 FILLER_78_2273 ();
 b15zdnd00an1n01x5 FILLER_78_2275 ();
 b15zdnd11an1n64x5 FILLER_79_0 ();
 b15zdnd11an1n64x5 FILLER_79_64 ();
 b15zdnd11an1n64x5 FILLER_79_128 ();
 b15zdnd11an1n64x5 FILLER_79_192 ();
 b15zdnd11an1n64x5 FILLER_79_256 ();
 b15zdnd11an1n64x5 FILLER_79_320 ();
 b15zdnd11an1n64x5 FILLER_79_384 ();
 b15zdnd11an1n64x5 FILLER_79_448 ();
 b15zdnd11an1n64x5 FILLER_79_512 ();
 b15zdnd11an1n64x5 FILLER_79_576 ();
 b15zdnd11an1n64x5 FILLER_79_640 ();
 b15zdnd11an1n64x5 FILLER_79_704 ();
 b15zdnd11an1n64x5 FILLER_79_768 ();
 b15zdnd11an1n64x5 FILLER_79_832 ();
 b15zdnd11an1n64x5 FILLER_79_896 ();
 b15zdnd11an1n08x5 FILLER_79_960 ();
 b15zdnd11an1n04x5 FILLER_79_1012 ();
 b15zdnd11an1n64x5 FILLER_79_1019 ();
 b15zdnd11an1n64x5 FILLER_79_1083 ();
 b15zdnd11an1n64x5 FILLER_79_1147 ();
 b15zdnd11an1n64x5 FILLER_79_1211 ();
 b15zdnd11an1n64x5 FILLER_79_1275 ();
 b15zdnd11an1n64x5 FILLER_79_1339 ();
 b15zdnd11an1n64x5 FILLER_79_1403 ();
 b15zdnd11an1n16x5 FILLER_79_1467 ();
 b15zdnd00an1n02x5 FILLER_79_1483 ();
 b15zdnd00an1n01x5 FILLER_79_1485 ();
 b15zdnd11an1n16x5 FILLER_79_2257 ();
 b15zdnd11an1n08x5 FILLER_79_2273 ();
 b15zdnd00an1n02x5 FILLER_79_2281 ();
 b15zdnd00an1n01x5 FILLER_79_2283 ();
 b15zdnd11an1n64x5 FILLER_80_8 ();
 b15zdnd11an1n64x5 FILLER_80_72 ();
 b15zdnd11an1n64x5 FILLER_80_136 ();
 b15zdnd11an1n64x5 FILLER_80_200 ();
 b15zdnd11an1n64x5 FILLER_80_264 ();
 b15zdnd11an1n64x5 FILLER_80_328 ();
 b15zdnd11an1n64x5 FILLER_80_392 ();
 b15zdnd11an1n64x5 FILLER_80_456 ();
 b15zdnd11an1n64x5 FILLER_80_520 ();
 b15zdnd11an1n64x5 FILLER_80_584 ();
 b15zdnd11an1n64x5 FILLER_80_648 ();
 b15zdnd11an1n04x5 FILLER_80_712 ();
 b15zdnd00an1n02x5 FILLER_80_716 ();
 b15zdnd11an1n16x5 FILLER_80_726 ();
 b15zdnd11an1n08x5 FILLER_80_742 ();
 b15zdnd11an1n64x5 FILLER_80_753 ();
 b15zdnd11an1n64x5 FILLER_80_817 ();
 b15zdnd11an1n64x5 FILLER_80_881 ();
 b15zdnd11an1n32x5 FILLER_80_945 ();
 b15zdnd11an1n16x5 FILLER_80_977 ();
 b15zdnd11an1n08x5 FILLER_80_993 ();
 b15zdnd00an1n01x5 FILLER_80_1001 ();
 b15zdnd11an1n04x5 FILLER_80_1005 ();
 b15zdnd11an1n04x5 FILLER_80_1012 ();
 b15zdnd00an1n02x5 FILLER_80_1016 ();
 b15zdnd00an1n01x5 FILLER_80_1018 ();
 b15zdnd11an1n64x5 FILLER_80_1022 ();
 b15zdnd11an1n64x5 FILLER_80_1086 ();
 b15zdnd11an1n64x5 FILLER_80_1150 ();
 b15zdnd11an1n64x5 FILLER_80_1214 ();
 b15zdnd11an1n64x5 FILLER_80_1278 ();
 b15zdnd11an1n64x5 FILLER_80_1342 ();
 b15zdnd11an1n64x5 FILLER_80_1406 ();
 b15zdnd11an1n08x5 FILLER_80_1470 ();
 b15zdnd11an1n08x5 FILLER_80_2265 ();
 b15zdnd00an1n02x5 FILLER_80_2273 ();
 b15zdnd00an1n01x5 FILLER_80_2275 ();
 b15zdnd11an1n64x5 FILLER_81_0 ();
 b15zdnd11an1n64x5 FILLER_81_64 ();
 b15zdnd11an1n64x5 FILLER_81_128 ();
 b15zdnd11an1n64x5 FILLER_81_192 ();
 b15zdnd11an1n64x5 FILLER_81_256 ();
 b15zdnd11an1n64x5 FILLER_81_320 ();
 b15zdnd11an1n64x5 FILLER_81_384 ();
 b15zdnd11an1n64x5 FILLER_81_448 ();
 b15zdnd11an1n64x5 FILLER_81_512 ();
 b15zdnd11an1n64x5 FILLER_81_576 ();
 b15zdnd11an1n64x5 FILLER_81_640 ();
 b15zdnd11an1n32x5 FILLER_81_704 ();
 b15zdnd11an1n08x5 FILLER_81_736 ();
 b15zdnd11an1n04x5 FILLER_81_747 ();
 b15zdnd11an1n64x5 FILLER_81_754 ();
 b15zdnd11an1n64x5 FILLER_81_818 ();
 b15zdnd11an1n64x5 FILLER_81_882 ();
 b15zdnd11an1n32x5 FILLER_81_946 ();
 b15zdnd11an1n16x5 FILLER_81_978 ();
 b15zdnd11an1n08x5 FILLER_81_994 ();
 b15zdnd00an1n01x5 FILLER_81_1002 ();
 b15zdnd11an1n04x5 FILLER_81_1006 ();
 b15zdnd00an1n02x5 FILLER_81_1010 ();
 b15zdnd00an1n01x5 FILLER_81_1012 ();
 b15zdnd11an1n64x5 FILLER_81_1016 ();
 b15zdnd11an1n64x5 FILLER_81_1080 ();
 b15zdnd11an1n64x5 FILLER_81_1144 ();
 b15zdnd11an1n64x5 FILLER_81_1208 ();
 b15zdnd11an1n64x5 FILLER_81_1272 ();
 b15zdnd11an1n64x5 FILLER_81_1336 ();
 b15zdnd11an1n64x5 FILLER_81_1400 ();
 b15zdnd11an1n16x5 FILLER_81_1464 ();
 b15zdnd11an1n04x5 FILLER_81_1480 ();
 b15zdnd00an1n02x5 FILLER_81_1484 ();
 b15zdnd11an1n16x5 FILLER_81_2257 ();
 b15zdnd11an1n08x5 FILLER_81_2273 ();
 b15zdnd00an1n02x5 FILLER_81_2281 ();
 b15zdnd00an1n01x5 FILLER_81_2283 ();
 b15zdnd11an1n64x5 FILLER_82_8 ();
 b15zdnd11an1n64x5 FILLER_82_72 ();
 b15zdnd11an1n64x5 FILLER_82_136 ();
 b15zdnd11an1n64x5 FILLER_82_200 ();
 b15zdnd11an1n64x5 FILLER_82_264 ();
 b15zdnd11an1n64x5 FILLER_82_328 ();
 b15zdnd11an1n64x5 FILLER_82_392 ();
 b15zdnd11an1n64x5 FILLER_82_456 ();
 b15zdnd11an1n64x5 FILLER_82_520 ();
 b15zdnd11an1n64x5 FILLER_82_584 ();
 b15zdnd11an1n64x5 FILLER_82_648 ();
 b15zdnd11an1n04x5 FILLER_82_712 ();
 b15zdnd00an1n02x5 FILLER_82_716 ();
 b15zdnd00an1n02x5 FILLER_82_726 ();
 b15zdnd11an1n64x5 FILLER_82_772 ();
 b15zdnd11an1n64x5 FILLER_82_836 ();
 b15zdnd11an1n64x5 FILLER_82_900 ();
 b15zdnd11an1n16x5 FILLER_82_964 ();
 b15zdnd00an1n01x5 FILLER_82_980 ();
 b15zdnd11an1n64x5 FILLER_82_984 ();
 b15zdnd11an1n08x5 FILLER_82_1048 ();
 b15zdnd00an1n02x5 FILLER_82_1056 ();
 b15zdnd00an1n01x5 FILLER_82_1058 ();
 b15zdnd11an1n64x5 FILLER_82_1101 ();
 b15zdnd11an1n64x5 FILLER_82_1165 ();
 b15zdnd11an1n64x5 FILLER_82_1229 ();
 b15zdnd11an1n64x5 FILLER_82_1293 ();
 b15zdnd11an1n64x5 FILLER_82_1357 ();
 b15zdnd11an1n32x5 FILLER_82_1421 ();
 b15zdnd11an1n16x5 FILLER_82_1453 ();
 b15zdnd11an1n08x5 FILLER_82_1469 ();
 b15zdnd00an1n01x5 FILLER_82_1477 ();
 b15zdnd11an1n08x5 FILLER_82_2265 ();
 b15zdnd00an1n02x5 FILLER_82_2273 ();
 b15zdnd00an1n01x5 FILLER_82_2275 ();
 b15zdnd11an1n64x5 FILLER_83_0 ();
 b15zdnd11an1n64x5 FILLER_83_64 ();
 b15zdnd11an1n64x5 FILLER_83_128 ();
 b15zdnd11an1n64x5 FILLER_83_192 ();
 b15zdnd11an1n64x5 FILLER_83_256 ();
 b15zdnd11an1n64x5 FILLER_83_320 ();
 b15zdnd11an1n64x5 FILLER_83_384 ();
 b15zdnd11an1n64x5 FILLER_83_448 ();
 b15zdnd11an1n64x5 FILLER_83_512 ();
 b15zdnd11an1n64x5 FILLER_83_576 ();
 b15zdnd11an1n64x5 FILLER_83_640 ();
 b15zdnd00an1n01x5 FILLER_83_704 ();
 b15zdnd11an1n64x5 FILLER_83_749 ();
 b15zdnd11an1n64x5 FILLER_83_813 ();
 b15zdnd11an1n64x5 FILLER_83_877 ();
 b15zdnd11an1n16x5 FILLER_83_941 ();
 b15zdnd11an1n64x5 FILLER_83_1001 ();
 b15zdnd11an1n64x5 FILLER_83_1065 ();
 b15zdnd11an1n64x5 FILLER_83_1129 ();
 b15zdnd11an1n64x5 FILLER_83_1193 ();
 b15zdnd11an1n08x5 FILLER_83_1257 ();
 b15zdnd00an1n01x5 FILLER_83_1265 ();
 b15zdnd11an1n64x5 FILLER_83_1275 ();
 b15zdnd11an1n64x5 FILLER_83_1339 ();
 b15zdnd11an1n64x5 FILLER_83_1403 ();
 b15zdnd11an1n16x5 FILLER_83_1467 ();
 b15zdnd00an1n02x5 FILLER_83_1483 ();
 b15zdnd00an1n01x5 FILLER_83_1485 ();
 b15zdnd11an1n16x5 FILLER_83_2257 ();
 b15zdnd11an1n08x5 FILLER_83_2273 ();
 b15zdnd00an1n02x5 FILLER_83_2281 ();
 b15zdnd00an1n01x5 FILLER_83_2283 ();
 b15zdnd11an1n64x5 FILLER_84_8 ();
 b15zdnd11an1n64x5 FILLER_84_72 ();
 b15zdnd11an1n64x5 FILLER_84_136 ();
 b15zdnd11an1n64x5 FILLER_84_200 ();
 b15zdnd11an1n64x5 FILLER_84_264 ();
 b15zdnd11an1n64x5 FILLER_84_328 ();
 b15zdnd11an1n32x5 FILLER_84_392 ();
 b15zdnd11an1n64x5 FILLER_84_439 ();
 b15zdnd11an1n64x5 FILLER_84_503 ();
 b15zdnd11an1n64x5 FILLER_84_567 ();
 b15zdnd11an1n64x5 FILLER_84_631 ();
 b15zdnd11an1n16x5 FILLER_84_695 ();
 b15zdnd11an1n04x5 FILLER_84_711 ();
 b15zdnd00an1n02x5 FILLER_84_715 ();
 b15zdnd00an1n01x5 FILLER_84_717 ();
 b15zdnd00an1n02x5 FILLER_84_726 ();
 b15zdnd11an1n04x5 FILLER_84_731 ();
 b15zdnd11an1n04x5 FILLER_84_738 ();
 b15zdnd00an1n01x5 FILLER_84_742 ();
 b15zdnd11an1n64x5 FILLER_84_746 ();
 b15zdnd11an1n64x5 FILLER_84_810 ();
 b15zdnd11an1n64x5 FILLER_84_874 ();
 b15zdnd11an1n32x5 FILLER_84_938 ();
 b15zdnd00an1n02x5 FILLER_84_970 ();
 b15zdnd00an1n01x5 FILLER_84_972 ();
 b15zdnd11an1n04x5 FILLER_84_976 ();
 b15zdnd11an1n64x5 FILLER_84_983 ();
 b15zdnd11an1n64x5 FILLER_84_1047 ();
 b15zdnd11an1n64x5 FILLER_84_1111 ();
 b15zdnd11an1n64x5 FILLER_84_1175 ();
 b15zdnd11an1n32x5 FILLER_84_1239 ();
 b15zdnd11an1n16x5 FILLER_84_1271 ();
 b15zdnd11an1n04x5 FILLER_84_1287 ();
 b15zdnd00an1n02x5 FILLER_84_1291 ();
 b15zdnd00an1n01x5 FILLER_84_1293 ();
 b15zdnd11an1n64x5 FILLER_84_1297 ();
 b15zdnd11an1n64x5 FILLER_84_1361 ();
 b15zdnd11an1n32x5 FILLER_84_1425 ();
 b15zdnd11an1n16x5 FILLER_84_1457 ();
 b15zdnd11an1n04x5 FILLER_84_1473 ();
 b15zdnd00an1n01x5 FILLER_84_1477 ();
 b15zdnd11an1n08x5 FILLER_84_2265 ();
 b15zdnd00an1n02x5 FILLER_84_2273 ();
 b15zdnd00an1n01x5 FILLER_84_2275 ();
 b15zdnd11an1n64x5 FILLER_85_0 ();
 b15zdnd11an1n64x5 FILLER_85_64 ();
 b15zdnd11an1n64x5 FILLER_85_128 ();
 b15zdnd11an1n64x5 FILLER_85_192 ();
 b15zdnd11an1n64x5 FILLER_85_256 ();
 b15zdnd11an1n64x5 FILLER_85_320 ();
 b15zdnd11an1n64x5 FILLER_85_384 ();
 b15zdnd11an1n64x5 FILLER_85_448 ();
 b15zdnd11an1n64x5 FILLER_85_512 ();
 b15zdnd11an1n64x5 FILLER_85_576 ();
 b15zdnd11an1n64x5 FILLER_85_640 ();
 b15zdnd11an1n64x5 FILLER_85_748 ();
 b15zdnd11an1n64x5 FILLER_85_812 ();
 b15zdnd11an1n64x5 FILLER_85_876 ();
 b15zdnd11an1n64x5 FILLER_85_940 ();
 b15zdnd11an1n64x5 FILLER_85_1004 ();
 b15zdnd11an1n64x5 FILLER_85_1068 ();
 b15zdnd11an1n64x5 FILLER_85_1132 ();
 b15zdnd11an1n64x5 FILLER_85_1196 ();
 b15zdnd11an1n16x5 FILLER_85_1260 ();
 b15zdnd11an1n08x5 FILLER_85_1276 ();
 b15zdnd00an1n02x5 FILLER_85_1284 ();
 b15zdnd11an1n04x5 FILLER_85_1289 ();
 b15zdnd11an1n04x5 FILLER_85_1296 ();
 b15zdnd11an1n64x5 FILLER_85_1303 ();
 b15zdnd11an1n64x5 FILLER_85_1367 ();
 b15zdnd11an1n32x5 FILLER_85_1431 ();
 b15zdnd11an1n16x5 FILLER_85_1463 ();
 b15zdnd11an1n04x5 FILLER_85_1479 ();
 b15zdnd00an1n02x5 FILLER_85_1483 ();
 b15zdnd00an1n01x5 FILLER_85_1485 ();
 b15zdnd11an1n16x5 FILLER_85_2257 ();
 b15zdnd11an1n08x5 FILLER_85_2273 ();
 b15zdnd00an1n02x5 FILLER_85_2281 ();
 b15zdnd00an1n01x5 FILLER_85_2283 ();
 b15zdnd11an1n64x5 FILLER_86_8 ();
 b15zdnd11an1n64x5 FILLER_86_72 ();
 b15zdnd11an1n64x5 FILLER_86_136 ();
 b15zdnd11an1n64x5 FILLER_86_200 ();
 b15zdnd11an1n64x5 FILLER_86_264 ();
 b15zdnd11an1n64x5 FILLER_86_328 ();
 b15zdnd11an1n64x5 FILLER_86_392 ();
 b15zdnd11an1n64x5 FILLER_86_456 ();
 b15zdnd11an1n64x5 FILLER_86_520 ();
 b15zdnd11an1n64x5 FILLER_86_584 ();
 b15zdnd11an1n64x5 FILLER_86_648 ();
 b15zdnd00an1n01x5 FILLER_86_712 ();
 b15zdnd00an1n02x5 FILLER_86_716 ();
 b15zdnd00an1n02x5 FILLER_86_726 ();
 b15zdnd11an1n04x5 FILLER_86_731 ();
 b15zdnd11an1n08x5 FILLER_86_738 ();
 b15zdnd11an1n64x5 FILLER_86_749 ();
 b15zdnd11an1n64x5 FILLER_86_813 ();
 b15zdnd11an1n64x5 FILLER_86_877 ();
 b15zdnd11an1n64x5 FILLER_86_941 ();
 b15zdnd11an1n64x5 FILLER_86_1005 ();
 b15zdnd11an1n64x5 FILLER_86_1069 ();
 b15zdnd11an1n64x5 FILLER_86_1133 ();
 b15zdnd11an1n64x5 FILLER_86_1197 ();
 b15zdnd11an1n08x5 FILLER_86_1261 ();
 b15zdnd11an1n04x5 FILLER_86_1269 ();
 b15zdnd00an1n01x5 FILLER_86_1273 ();
 b15zdnd11an1n04x5 FILLER_86_1318 ();
 b15zdnd11an1n64x5 FILLER_86_1325 ();
 b15zdnd11an1n64x5 FILLER_86_1389 ();
 b15zdnd11an1n16x5 FILLER_86_1453 ();
 b15zdnd11an1n08x5 FILLER_86_1469 ();
 b15zdnd00an1n01x5 FILLER_86_1477 ();
 b15zdnd11an1n08x5 FILLER_86_2265 ();
 b15zdnd00an1n02x5 FILLER_86_2273 ();
 b15zdnd00an1n01x5 FILLER_86_2275 ();
 b15zdnd11an1n64x5 FILLER_87_0 ();
 b15zdnd11an1n64x5 FILLER_87_64 ();
 b15zdnd11an1n64x5 FILLER_87_128 ();
 b15zdnd11an1n64x5 FILLER_87_192 ();
 b15zdnd11an1n64x5 FILLER_87_256 ();
 b15zdnd11an1n64x5 FILLER_87_320 ();
 b15zdnd11an1n64x5 FILLER_87_384 ();
 b15zdnd11an1n64x5 FILLER_87_448 ();
 b15zdnd11an1n64x5 FILLER_87_512 ();
 b15zdnd11an1n64x5 FILLER_87_576 ();
 b15zdnd11an1n64x5 FILLER_87_640 ();
 b15zdnd11an1n04x5 FILLER_87_704 ();
 b15zdnd11an1n64x5 FILLER_87_752 ();
 b15zdnd11an1n64x5 FILLER_87_816 ();
 b15zdnd11an1n64x5 FILLER_87_880 ();
 b15zdnd11an1n64x5 FILLER_87_944 ();
 b15zdnd11an1n64x5 FILLER_87_1008 ();
 b15zdnd11an1n64x5 FILLER_87_1072 ();
 b15zdnd11an1n64x5 FILLER_87_1136 ();
 b15zdnd11an1n64x5 FILLER_87_1200 ();
 b15zdnd11an1n08x5 FILLER_87_1264 ();
 b15zdnd00an1n02x5 FILLER_87_1272 ();
 b15zdnd11an1n04x5 FILLER_87_1318 ();
 b15zdnd11an1n04x5 FILLER_87_1325 ();
 b15zdnd11an1n64x5 FILLER_87_1332 ();
 b15zdnd11an1n64x5 FILLER_87_1396 ();
 b15zdnd11an1n16x5 FILLER_87_1460 ();
 b15zdnd11an1n08x5 FILLER_87_1476 ();
 b15zdnd00an1n02x5 FILLER_87_1484 ();
 b15zdnd11an1n16x5 FILLER_87_2257 ();
 b15zdnd11an1n08x5 FILLER_87_2273 ();
 b15zdnd00an1n02x5 FILLER_87_2281 ();
 b15zdnd00an1n01x5 FILLER_87_2283 ();
 b15zdnd11an1n64x5 FILLER_88_8 ();
 b15zdnd11an1n64x5 FILLER_88_72 ();
 b15zdnd11an1n64x5 FILLER_88_136 ();
 b15zdnd11an1n64x5 FILLER_88_200 ();
 b15zdnd11an1n64x5 FILLER_88_264 ();
 b15zdnd11an1n64x5 FILLER_88_328 ();
 b15zdnd11an1n16x5 FILLER_88_392 ();
 b15zdnd11an1n08x5 FILLER_88_408 ();
 b15zdnd11an1n04x5 FILLER_88_416 ();
 b15zdnd11an1n64x5 FILLER_88_433 ();
 b15zdnd11an1n64x5 FILLER_88_497 ();
 b15zdnd11an1n64x5 FILLER_88_561 ();
 b15zdnd11an1n64x5 FILLER_88_625 ();
 b15zdnd11an1n16x5 FILLER_88_689 ();
 b15zdnd11an1n08x5 FILLER_88_705 ();
 b15zdnd11an1n04x5 FILLER_88_713 ();
 b15zdnd00an1n01x5 FILLER_88_717 ();
 b15zdnd11an1n04x5 FILLER_88_726 ();
 b15zdnd00an1n01x5 FILLER_88_730 ();
 b15zdnd11an1n64x5 FILLER_88_734 ();
 b15zdnd11an1n64x5 FILLER_88_798 ();
 b15zdnd11an1n64x5 FILLER_88_862 ();
 b15zdnd11an1n64x5 FILLER_88_926 ();
 b15zdnd11an1n64x5 FILLER_88_990 ();
 b15zdnd11an1n64x5 FILLER_88_1054 ();
 b15zdnd11an1n64x5 FILLER_88_1118 ();
 b15zdnd11an1n64x5 FILLER_88_1182 ();
 b15zdnd11an1n16x5 FILLER_88_1246 ();
 b15zdnd11an1n04x5 FILLER_88_1262 ();
 b15zdnd00an1n01x5 FILLER_88_1266 ();
 b15zdnd11an1n04x5 FILLER_88_1270 ();
 b15zdnd11an1n04x5 FILLER_88_1318 ();
 b15zdnd11an1n04x5 FILLER_88_1325 ();
 b15zdnd11an1n64x5 FILLER_88_1332 ();
 b15zdnd11an1n64x5 FILLER_88_1396 ();
 b15zdnd11an1n16x5 FILLER_88_1460 ();
 b15zdnd00an1n02x5 FILLER_88_1476 ();
 b15zdnd11an1n08x5 FILLER_88_2265 ();
 b15zdnd00an1n02x5 FILLER_88_2273 ();
 b15zdnd00an1n01x5 FILLER_88_2275 ();
 b15zdnd11an1n64x5 FILLER_89_0 ();
 b15zdnd11an1n64x5 FILLER_89_64 ();
 b15zdnd11an1n64x5 FILLER_89_128 ();
 b15zdnd11an1n64x5 FILLER_89_192 ();
 b15zdnd11an1n64x5 FILLER_89_256 ();
 b15zdnd11an1n64x5 FILLER_89_320 ();
 b15zdnd11an1n32x5 FILLER_89_384 ();
 b15zdnd00an1n02x5 FILLER_89_416 ();
 b15zdnd00an1n01x5 FILLER_89_418 ();
 b15zdnd11an1n64x5 FILLER_89_435 ();
 b15zdnd11an1n64x5 FILLER_89_499 ();
 b15zdnd11an1n64x5 FILLER_89_563 ();
 b15zdnd11an1n64x5 FILLER_89_627 ();
 b15zdnd11an1n32x5 FILLER_89_691 ();
 b15zdnd11an1n04x5 FILLER_89_723 ();
 b15zdnd00an1n02x5 FILLER_89_727 ();
 b15zdnd11an1n64x5 FILLER_89_732 ();
 b15zdnd11an1n64x5 FILLER_89_796 ();
 b15zdnd11an1n64x5 FILLER_89_860 ();
 b15zdnd11an1n64x5 FILLER_89_924 ();
 b15zdnd11an1n64x5 FILLER_89_988 ();
 b15zdnd11an1n64x5 FILLER_89_1052 ();
 b15zdnd11an1n64x5 FILLER_89_1116 ();
 b15zdnd11an1n64x5 FILLER_89_1180 ();
 b15zdnd11an1n16x5 FILLER_89_1244 ();
 b15zdnd11an1n08x5 FILLER_89_1260 ();
 b15zdnd11an1n04x5 FILLER_89_1268 ();
 b15zdnd00an1n02x5 FILLER_89_1272 ();
 b15zdnd11an1n04x5 FILLER_89_1318 ();
 b15zdnd11an1n04x5 FILLER_89_1325 ();
 b15zdnd11an1n64x5 FILLER_89_1332 ();
 b15zdnd11an1n64x5 FILLER_89_1396 ();
 b15zdnd11an1n16x5 FILLER_89_1460 ();
 b15zdnd11an1n08x5 FILLER_89_1476 ();
 b15zdnd00an1n02x5 FILLER_89_1484 ();
 b15zdnd11an1n16x5 FILLER_89_2257 ();
 b15zdnd11an1n08x5 FILLER_89_2273 ();
 b15zdnd00an1n02x5 FILLER_89_2281 ();
 b15zdnd00an1n01x5 FILLER_89_2283 ();
 b15zdnd11an1n64x5 FILLER_90_8 ();
 b15zdnd11an1n64x5 FILLER_90_72 ();
 b15zdnd11an1n64x5 FILLER_90_136 ();
 b15zdnd11an1n64x5 FILLER_90_200 ();
 b15zdnd11an1n64x5 FILLER_90_264 ();
 b15zdnd11an1n64x5 FILLER_90_328 ();
 b15zdnd11an1n64x5 FILLER_90_392 ();
 b15zdnd11an1n64x5 FILLER_90_456 ();
 b15zdnd11an1n64x5 FILLER_90_520 ();
 b15zdnd11an1n64x5 FILLER_90_584 ();
 b15zdnd11an1n64x5 FILLER_90_648 ();
 b15zdnd11an1n04x5 FILLER_90_712 ();
 b15zdnd00an1n02x5 FILLER_90_716 ();
 b15zdnd11an1n64x5 FILLER_90_726 ();
 b15zdnd11an1n64x5 FILLER_90_790 ();
 b15zdnd11an1n64x5 FILLER_90_854 ();
 b15zdnd11an1n64x5 FILLER_90_918 ();
 b15zdnd11an1n64x5 FILLER_90_982 ();
 b15zdnd11an1n64x5 FILLER_90_1046 ();
 b15zdnd11an1n64x5 FILLER_90_1110 ();
 b15zdnd11an1n64x5 FILLER_90_1174 ();
 b15zdnd11an1n32x5 FILLER_90_1238 ();
 b15zdnd11an1n16x5 FILLER_90_1270 ();
 b15zdnd11an1n04x5 FILLER_90_1289 ();
 b15zdnd11an1n04x5 FILLER_90_1296 ();
 b15zdnd11an1n04x5 FILLER_90_1303 ();
 b15zdnd11an1n04x5 FILLER_90_1310 ();
 b15zdnd11an1n64x5 FILLER_90_1317 ();
 b15zdnd11an1n64x5 FILLER_90_1381 ();
 b15zdnd11an1n32x5 FILLER_90_1445 ();
 b15zdnd00an1n01x5 FILLER_90_1477 ();
 b15zdnd11an1n08x5 FILLER_90_2265 ();
 b15zdnd00an1n02x5 FILLER_90_2273 ();
 b15zdnd00an1n01x5 FILLER_90_2275 ();
 b15zdnd00an1n02x5 FILLER_91_0 ();
 b15zdnd00an1n01x5 FILLER_91_2 ();
 b15zdnd11an1n08x5 FILLER_91_10 ();
 b15zdnd11an1n04x5 FILLER_91_25 ();
 b15zdnd11an1n04x5 FILLER_91_33 ();
 b15zdnd11an1n64x5 FILLER_91_41 ();
 b15zdnd11an1n64x5 FILLER_91_105 ();
 b15zdnd11an1n64x5 FILLER_91_169 ();
 b15zdnd11an1n64x5 FILLER_91_233 ();
 b15zdnd11an1n64x5 FILLER_91_297 ();
 b15zdnd11an1n64x5 FILLER_91_361 ();
 b15zdnd11an1n64x5 FILLER_91_425 ();
 b15zdnd11an1n64x5 FILLER_91_489 ();
 b15zdnd11an1n64x5 FILLER_91_553 ();
 b15zdnd11an1n64x5 FILLER_91_617 ();
 b15zdnd11an1n64x5 FILLER_91_681 ();
 b15zdnd11an1n64x5 FILLER_91_745 ();
 b15zdnd11an1n64x5 FILLER_91_809 ();
 b15zdnd11an1n64x5 FILLER_91_873 ();
 b15zdnd11an1n64x5 FILLER_91_937 ();
 b15zdnd11an1n64x5 FILLER_91_1001 ();
 b15zdnd11an1n64x5 FILLER_91_1065 ();
 b15zdnd11an1n64x5 FILLER_91_1129 ();
 b15zdnd11an1n32x5 FILLER_91_1193 ();
 b15zdnd11an1n16x5 FILLER_91_1225 ();
 b15zdnd11an1n08x5 FILLER_91_1241 ();
 b15zdnd00an1n02x5 FILLER_91_1249 ();
 b15zdnd11an1n16x5 FILLER_91_1258 ();
 b15zdnd11an1n08x5 FILLER_91_1274 ();
 b15zdnd00an1n02x5 FILLER_91_1282 ();
 b15zdnd11an1n04x5 FILLER_91_1293 ();
 b15zdnd11an1n04x5 FILLER_91_1300 ();
 b15zdnd11an1n64x5 FILLER_91_1307 ();
 b15zdnd11an1n64x5 FILLER_91_1371 ();
 b15zdnd11an1n32x5 FILLER_91_1435 ();
 b15zdnd11an1n16x5 FILLER_91_1467 ();
 b15zdnd00an1n02x5 FILLER_91_1483 ();
 b15zdnd00an1n01x5 FILLER_91_1485 ();
 b15zdnd11an1n16x5 FILLER_91_2257 ();
 b15zdnd11an1n08x5 FILLER_91_2273 ();
 b15zdnd00an1n02x5 FILLER_91_2281 ();
 b15zdnd00an1n01x5 FILLER_91_2283 ();
 b15zdnd00an1n02x5 FILLER_92_8 ();
 b15zdnd00an1n01x5 FILLER_92_10 ();
 b15zdnd11an1n64x5 FILLER_92_53 ();
 b15zdnd11an1n64x5 FILLER_92_117 ();
 b15zdnd11an1n64x5 FILLER_92_181 ();
 b15zdnd11an1n64x5 FILLER_92_245 ();
 b15zdnd11an1n64x5 FILLER_92_309 ();
 b15zdnd11an1n32x5 FILLER_92_373 ();
 b15zdnd11an1n08x5 FILLER_92_405 ();
 b15zdnd00an1n02x5 FILLER_92_413 ();
 b15zdnd11an1n64x5 FILLER_92_427 ();
 b15zdnd11an1n64x5 FILLER_92_491 ();
 b15zdnd11an1n64x5 FILLER_92_555 ();
 b15zdnd11an1n64x5 FILLER_92_619 ();
 b15zdnd11an1n32x5 FILLER_92_683 ();
 b15zdnd00an1n02x5 FILLER_92_715 ();
 b15zdnd00an1n01x5 FILLER_92_717 ();
 b15zdnd00an1n02x5 FILLER_92_726 ();
 b15zdnd11an1n16x5 FILLER_92_772 ();
 b15zdnd11an1n04x5 FILLER_92_788 ();
 b15zdnd00an1n02x5 FILLER_92_792 ();
 b15zdnd11an1n64x5 FILLER_92_803 ();
 b15zdnd11an1n64x5 FILLER_92_867 ();
 b15zdnd11an1n64x5 FILLER_92_931 ();
 b15zdnd11an1n64x5 FILLER_92_995 ();
 b15zdnd11an1n64x5 FILLER_92_1059 ();
 b15zdnd11an1n64x5 FILLER_92_1123 ();
 b15zdnd11an1n64x5 FILLER_92_1187 ();
 b15zdnd11an1n08x5 FILLER_92_1251 ();
 b15zdnd11an1n04x5 FILLER_92_1259 ();
 b15zdnd00an1n02x5 FILLER_92_1263 ();
 b15zdnd00an1n01x5 FILLER_92_1265 ();
 b15zdnd11an1n16x5 FILLER_92_1275 ();
 b15zdnd11an1n04x5 FILLER_92_1291 ();
 b15zdnd00an1n01x5 FILLER_92_1295 ();
 b15zdnd11an1n04x5 FILLER_92_1299 ();
 b15zdnd11an1n64x5 FILLER_92_1306 ();
 b15zdnd11an1n64x5 FILLER_92_1370 ();
 b15zdnd11an1n08x5 FILLER_92_1434 ();
 b15zdnd11an1n04x5 FILLER_92_1442 ();
 b15zdnd11an1n16x5 FILLER_92_1460 ();
 b15zdnd00an1n02x5 FILLER_92_1476 ();
 b15zdnd11an1n08x5 FILLER_92_2265 ();
 b15zdnd00an1n02x5 FILLER_92_2273 ();
 b15zdnd00an1n01x5 FILLER_92_2275 ();
 b15zdnd11an1n08x5 FILLER_93_0 ();
 b15zdnd00an1n01x5 FILLER_93_8 ();
 b15zdnd11an1n64x5 FILLER_93_51 ();
 b15zdnd11an1n64x5 FILLER_93_115 ();
 b15zdnd11an1n64x5 FILLER_93_179 ();
 b15zdnd11an1n64x5 FILLER_93_243 ();
 b15zdnd11an1n64x5 FILLER_93_307 ();
 b15zdnd11an1n64x5 FILLER_93_371 ();
 b15zdnd11an1n64x5 FILLER_93_435 ();
 b15zdnd11an1n64x5 FILLER_93_499 ();
 b15zdnd11an1n64x5 FILLER_93_563 ();
 b15zdnd11an1n64x5 FILLER_93_627 ();
 b15zdnd11an1n16x5 FILLER_93_691 ();
 b15zdnd11an1n08x5 FILLER_93_707 ();
 b15zdnd11an1n04x5 FILLER_93_715 ();
 b15zdnd00an1n02x5 FILLER_93_719 ();
 b15zdnd11an1n64x5 FILLER_93_724 ();
 b15zdnd11an1n64x5 FILLER_93_788 ();
 b15zdnd11an1n64x5 FILLER_93_852 ();
 b15zdnd11an1n64x5 FILLER_93_916 ();
 b15zdnd11an1n64x5 FILLER_93_980 ();
 b15zdnd11an1n64x5 FILLER_93_1044 ();
 b15zdnd11an1n64x5 FILLER_93_1108 ();
 b15zdnd11an1n64x5 FILLER_93_1172 ();
 b15zdnd11an1n32x5 FILLER_93_1236 ();
 b15zdnd11an1n08x5 FILLER_93_1268 ();
 b15zdnd00an1n02x5 FILLER_93_1276 ();
 b15zdnd00an1n01x5 FILLER_93_1278 ();
 b15zdnd11an1n64x5 FILLER_93_1323 ();
 b15zdnd11an1n64x5 FILLER_93_1387 ();
 b15zdnd11an1n32x5 FILLER_93_1451 ();
 b15zdnd00an1n02x5 FILLER_93_1483 ();
 b15zdnd00an1n01x5 FILLER_93_1485 ();
 b15zdnd11an1n16x5 FILLER_93_2257 ();
 b15zdnd11an1n08x5 FILLER_93_2273 ();
 b15zdnd00an1n02x5 FILLER_93_2281 ();
 b15zdnd00an1n01x5 FILLER_93_2283 ();
 b15zdnd00an1n02x5 FILLER_94_8 ();
 b15zdnd00an1n01x5 FILLER_94_10 ();
 b15zdnd11an1n04x5 FILLER_94_18 ();
 b15zdnd11an1n04x5 FILLER_94_29 ();
 b15zdnd11an1n64x5 FILLER_94_37 ();
 b15zdnd11an1n64x5 FILLER_94_101 ();
 b15zdnd11an1n64x5 FILLER_94_165 ();
 b15zdnd11an1n64x5 FILLER_94_229 ();
 b15zdnd11an1n64x5 FILLER_94_293 ();
 b15zdnd11an1n32x5 FILLER_94_357 ();
 b15zdnd11an1n16x5 FILLER_94_389 ();
 b15zdnd11an1n08x5 FILLER_94_405 ();
 b15zdnd00an1n02x5 FILLER_94_413 ();
 b15zdnd00an1n01x5 FILLER_94_415 ();
 b15zdnd11an1n64x5 FILLER_94_423 ();
 b15zdnd11an1n64x5 FILLER_94_487 ();
 b15zdnd11an1n64x5 FILLER_94_551 ();
 b15zdnd11an1n16x5 FILLER_94_615 ();
 b15zdnd11an1n32x5 FILLER_94_673 ();
 b15zdnd11an1n08x5 FILLER_94_705 ();
 b15zdnd11an1n04x5 FILLER_94_713 ();
 b15zdnd00an1n01x5 FILLER_94_717 ();
 b15zdnd00an1n02x5 FILLER_94_726 ();
 b15zdnd11an1n64x5 FILLER_94_731 ();
 b15zdnd11an1n64x5 FILLER_94_795 ();
 b15zdnd11an1n64x5 FILLER_94_859 ();
 b15zdnd11an1n64x5 FILLER_94_923 ();
 b15zdnd11an1n64x5 FILLER_94_987 ();
 b15zdnd11an1n64x5 FILLER_94_1051 ();
 b15zdnd11an1n64x5 FILLER_94_1115 ();
 b15zdnd11an1n64x5 FILLER_94_1179 ();
 b15zdnd11an1n32x5 FILLER_94_1243 ();
 b15zdnd11an1n04x5 FILLER_94_1275 ();
 b15zdnd11an1n04x5 FILLER_94_1323 ();
 b15zdnd11an1n64x5 FILLER_94_1330 ();
 b15zdnd11an1n64x5 FILLER_94_1394 ();
 b15zdnd11an1n16x5 FILLER_94_1458 ();
 b15zdnd11an1n04x5 FILLER_94_1474 ();
 b15zdnd11an1n08x5 FILLER_94_2265 ();
 b15zdnd00an1n02x5 FILLER_94_2273 ();
 b15zdnd00an1n01x5 FILLER_94_2275 ();
 b15zdnd11an1n08x5 FILLER_95_0 ();
 b15zdnd11an1n04x5 FILLER_95_8 ();
 b15zdnd11an1n64x5 FILLER_95_54 ();
 b15zdnd11an1n64x5 FILLER_95_118 ();
 b15zdnd11an1n64x5 FILLER_95_182 ();
 b15zdnd11an1n64x5 FILLER_95_246 ();
 b15zdnd11an1n64x5 FILLER_95_310 ();
 b15zdnd11an1n32x5 FILLER_95_374 ();
 b15zdnd11an1n08x5 FILLER_95_406 ();
 b15zdnd11an1n04x5 FILLER_95_414 ();
 b15zdnd00an1n01x5 FILLER_95_418 ();
 b15zdnd11an1n64x5 FILLER_95_423 ();
 b15zdnd11an1n64x5 FILLER_95_487 ();
 b15zdnd11an1n64x5 FILLER_95_551 ();
 b15zdnd11an1n16x5 FILLER_95_615 ();
 b15zdnd11an1n08x5 FILLER_95_631 ();
 b15zdnd00an1n01x5 FILLER_95_639 ();
 b15zdnd11an1n08x5 FILLER_95_682 ();
 b15zdnd00an1n02x5 FILLER_95_690 ();
 b15zdnd11an1n64x5 FILLER_95_734 ();
 b15zdnd11an1n64x5 FILLER_95_798 ();
 b15zdnd11an1n64x5 FILLER_95_862 ();
 b15zdnd11an1n64x5 FILLER_95_926 ();
 b15zdnd11an1n64x5 FILLER_95_990 ();
 b15zdnd11an1n64x5 FILLER_95_1054 ();
 b15zdnd11an1n64x5 FILLER_95_1118 ();
 b15zdnd11an1n64x5 FILLER_95_1182 ();
 b15zdnd11an1n32x5 FILLER_95_1246 ();
 b15zdnd00an1n02x5 FILLER_95_1278 ();
 b15zdnd00an1n01x5 FILLER_95_1280 ();
 b15zdnd11an1n64x5 FILLER_95_1325 ();
 b15zdnd11an1n64x5 FILLER_95_1389 ();
 b15zdnd11an1n32x5 FILLER_95_1453 ();
 b15zdnd00an1n01x5 FILLER_95_1485 ();
 b15zdnd00an1n02x5 FILLER_95_2257 ();
 b15zdnd11an1n08x5 FILLER_95_2262 ();
 b15zdnd00an1n01x5 FILLER_95_2270 ();
 b15zdnd00an1n02x5 FILLER_95_2282 ();
 b15zdnd00an1n02x5 FILLER_96_8 ();
 b15zdnd11an1n64x5 FILLER_96_52 ();
 b15zdnd11an1n64x5 FILLER_96_116 ();
 b15zdnd11an1n64x5 FILLER_96_180 ();
 b15zdnd11an1n64x5 FILLER_96_244 ();
 b15zdnd11an1n64x5 FILLER_96_308 ();
 b15zdnd11an1n32x5 FILLER_96_372 ();
 b15zdnd11an1n08x5 FILLER_96_404 ();
 b15zdnd00an1n02x5 FILLER_96_412 ();
 b15zdnd00an1n01x5 FILLER_96_414 ();
 b15zdnd11an1n04x5 FILLER_96_419 ();
 b15zdnd00an1n01x5 FILLER_96_423 ();
 b15zdnd11an1n64x5 FILLER_96_427 ();
 b15zdnd11an1n64x5 FILLER_96_491 ();
 b15zdnd11an1n64x5 FILLER_96_555 ();
 b15zdnd11an1n04x5 FILLER_96_619 ();
 b15zdnd00an1n02x5 FILLER_96_623 ();
 b15zdnd11an1n32x5 FILLER_96_667 ();
 b15zdnd11an1n16x5 FILLER_96_699 ();
 b15zdnd00an1n02x5 FILLER_96_715 ();
 b15zdnd00an1n01x5 FILLER_96_717 ();
 b15zdnd00an1n02x5 FILLER_96_726 ();
 b15zdnd11an1n64x5 FILLER_96_731 ();
 b15zdnd11an1n64x5 FILLER_96_795 ();
 b15zdnd11an1n64x5 FILLER_96_859 ();
 b15zdnd11an1n64x5 FILLER_96_923 ();
 b15zdnd11an1n64x5 FILLER_96_987 ();
 b15zdnd11an1n64x5 FILLER_96_1051 ();
 b15zdnd11an1n64x5 FILLER_96_1115 ();
 b15zdnd11an1n64x5 FILLER_96_1179 ();
 b15zdnd11an1n32x5 FILLER_96_1243 ();
 b15zdnd11an1n16x5 FILLER_96_1275 ();
 b15zdnd11an1n04x5 FILLER_96_1291 ();
 b15zdnd00an1n01x5 FILLER_96_1295 ();
 b15zdnd11an1n04x5 FILLER_96_1299 ();
 b15zdnd11an1n04x5 FILLER_96_1306 ();
 b15zdnd11an1n04x5 FILLER_96_1313 ();
 b15zdnd11an1n64x5 FILLER_96_1320 ();
 b15zdnd11an1n64x5 FILLER_96_1384 ();
 b15zdnd11an1n16x5 FILLER_96_1448 ();
 b15zdnd11an1n08x5 FILLER_96_1464 ();
 b15zdnd11an1n04x5 FILLER_96_1472 ();
 b15zdnd00an1n02x5 FILLER_96_1476 ();
 b15zdnd00an1n02x5 FILLER_96_2265 ();
 b15zdnd11an1n04x5 FILLER_96_2270 ();
 b15zdnd00an1n02x5 FILLER_96_2274 ();
 b15zdnd11an1n16x5 FILLER_97_0 ();
 b15zdnd00an1n01x5 FILLER_97_16 ();
 b15zdnd11an1n64x5 FILLER_97_21 ();
 b15zdnd11an1n64x5 FILLER_97_85 ();
 b15zdnd11an1n64x5 FILLER_97_149 ();
 b15zdnd11an1n64x5 FILLER_97_213 ();
 b15zdnd11an1n64x5 FILLER_97_277 ();
 b15zdnd11an1n64x5 FILLER_97_341 ();
 b15zdnd11an1n08x5 FILLER_97_405 ();
 b15zdnd00an1n02x5 FILLER_97_413 ();
 b15zdnd11an1n64x5 FILLER_97_422 ();
 b15zdnd11an1n64x5 FILLER_97_486 ();
 b15zdnd11an1n64x5 FILLER_97_550 ();
 b15zdnd11an1n64x5 FILLER_97_614 ();
 b15zdnd11an1n08x5 FILLER_97_678 ();
 b15zdnd00an1n02x5 FILLER_97_686 ();
 b15zdnd11an1n64x5 FILLER_97_730 ();
 b15zdnd11an1n64x5 FILLER_97_794 ();
 b15zdnd11an1n32x5 FILLER_97_858 ();
 b15zdnd11an1n08x5 FILLER_97_890 ();
 b15zdnd11an1n04x5 FILLER_97_898 ();
 b15zdnd00an1n02x5 FILLER_97_902 ();
 b15zdnd00an1n01x5 FILLER_97_904 ();
 b15zdnd11an1n64x5 FILLER_97_914 ();
 b15zdnd11an1n64x5 FILLER_97_978 ();
 b15zdnd11an1n64x5 FILLER_97_1042 ();
 b15zdnd11an1n64x5 FILLER_97_1106 ();
 b15zdnd11an1n64x5 FILLER_97_1170 ();
 b15zdnd11an1n64x5 FILLER_97_1234 ();
 b15zdnd00an1n02x5 FILLER_97_1298 ();
 b15zdnd00an1n01x5 FILLER_97_1300 ();
 b15zdnd11an1n04x5 FILLER_97_1304 ();
 b15zdnd11an1n64x5 FILLER_97_1311 ();
 b15zdnd11an1n64x5 FILLER_97_1375 ();
 b15zdnd11an1n32x5 FILLER_97_1439 ();
 b15zdnd11an1n08x5 FILLER_97_1471 ();
 b15zdnd11an1n04x5 FILLER_97_1479 ();
 b15zdnd00an1n02x5 FILLER_97_1483 ();
 b15zdnd00an1n01x5 FILLER_97_1485 ();
 b15zdnd00an1n02x5 FILLER_97_2257 ();
 b15zdnd11an1n04x5 FILLER_97_2262 ();
 b15zdnd11an1n08x5 FILLER_97_2269 ();
 b15zdnd11an1n04x5 FILLER_97_2277 ();
 b15zdnd00an1n02x5 FILLER_97_2281 ();
 b15zdnd00an1n01x5 FILLER_97_2283 ();
 b15zdnd11an1n64x5 FILLER_98_8 ();
 b15zdnd11an1n64x5 FILLER_98_72 ();
 b15zdnd11an1n64x5 FILLER_98_136 ();
 b15zdnd11an1n64x5 FILLER_98_200 ();
 b15zdnd11an1n64x5 FILLER_98_264 ();
 b15zdnd11an1n64x5 FILLER_98_328 ();
 b15zdnd11an1n64x5 FILLER_98_392 ();
 b15zdnd11an1n64x5 FILLER_98_456 ();
 b15zdnd11an1n64x5 FILLER_98_520 ();
 b15zdnd11an1n64x5 FILLER_98_584 ();
 b15zdnd11an1n64x5 FILLER_98_648 ();
 b15zdnd11an1n04x5 FILLER_98_712 ();
 b15zdnd00an1n02x5 FILLER_98_716 ();
 b15zdnd11an1n64x5 FILLER_98_726 ();
 b15zdnd11an1n64x5 FILLER_98_790 ();
 b15zdnd11an1n64x5 FILLER_98_854 ();
 b15zdnd11an1n64x5 FILLER_98_918 ();
 b15zdnd11an1n64x5 FILLER_98_982 ();
 b15zdnd11an1n64x5 FILLER_98_1046 ();
 b15zdnd11an1n64x5 FILLER_98_1110 ();
 b15zdnd11an1n64x5 FILLER_98_1174 ();
 b15zdnd11an1n64x5 FILLER_98_1238 ();
 b15zdnd11an1n64x5 FILLER_98_1305 ();
 b15zdnd11an1n64x5 FILLER_98_1369 ();
 b15zdnd11an1n32x5 FILLER_98_1433 ();
 b15zdnd11an1n08x5 FILLER_98_1465 ();
 b15zdnd11an1n04x5 FILLER_98_1473 ();
 b15zdnd00an1n01x5 FILLER_98_1477 ();
 b15zdnd00an1n02x5 FILLER_98_2265 ();
 b15zdnd00an1n01x5 FILLER_98_2267 ();
 b15zdnd00an1n02x5 FILLER_98_2274 ();
 b15zdnd11an1n64x5 FILLER_99_0 ();
 b15zdnd11an1n64x5 FILLER_99_64 ();
 b15zdnd11an1n64x5 FILLER_99_128 ();
 b15zdnd11an1n32x5 FILLER_99_192 ();
 b15zdnd11an1n16x5 FILLER_99_224 ();
 b15zdnd11an1n64x5 FILLER_99_282 ();
 b15zdnd11an1n64x5 FILLER_99_346 ();
 b15zdnd11an1n64x5 FILLER_99_410 ();
 b15zdnd11an1n64x5 FILLER_99_474 ();
 b15zdnd11an1n64x5 FILLER_99_538 ();
 b15zdnd11an1n64x5 FILLER_99_602 ();
 b15zdnd11an1n64x5 FILLER_99_666 ();
 b15zdnd11an1n64x5 FILLER_99_730 ();
 b15zdnd11an1n64x5 FILLER_99_794 ();
 b15zdnd11an1n64x5 FILLER_99_867 ();
 b15zdnd11an1n64x5 FILLER_99_931 ();
 b15zdnd11an1n64x5 FILLER_99_995 ();
 b15zdnd11an1n64x5 FILLER_99_1059 ();
 b15zdnd11an1n64x5 FILLER_99_1123 ();
 b15zdnd11an1n64x5 FILLER_99_1187 ();
 b15zdnd11an1n64x5 FILLER_99_1251 ();
 b15zdnd11an1n64x5 FILLER_99_1315 ();
 b15zdnd11an1n64x5 FILLER_99_1379 ();
 b15zdnd11an1n32x5 FILLER_99_1443 ();
 b15zdnd11an1n08x5 FILLER_99_1475 ();
 b15zdnd00an1n02x5 FILLER_99_1483 ();
 b15zdnd00an1n01x5 FILLER_99_1485 ();
 b15zdnd00an1n02x5 FILLER_99_2257 ();
 b15zdnd11an1n08x5 FILLER_99_2271 ();
 b15zdnd11an1n04x5 FILLER_99_2279 ();
 b15zdnd00an1n01x5 FILLER_99_2283 ();
 b15zdnd11an1n64x5 FILLER_100_8 ();
 b15zdnd11an1n64x5 FILLER_100_72 ();
 b15zdnd11an1n64x5 FILLER_100_136 ();
 b15zdnd11an1n32x5 FILLER_100_200 ();
 b15zdnd11an1n08x5 FILLER_100_232 ();
 b15zdnd00an1n01x5 FILLER_100_240 ();
 b15zdnd11an1n64x5 FILLER_100_283 ();
 b15zdnd11an1n64x5 FILLER_100_347 ();
 b15zdnd11an1n08x5 FILLER_100_411 ();
 b15zdnd11an1n04x5 FILLER_100_419 ();
 b15zdnd00an1n02x5 FILLER_100_423 ();
 b15zdnd11an1n64x5 FILLER_100_431 ();
 b15zdnd11an1n64x5 FILLER_100_495 ();
 b15zdnd11an1n64x5 FILLER_100_559 ();
 b15zdnd11an1n64x5 FILLER_100_623 ();
 b15zdnd11an1n16x5 FILLER_100_687 ();
 b15zdnd11an1n08x5 FILLER_100_703 ();
 b15zdnd11an1n04x5 FILLER_100_711 ();
 b15zdnd00an1n02x5 FILLER_100_715 ();
 b15zdnd00an1n01x5 FILLER_100_717 ();
 b15zdnd11an1n64x5 FILLER_100_726 ();
 b15zdnd11an1n64x5 FILLER_100_790 ();
 b15zdnd11an1n64x5 FILLER_100_854 ();
 b15zdnd11an1n64x5 FILLER_100_918 ();
 b15zdnd11an1n64x5 FILLER_100_982 ();
 b15zdnd11an1n64x5 FILLER_100_1046 ();
 b15zdnd11an1n64x5 FILLER_100_1110 ();
 b15zdnd11an1n64x5 FILLER_100_1174 ();
 b15zdnd11an1n64x5 FILLER_100_1238 ();
 b15zdnd11an1n64x5 FILLER_100_1302 ();
 b15zdnd11an1n64x5 FILLER_100_1366 ();
 b15zdnd11an1n32x5 FILLER_100_1430 ();
 b15zdnd11an1n16x5 FILLER_100_1462 ();
 b15zdnd11an1n08x5 FILLER_100_2265 ();
 b15zdnd00an1n02x5 FILLER_100_2273 ();
 b15zdnd00an1n01x5 FILLER_100_2275 ();
 b15zdnd11an1n64x5 FILLER_101_0 ();
 b15zdnd11an1n64x5 FILLER_101_64 ();
 b15zdnd11an1n64x5 FILLER_101_128 ();
 b15zdnd11an1n32x5 FILLER_101_192 ();
 b15zdnd11an1n08x5 FILLER_101_224 ();
 b15zdnd11an1n04x5 FILLER_101_232 ();
 b15zdnd00an1n01x5 FILLER_101_236 ();
 b15zdnd11an1n64x5 FILLER_101_279 ();
 b15zdnd11an1n64x5 FILLER_101_343 ();
 b15zdnd11an1n64x5 FILLER_101_407 ();
 b15zdnd11an1n64x5 FILLER_101_471 ();
 b15zdnd11an1n64x5 FILLER_101_535 ();
 b15zdnd11an1n64x5 FILLER_101_599 ();
 b15zdnd11an1n64x5 FILLER_101_663 ();
 b15zdnd11an1n64x5 FILLER_101_727 ();
 b15zdnd11an1n64x5 FILLER_101_791 ();
 b15zdnd11an1n64x5 FILLER_101_855 ();
 b15zdnd11an1n64x5 FILLER_101_919 ();
 b15zdnd11an1n64x5 FILLER_101_983 ();
 b15zdnd11an1n64x5 FILLER_101_1047 ();
 b15zdnd11an1n64x5 FILLER_101_1111 ();
 b15zdnd11an1n64x5 FILLER_101_1175 ();
 b15zdnd11an1n64x5 FILLER_101_1239 ();
 b15zdnd11an1n08x5 FILLER_101_1303 ();
 b15zdnd11an1n64x5 FILLER_101_1353 ();
 b15zdnd11an1n64x5 FILLER_101_1417 ();
 b15zdnd11an1n04x5 FILLER_101_1481 ();
 b15zdnd00an1n01x5 FILLER_101_1485 ();
 b15zdnd00an1n02x5 FILLER_101_2257 ();
 b15zdnd11an1n16x5 FILLER_101_2262 ();
 b15zdnd11an1n04x5 FILLER_101_2278 ();
 b15zdnd00an1n02x5 FILLER_101_2282 ();
 b15zdnd11an1n64x5 FILLER_102_8 ();
 b15zdnd11an1n64x5 FILLER_102_72 ();
 b15zdnd11an1n64x5 FILLER_102_136 ();
 b15zdnd11an1n32x5 FILLER_102_200 ();
 b15zdnd11an1n08x5 FILLER_102_232 ();
 b15zdnd11an1n64x5 FILLER_102_282 ();
 b15zdnd11an1n64x5 FILLER_102_346 ();
 b15zdnd11an1n64x5 FILLER_102_410 ();
 b15zdnd11an1n64x5 FILLER_102_474 ();
 b15zdnd11an1n64x5 FILLER_102_538 ();
 b15zdnd11an1n16x5 FILLER_102_602 ();
 b15zdnd11an1n04x5 FILLER_102_618 ();
 b15zdnd00an1n02x5 FILLER_102_622 ();
 b15zdnd00an1n01x5 FILLER_102_624 ();
 b15zdnd11an1n64x5 FILLER_102_651 ();
 b15zdnd00an1n02x5 FILLER_102_715 ();
 b15zdnd00an1n01x5 FILLER_102_717 ();
 b15zdnd11an1n64x5 FILLER_102_726 ();
 b15zdnd11an1n64x5 FILLER_102_790 ();
 b15zdnd11an1n64x5 FILLER_102_854 ();
 b15zdnd11an1n64x5 FILLER_102_918 ();
 b15zdnd11an1n64x5 FILLER_102_982 ();
 b15zdnd11an1n64x5 FILLER_102_1046 ();
 b15zdnd11an1n64x5 FILLER_102_1110 ();
 b15zdnd11an1n64x5 FILLER_102_1174 ();
 b15zdnd11an1n64x5 FILLER_102_1238 ();
 b15zdnd11an1n16x5 FILLER_102_1302 ();
 b15zdnd00an1n01x5 FILLER_102_1318 ();
 b15zdnd11an1n64x5 FILLER_102_1361 ();
 b15zdnd11an1n32x5 FILLER_102_1425 ();
 b15zdnd11an1n16x5 FILLER_102_1457 ();
 b15zdnd11an1n04x5 FILLER_102_1473 ();
 b15zdnd00an1n01x5 FILLER_102_1477 ();
 b15zdnd00an1n02x5 FILLER_102_2265 ();
 b15zdnd00an1n01x5 FILLER_102_2267 ();
 b15zdnd11an1n04x5 FILLER_102_2271 ();
 b15zdnd00an1n01x5 FILLER_102_2275 ();
 b15zdnd11an1n64x5 FILLER_103_0 ();
 b15zdnd11an1n64x5 FILLER_103_64 ();
 b15zdnd11an1n64x5 FILLER_103_128 ();
 b15zdnd11an1n64x5 FILLER_103_192 ();
 b15zdnd11an1n64x5 FILLER_103_256 ();
 b15zdnd11an1n64x5 FILLER_103_320 ();
 b15zdnd11an1n64x5 FILLER_103_384 ();
 b15zdnd11an1n64x5 FILLER_103_448 ();
 b15zdnd11an1n64x5 FILLER_103_512 ();
 b15zdnd11an1n64x5 FILLER_103_576 ();
 b15zdnd11an1n64x5 FILLER_103_640 ();
 b15zdnd11an1n64x5 FILLER_103_704 ();
 b15zdnd11an1n64x5 FILLER_103_768 ();
 b15zdnd11an1n64x5 FILLER_103_832 ();
 b15zdnd11an1n64x5 FILLER_103_896 ();
 b15zdnd11an1n64x5 FILLER_103_960 ();
 b15zdnd11an1n64x5 FILLER_103_1024 ();
 b15zdnd11an1n64x5 FILLER_103_1088 ();
 b15zdnd11an1n64x5 FILLER_103_1152 ();
 b15zdnd11an1n64x5 FILLER_103_1216 ();
 b15zdnd11an1n64x5 FILLER_103_1280 ();
 b15zdnd11an1n64x5 FILLER_103_1344 ();
 b15zdnd11an1n64x5 FILLER_103_1408 ();
 b15zdnd11an1n08x5 FILLER_103_1472 ();
 b15zdnd00an1n01x5 FILLER_103_1480 ();
 b15zdnd00an1n02x5 FILLER_103_1484 ();
 b15zdnd00an1n02x5 FILLER_103_2257 ();
 b15zdnd11an1n16x5 FILLER_103_2262 ();
 b15zdnd11an1n04x5 FILLER_103_2278 ();
 b15zdnd00an1n02x5 FILLER_103_2282 ();
 b15zdnd11an1n64x5 FILLER_104_8 ();
 b15zdnd11an1n64x5 FILLER_104_72 ();
 b15zdnd11an1n64x5 FILLER_104_136 ();
 b15zdnd11an1n64x5 FILLER_104_200 ();
 b15zdnd11an1n64x5 FILLER_104_264 ();
 b15zdnd11an1n64x5 FILLER_104_328 ();
 b15zdnd11an1n32x5 FILLER_104_392 ();
 b15zdnd11an1n08x5 FILLER_104_424 ();
 b15zdnd11an1n64x5 FILLER_104_442 ();
 b15zdnd11an1n64x5 FILLER_104_506 ();
 b15zdnd11an1n64x5 FILLER_104_570 ();
 b15zdnd11an1n64x5 FILLER_104_634 ();
 b15zdnd11an1n16x5 FILLER_104_698 ();
 b15zdnd11an1n04x5 FILLER_104_714 ();
 b15zdnd11an1n64x5 FILLER_104_726 ();
 b15zdnd11an1n64x5 FILLER_104_790 ();
 b15zdnd11an1n64x5 FILLER_104_854 ();
 b15zdnd11an1n64x5 FILLER_104_918 ();
 b15zdnd11an1n64x5 FILLER_104_982 ();
 b15zdnd11an1n64x5 FILLER_104_1046 ();
 b15zdnd11an1n64x5 FILLER_104_1110 ();
 b15zdnd11an1n64x5 FILLER_104_1174 ();
 b15zdnd11an1n64x5 FILLER_104_1238 ();
 b15zdnd11an1n64x5 FILLER_104_1302 ();
 b15zdnd11an1n64x5 FILLER_104_1366 ();
 b15zdnd11an1n32x5 FILLER_104_1430 ();
 b15zdnd11an1n16x5 FILLER_104_1462 ();
 b15zdnd11an1n08x5 FILLER_104_2265 ();
 b15zdnd00an1n02x5 FILLER_104_2273 ();
 b15zdnd00an1n01x5 FILLER_104_2275 ();
 b15zdnd11an1n64x5 FILLER_105_0 ();
 b15zdnd11an1n64x5 FILLER_105_64 ();
 b15zdnd11an1n64x5 FILLER_105_128 ();
 b15zdnd11an1n64x5 FILLER_105_192 ();
 b15zdnd11an1n64x5 FILLER_105_256 ();
 b15zdnd11an1n64x5 FILLER_105_320 ();
 b15zdnd11an1n64x5 FILLER_105_384 ();
 b15zdnd11an1n64x5 FILLER_105_448 ();
 b15zdnd11an1n64x5 FILLER_105_512 ();
 b15zdnd11an1n64x5 FILLER_105_576 ();
 b15zdnd11an1n64x5 FILLER_105_640 ();
 b15zdnd11an1n64x5 FILLER_105_729 ();
 b15zdnd11an1n64x5 FILLER_105_793 ();
 b15zdnd11an1n64x5 FILLER_105_857 ();
 b15zdnd11an1n64x5 FILLER_105_921 ();
 b15zdnd11an1n64x5 FILLER_105_985 ();
 b15zdnd11an1n64x5 FILLER_105_1049 ();
 b15zdnd11an1n64x5 FILLER_105_1113 ();
 b15zdnd11an1n32x5 FILLER_105_1177 ();
 b15zdnd11an1n16x5 FILLER_105_1209 ();
 b15zdnd11an1n08x5 FILLER_105_1225 ();
 b15zdnd00an1n02x5 FILLER_105_1233 ();
 b15zdnd00an1n01x5 FILLER_105_1235 ();
 b15zdnd11an1n04x5 FILLER_105_1239 ();
 b15zdnd11an1n64x5 FILLER_105_1270 ();
 b15zdnd11an1n64x5 FILLER_105_1334 ();
 b15zdnd11an1n64x5 FILLER_105_1398 ();
 b15zdnd11an1n08x5 FILLER_105_1462 ();
 b15zdnd11an1n04x5 FILLER_105_1470 ();
 b15zdnd11an1n04x5 FILLER_105_1477 ();
 b15zdnd00an1n02x5 FILLER_105_1484 ();
 b15zdnd11an1n16x5 FILLER_105_2257 ();
 b15zdnd00an1n02x5 FILLER_105_2273 ();
 b15zdnd00an1n02x5 FILLER_105_2282 ();
 b15zdnd11an1n64x5 FILLER_106_8 ();
 b15zdnd11an1n64x5 FILLER_106_72 ();
 b15zdnd11an1n64x5 FILLER_106_136 ();
 b15zdnd11an1n64x5 FILLER_106_200 ();
 b15zdnd11an1n64x5 FILLER_106_264 ();
 b15zdnd11an1n64x5 FILLER_106_328 ();
 b15zdnd11an1n16x5 FILLER_106_392 ();
 b15zdnd11an1n16x5 FILLER_106_420 ();
 b15zdnd11an1n04x5 FILLER_106_436 ();
 b15zdnd00an1n01x5 FILLER_106_440 ();
 b15zdnd11an1n04x5 FILLER_106_451 ();
 b15zdnd11an1n64x5 FILLER_106_465 ();
 b15zdnd11an1n64x5 FILLER_106_529 ();
 b15zdnd11an1n64x5 FILLER_106_593 ();
 b15zdnd11an1n32x5 FILLER_106_657 ();
 b15zdnd11an1n08x5 FILLER_106_689 ();
 b15zdnd11an1n04x5 FILLER_106_697 ();
 b15zdnd11an1n04x5 FILLER_106_704 ();
 b15zdnd11an1n04x5 FILLER_106_711 ();
 b15zdnd00an1n02x5 FILLER_106_715 ();
 b15zdnd00an1n01x5 FILLER_106_717 ();
 b15zdnd11an1n64x5 FILLER_106_726 ();
 b15zdnd11an1n64x5 FILLER_106_790 ();
 b15zdnd11an1n64x5 FILLER_106_854 ();
 b15zdnd11an1n64x5 FILLER_106_918 ();
 b15zdnd11an1n64x5 FILLER_106_982 ();
 b15zdnd11an1n64x5 FILLER_106_1046 ();
 b15zdnd11an1n64x5 FILLER_106_1110 ();
 b15zdnd11an1n64x5 FILLER_106_1174 ();
 b15zdnd11an1n64x5 FILLER_106_1238 ();
 b15zdnd11an1n64x5 FILLER_106_1302 ();
 b15zdnd11an1n64x5 FILLER_106_1366 ();
 b15zdnd11an1n32x5 FILLER_106_1430 ();
 b15zdnd11an1n08x5 FILLER_106_1462 ();
 b15zdnd00an1n02x5 FILLER_106_1470 ();
 b15zdnd00an1n01x5 FILLER_106_1472 ();
 b15zdnd00an1n02x5 FILLER_106_1476 ();
 b15zdnd11an1n08x5 FILLER_106_2265 ();
 b15zdnd00an1n02x5 FILLER_106_2273 ();
 b15zdnd00an1n01x5 FILLER_106_2275 ();
 b15zdnd11an1n64x5 FILLER_107_0 ();
 b15zdnd11an1n64x5 FILLER_107_64 ();
 b15zdnd11an1n64x5 FILLER_107_128 ();
 b15zdnd11an1n64x5 FILLER_107_192 ();
 b15zdnd11an1n64x5 FILLER_107_256 ();
 b15zdnd11an1n64x5 FILLER_107_320 ();
 b15zdnd11an1n16x5 FILLER_107_384 ();
 b15zdnd11an1n08x5 FILLER_107_400 ();
 b15zdnd11an1n04x5 FILLER_107_408 ();
 b15zdnd11an1n16x5 FILLER_107_422 ();
 b15zdnd11an1n08x5 FILLER_107_438 ();
 b15zdnd11an1n64x5 FILLER_107_456 ();
 b15zdnd11an1n64x5 FILLER_107_520 ();
 b15zdnd11an1n64x5 FILLER_107_584 ();
 b15zdnd11an1n32x5 FILLER_107_648 ();
 b15zdnd11an1n16x5 FILLER_107_680 ();
 b15zdnd11an1n08x5 FILLER_107_696 ();
 b15zdnd11an1n04x5 FILLER_107_704 ();
 b15zdnd00an1n01x5 FILLER_107_708 ();
 b15zdnd11an1n08x5 FILLER_107_712 ();
 b15zdnd00an1n01x5 FILLER_107_720 ();
 b15zdnd11an1n08x5 FILLER_107_724 ();
 b15zdnd00an1n02x5 FILLER_107_732 ();
 b15zdnd11an1n64x5 FILLER_107_759 ();
 b15zdnd11an1n64x5 FILLER_107_823 ();
 b15zdnd11an1n64x5 FILLER_107_887 ();
 b15zdnd11an1n64x5 FILLER_107_951 ();
 b15zdnd11an1n64x5 FILLER_107_1015 ();
 b15zdnd11an1n64x5 FILLER_107_1079 ();
 b15zdnd11an1n64x5 FILLER_107_1143 ();
 b15zdnd11an1n64x5 FILLER_107_1207 ();
 b15zdnd11an1n64x5 FILLER_107_1271 ();
 b15zdnd11an1n64x5 FILLER_107_1335 ();
 b15zdnd11an1n64x5 FILLER_107_1399 ();
 b15zdnd11an1n16x5 FILLER_107_1463 ();
 b15zdnd11an1n04x5 FILLER_107_1479 ();
 b15zdnd00an1n02x5 FILLER_107_1483 ();
 b15zdnd00an1n01x5 FILLER_107_1485 ();
 b15zdnd11an1n16x5 FILLER_107_2257 ();
 b15zdnd00an1n01x5 FILLER_107_2273 ();
 b15zdnd00an1n02x5 FILLER_107_2282 ();
 b15zdnd11an1n64x5 FILLER_108_8 ();
 b15zdnd11an1n64x5 FILLER_108_72 ();
 b15zdnd11an1n64x5 FILLER_108_136 ();
 b15zdnd11an1n64x5 FILLER_108_200 ();
 b15zdnd11an1n64x5 FILLER_108_264 ();
 b15zdnd11an1n64x5 FILLER_108_328 ();
 b15zdnd11an1n08x5 FILLER_108_392 ();
 b15zdnd00an1n02x5 FILLER_108_400 ();
 b15zdnd11an1n04x5 FILLER_108_405 ();
 b15zdnd11an1n64x5 FILLER_108_418 ();
 b15zdnd11an1n64x5 FILLER_108_482 ();
 b15zdnd11an1n64x5 FILLER_108_546 ();
 b15zdnd11an1n64x5 FILLER_108_610 ();
 b15zdnd11an1n32x5 FILLER_108_674 ();
 b15zdnd11an1n08x5 FILLER_108_706 ();
 b15zdnd11an1n04x5 FILLER_108_714 ();
 b15zdnd11an1n64x5 FILLER_108_726 ();
 b15zdnd11an1n64x5 FILLER_108_790 ();
 b15zdnd11an1n64x5 FILLER_108_854 ();
 b15zdnd11an1n64x5 FILLER_108_918 ();
 b15zdnd11an1n64x5 FILLER_108_982 ();
 b15zdnd11an1n64x5 FILLER_108_1046 ();
 b15zdnd11an1n64x5 FILLER_108_1110 ();
 b15zdnd11an1n64x5 FILLER_108_1174 ();
 b15zdnd11an1n64x5 FILLER_108_1238 ();
 b15zdnd11an1n08x5 FILLER_108_1302 ();
 b15zdnd11an1n04x5 FILLER_108_1310 ();
 b15zdnd11an1n64x5 FILLER_108_1322 ();
 b15zdnd11an1n64x5 FILLER_108_1386 ();
 b15zdnd11an1n16x5 FILLER_108_1450 ();
 b15zdnd11an1n08x5 FILLER_108_1466 ();
 b15zdnd11an1n04x5 FILLER_108_1474 ();
 b15zdnd11an1n04x5 FILLER_108_2265 ();
 b15zdnd00an1n02x5 FILLER_108_2274 ();
 b15zdnd11an1n64x5 FILLER_109_0 ();
 b15zdnd11an1n64x5 FILLER_109_64 ();
 b15zdnd11an1n64x5 FILLER_109_128 ();
 b15zdnd11an1n64x5 FILLER_109_192 ();
 b15zdnd11an1n64x5 FILLER_109_256 ();
 b15zdnd11an1n64x5 FILLER_109_320 ();
 b15zdnd11an1n64x5 FILLER_109_384 ();
 b15zdnd11an1n64x5 FILLER_109_448 ();
 b15zdnd11an1n64x5 FILLER_109_512 ();
 b15zdnd11an1n64x5 FILLER_109_576 ();
 b15zdnd11an1n64x5 FILLER_109_640 ();
 b15zdnd11an1n64x5 FILLER_109_704 ();
 b15zdnd11an1n64x5 FILLER_109_768 ();
 b15zdnd11an1n64x5 FILLER_109_832 ();
 b15zdnd11an1n64x5 FILLER_109_896 ();
 b15zdnd11an1n64x5 FILLER_109_960 ();
 b15zdnd11an1n64x5 FILLER_109_1024 ();
 b15zdnd11an1n64x5 FILLER_109_1088 ();
 b15zdnd11an1n64x5 FILLER_109_1152 ();
 b15zdnd11an1n64x5 FILLER_109_1216 ();
 b15zdnd11an1n16x5 FILLER_109_1280 ();
 b15zdnd00an1n02x5 FILLER_109_1296 ();
 b15zdnd11an1n64x5 FILLER_109_1306 ();
 b15zdnd11an1n64x5 FILLER_109_1370 ();
 b15zdnd11an1n32x5 FILLER_109_1434 ();
 b15zdnd11an1n16x5 FILLER_109_1466 ();
 b15zdnd11an1n04x5 FILLER_109_1482 ();
 b15zdnd11an1n16x5 FILLER_109_2257 ();
 b15zdnd11an1n08x5 FILLER_109_2273 ();
 b15zdnd00an1n02x5 FILLER_109_2281 ();
 b15zdnd00an1n01x5 FILLER_109_2283 ();
 b15zdnd11an1n64x5 FILLER_110_8 ();
 b15zdnd11an1n64x5 FILLER_110_72 ();
 b15zdnd11an1n64x5 FILLER_110_136 ();
 b15zdnd11an1n64x5 FILLER_110_200 ();
 b15zdnd11an1n64x5 FILLER_110_264 ();
 b15zdnd11an1n64x5 FILLER_110_328 ();
 b15zdnd11an1n64x5 FILLER_110_392 ();
 b15zdnd11an1n64x5 FILLER_110_456 ();
 b15zdnd11an1n64x5 FILLER_110_520 ();
 b15zdnd11an1n64x5 FILLER_110_584 ();
 b15zdnd11an1n64x5 FILLER_110_648 ();
 b15zdnd11an1n04x5 FILLER_110_712 ();
 b15zdnd00an1n02x5 FILLER_110_716 ();
 b15zdnd11an1n64x5 FILLER_110_726 ();
 b15zdnd11an1n64x5 FILLER_110_790 ();
 b15zdnd11an1n64x5 FILLER_110_854 ();
 b15zdnd11an1n64x5 FILLER_110_918 ();
 b15zdnd11an1n64x5 FILLER_110_982 ();
 b15zdnd11an1n64x5 FILLER_110_1046 ();
 b15zdnd11an1n64x5 FILLER_110_1110 ();
 b15zdnd11an1n64x5 FILLER_110_1174 ();
 b15zdnd11an1n64x5 FILLER_110_1238 ();
 b15zdnd11an1n64x5 FILLER_110_1302 ();
 b15zdnd11an1n64x5 FILLER_110_1366 ();
 b15zdnd11an1n32x5 FILLER_110_1430 ();
 b15zdnd11an1n16x5 FILLER_110_1462 ();
 b15zdnd11an1n08x5 FILLER_110_2265 ();
 b15zdnd00an1n02x5 FILLER_110_2273 ();
 b15zdnd00an1n01x5 FILLER_110_2275 ();
 b15zdnd11an1n64x5 FILLER_111_0 ();
 b15zdnd11an1n64x5 FILLER_111_64 ();
 b15zdnd11an1n64x5 FILLER_111_128 ();
 b15zdnd11an1n64x5 FILLER_111_192 ();
 b15zdnd11an1n64x5 FILLER_111_256 ();
 b15zdnd11an1n64x5 FILLER_111_320 ();
 b15zdnd11an1n64x5 FILLER_111_384 ();
 b15zdnd11an1n64x5 FILLER_111_448 ();
 b15zdnd11an1n64x5 FILLER_111_512 ();
 b15zdnd11an1n64x5 FILLER_111_576 ();
 b15zdnd11an1n64x5 FILLER_111_640 ();
 b15zdnd11an1n64x5 FILLER_111_704 ();
 b15zdnd11an1n64x5 FILLER_111_768 ();
 b15zdnd11an1n64x5 FILLER_111_832 ();
 b15zdnd11an1n64x5 FILLER_111_896 ();
 b15zdnd11an1n64x5 FILLER_111_960 ();
 b15zdnd11an1n64x5 FILLER_111_1024 ();
 b15zdnd11an1n64x5 FILLER_111_1088 ();
 b15zdnd11an1n64x5 FILLER_111_1152 ();
 b15zdnd11an1n64x5 FILLER_111_1216 ();
 b15zdnd11an1n64x5 FILLER_111_1280 ();
 b15zdnd11an1n64x5 FILLER_111_1344 ();
 b15zdnd11an1n64x5 FILLER_111_1408 ();
 b15zdnd11an1n08x5 FILLER_111_1472 ();
 b15zdnd11an1n04x5 FILLER_111_1480 ();
 b15zdnd00an1n02x5 FILLER_111_1484 ();
 b15zdnd11an1n08x5 FILLER_111_2257 ();
 b15zdnd11an1n04x5 FILLER_111_2265 ();
 b15zdnd00an1n02x5 FILLER_111_2269 ();
 b15zdnd00an1n01x5 FILLER_111_2271 ();
 b15zdnd11an1n04x5 FILLER_111_2280 ();
 b15zdnd11an1n64x5 FILLER_112_8 ();
 b15zdnd11an1n64x5 FILLER_112_72 ();
 b15zdnd11an1n64x5 FILLER_112_136 ();
 b15zdnd11an1n64x5 FILLER_112_200 ();
 b15zdnd11an1n64x5 FILLER_112_264 ();
 b15zdnd11an1n64x5 FILLER_112_328 ();
 b15zdnd11an1n64x5 FILLER_112_392 ();
 b15zdnd11an1n64x5 FILLER_112_456 ();
 b15zdnd11an1n64x5 FILLER_112_520 ();
 b15zdnd11an1n64x5 FILLER_112_584 ();
 b15zdnd11an1n64x5 FILLER_112_648 ();
 b15zdnd11an1n04x5 FILLER_112_712 ();
 b15zdnd00an1n02x5 FILLER_112_716 ();
 b15zdnd11an1n64x5 FILLER_112_726 ();
 b15zdnd11an1n64x5 FILLER_112_790 ();
 b15zdnd11an1n64x5 FILLER_112_854 ();
 b15zdnd11an1n64x5 FILLER_112_918 ();
 b15zdnd11an1n64x5 FILLER_112_982 ();
 b15zdnd11an1n64x5 FILLER_112_1046 ();
 b15zdnd11an1n64x5 FILLER_112_1110 ();
 b15zdnd11an1n64x5 FILLER_112_1174 ();
 b15zdnd11an1n64x5 FILLER_112_1238 ();
 b15zdnd11an1n64x5 FILLER_112_1302 ();
 b15zdnd11an1n64x5 FILLER_112_1366 ();
 b15zdnd11an1n32x5 FILLER_112_1430 ();
 b15zdnd11an1n16x5 FILLER_112_1462 ();
 b15zdnd11an1n08x5 FILLER_112_2265 ();
 b15zdnd00an1n02x5 FILLER_112_2273 ();
 b15zdnd00an1n01x5 FILLER_112_2275 ();
 b15zdnd11an1n64x5 FILLER_113_0 ();
 b15zdnd11an1n64x5 FILLER_113_64 ();
 b15zdnd11an1n64x5 FILLER_113_128 ();
 b15zdnd11an1n64x5 FILLER_113_192 ();
 b15zdnd11an1n64x5 FILLER_113_256 ();
 b15zdnd11an1n64x5 FILLER_113_320 ();
 b15zdnd11an1n64x5 FILLER_113_384 ();
 b15zdnd11an1n64x5 FILLER_113_448 ();
 b15zdnd11an1n64x5 FILLER_113_512 ();
 b15zdnd11an1n64x5 FILLER_113_576 ();
 b15zdnd11an1n64x5 FILLER_113_640 ();
 b15zdnd11an1n64x5 FILLER_113_704 ();
 b15zdnd11an1n64x5 FILLER_113_768 ();
 b15zdnd11an1n64x5 FILLER_113_832 ();
 b15zdnd11an1n64x5 FILLER_113_896 ();
 b15zdnd11an1n64x5 FILLER_113_960 ();
 b15zdnd11an1n64x5 FILLER_113_1024 ();
 b15zdnd11an1n64x5 FILLER_113_1088 ();
 b15zdnd11an1n64x5 FILLER_113_1152 ();
 b15zdnd11an1n64x5 FILLER_113_1216 ();
 b15zdnd11an1n64x5 FILLER_113_1280 ();
 b15zdnd11an1n64x5 FILLER_113_1344 ();
 b15zdnd11an1n64x5 FILLER_113_1408 ();
 b15zdnd11an1n08x5 FILLER_113_1472 ();
 b15zdnd11an1n04x5 FILLER_113_1480 ();
 b15zdnd00an1n02x5 FILLER_113_1484 ();
 b15zdnd11an1n16x5 FILLER_113_2257 ();
 b15zdnd11an1n08x5 FILLER_113_2273 ();
 b15zdnd00an1n02x5 FILLER_113_2281 ();
 b15zdnd00an1n01x5 FILLER_113_2283 ();
 b15zdnd11an1n64x5 FILLER_114_8 ();
 b15zdnd11an1n64x5 FILLER_114_72 ();
 b15zdnd11an1n64x5 FILLER_114_136 ();
 b15zdnd11an1n64x5 FILLER_114_200 ();
 b15zdnd11an1n64x5 FILLER_114_264 ();
 b15zdnd11an1n64x5 FILLER_114_328 ();
 b15zdnd11an1n64x5 FILLER_114_392 ();
 b15zdnd11an1n64x5 FILLER_114_456 ();
 b15zdnd11an1n64x5 FILLER_114_520 ();
 b15zdnd11an1n64x5 FILLER_114_584 ();
 b15zdnd11an1n64x5 FILLER_114_648 ();
 b15zdnd11an1n04x5 FILLER_114_712 ();
 b15zdnd00an1n02x5 FILLER_114_716 ();
 b15zdnd11an1n64x5 FILLER_114_726 ();
 b15zdnd11an1n64x5 FILLER_114_790 ();
 b15zdnd11an1n64x5 FILLER_114_854 ();
 b15zdnd11an1n64x5 FILLER_114_918 ();
 b15zdnd11an1n64x5 FILLER_114_982 ();
 b15zdnd11an1n64x5 FILLER_114_1046 ();
 b15zdnd11an1n64x5 FILLER_114_1110 ();
 b15zdnd11an1n64x5 FILLER_114_1174 ();
 b15zdnd11an1n64x5 FILLER_114_1238 ();
 b15zdnd11an1n64x5 FILLER_114_1302 ();
 b15zdnd11an1n64x5 FILLER_114_1366 ();
 b15zdnd11an1n32x5 FILLER_114_1430 ();
 b15zdnd11an1n16x5 FILLER_114_1462 ();
 b15zdnd11an1n08x5 FILLER_114_2265 ();
 b15zdnd00an1n02x5 FILLER_114_2273 ();
 b15zdnd00an1n01x5 FILLER_114_2275 ();
 b15zdnd11an1n64x5 FILLER_115_0 ();
 b15zdnd11an1n64x5 FILLER_115_64 ();
 b15zdnd11an1n64x5 FILLER_115_128 ();
 b15zdnd11an1n64x5 FILLER_115_192 ();
 b15zdnd11an1n64x5 FILLER_115_256 ();
 b15zdnd11an1n64x5 FILLER_115_320 ();
 b15zdnd11an1n64x5 FILLER_115_384 ();
 b15zdnd11an1n64x5 FILLER_115_448 ();
 b15zdnd11an1n64x5 FILLER_115_512 ();
 b15zdnd11an1n64x5 FILLER_115_576 ();
 b15zdnd11an1n64x5 FILLER_115_640 ();
 b15zdnd11an1n64x5 FILLER_115_704 ();
 b15zdnd11an1n64x5 FILLER_115_768 ();
 b15zdnd11an1n64x5 FILLER_115_832 ();
 b15zdnd11an1n64x5 FILLER_115_896 ();
 b15zdnd11an1n64x5 FILLER_115_960 ();
 b15zdnd11an1n64x5 FILLER_115_1024 ();
 b15zdnd11an1n64x5 FILLER_115_1088 ();
 b15zdnd11an1n64x5 FILLER_115_1152 ();
 b15zdnd11an1n32x5 FILLER_115_1216 ();
 b15zdnd11an1n16x5 FILLER_115_1248 ();
 b15zdnd00an1n02x5 FILLER_115_1264 ();
 b15zdnd00an1n01x5 FILLER_115_1266 ();
 b15zdnd11an1n64x5 FILLER_115_1309 ();
 b15zdnd11an1n64x5 FILLER_115_1373 ();
 b15zdnd11an1n32x5 FILLER_115_1437 ();
 b15zdnd11an1n16x5 FILLER_115_1469 ();
 b15zdnd00an1n01x5 FILLER_115_1485 ();
 b15zdnd11an1n16x5 FILLER_115_2257 ();
 b15zdnd11an1n08x5 FILLER_115_2273 ();
 b15zdnd00an1n02x5 FILLER_115_2281 ();
 b15zdnd00an1n01x5 FILLER_115_2283 ();
 b15zdnd11an1n64x5 FILLER_116_8 ();
 b15zdnd11an1n64x5 FILLER_116_72 ();
 b15zdnd11an1n64x5 FILLER_116_136 ();
 b15zdnd11an1n64x5 FILLER_116_200 ();
 b15zdnd11an1n64x5 FILLER_116_264 ();
 b15zdnd11an1n64x5 FILLER_116_328 ();
 b15zdnd11an1n64x5 FILLER_116_392 ();
 b15zdnd11an1n64x5 FILLER_116_456 ();
 b15zdnd11an1n64x5 FILLER_116_520 ();
 b15zdnd11an1n64x5 FILLER_116_584 ();
 b15zdnd11an1n64x5 FILLER_116_648 ();
 b15zdnd11an1n04x5 FILLER_116_712 ();
 b15zdnd00an1n02x5 FILLER_116_716 ();
 b15zdnd11an1n64x5 FILLER_116_726 ();
 b15zdnd11an1n64x5 FILLER_116_790 ();
 b15zdnd11an1n64x5 FILLER_116_854 ();
 b15zdnd11an1n32x5 FILLER_116_918 ();
 b15zdnd00an1n02x5 FILLER_116_950 ();
 b15zdnd00an1n01x5 FILLER_116_952 ();
 b15zdnd11an1n64x5 FILLER_116_956 ();
 b15zdnd11an1n64x5 FILLER_116_1020 ();
 b15zdnd11an1n64x5 FILLER_116_1084 ();
 b15zdnd11an1n64x5 FILLER_116_1148 ();
 b15zdnd11an1n64x5 FILLER_116_1212 ();
 b15zdnd11an1n64x5 FILLER_116_1276 ();
 b15zdnd11an1n64x5 FILLER_116_1340 ();
 b15zdnd11an1n64x5 FILLER_116_1404 ();
 b15zdnd11an1n08x5 FILLER_116_1468 ();
 b15zdnd00an1n02x5 FILLER_116_1476 ();
 b15zdnd11an1n08x5 FILLER_116_2265 ();
 b15zdnd00an1n02x5 FILLER_116_2273 ();
 b15zdnd00an1n01x5 FILLER_116_2275 ();
 b15zdnd11an1n64x5 FILLER_117_0 ();
 b15zdnd11an1n64x5 FILLER_117_64 ();
 b15zdnd11an1n64x5 FILLER_117_128 ();
 b15zdnd11an1n64x5 FILLER_117_192 ();
 b15zdnd11an1n64x5 FILLER_117_256 ();
 b15zdnd11an1n64x5 FILLER_117_320 ();
 b15zdnd11an1n64x5 FILLER_117_384 ();
 b15zdnd11an1n64x5 FILLER_117_448 ();
 b15zdnd11an1n64x5 FILLER_117_512 ();
 b15zdnd11an1n64x5 FILLER_117_576 ();
 b15zdnd11an1n64x5 FILLER_117_640 ();
 b15zdnd00an1n02x5 FILLER_117_704 ();
 b15zdnd11an1n64x5 FILLER_117_748 ();
 b15zdnd11an1n64x5 FILLER_117_812 ();
 b15zdnd11an1n64x5 FILLER_117_876 ();
 b15zdnd11an1n08x5 FILLER_117_940 ();
 b15zdnd11an1n04x5 FILLER_117_948 ();
 b15zdnd11an1n16x5 FILLER_117_979 ();
 b15zdnd00an1n01x5 FILLER_117_995 ();
 b15zdnd11an1n04x5 FILLER_117_999 ();
 b15zdnd00an1n02x5 FILLER_117_1003 ();
 b15zdnd11an1n64x5 FILLER_117_1008 ();
 b15zdnd11an1n64x5 FILLER_117_1072 ();
 b15zdnd11an1n64x5 FILLER_117_1136 ();
 b15zdnd11an1n64x5 FILLER_117_1200 ();
 b15zdnd11an1n64x5 FILLER_117_1264 ();
 b15zdnd11an1n64x5 FILLER_117_1328 ();
 b15zdnd11an1n64x5 FILLER_117_1392 ();
 b15zdnd11an1n16x5 FILLER_117_1456 ();
 b15zdnd11an1n08x5 FILLER_117_1472 ();
 b15zdnd11an1n04x5 FILLER_117_1480 ();
 b15zdnd00an1n02x5 FILLER_117_1484 ();
 b15zdnd11an1n16x5 FILLER_117_2257 ();
 b15zdnd11an1n08x5 FILLER_117_2273 ();
 b15zdnd00an1n02x5 FILLER_117_2281 ();
 b15zdnd00an1n01x5 FILLER_117_2283 ();
 b15zdnd11an1n64x5 FILLER_118_8 ();
 b15zdnd11an1n64x5 FILLER_118_72 ();
 b15zdnd11an1n64x5 FILLER_118_136 ();
 b15zdnd11an1n64x5 FILLER_118_200 ();
 b15zdnd11an1n64x5 FILLER_118_264 ();
 b15zdnd11an1n64x5 FILLER_118_328 ();
 b15zdnd11an1n64x5 FILLER_118_392 ();
 b15zdnd11an1n64x5 FILLER_118_456 ();
 b15zdnd11an1n64x5 FILLER_118_520 ();
 b15zdnd11an1n64x5 FILLER_118_584 ();
 b15zdnd11an1n64x5 FILLER_118_648 ();
 b15zdnd11an1n04x5 FILLER_118_712 ();
 b15zdnd00an1n02x5 FILLER_118_716 ();
 b15zdnd11an1n64x5 FILLER_118_726 ();
 b15zdnd11an1n64x5 FILLER_118_790 ();
 b15zdnd11an1n64x5 FILLER_118_854 ();
 b15zdnd11an1n64x5 FILLER_118_918 ();
 b15zdnd11an1n08x5 FILLER_118_982 ();
 b15zdnd11an1n64x5 FILLER_118_1034 ();
 b15zdnd11an1n64x5 FILLER_118_1098 ();
 b15zdnd11an1n64x5 FILLER_118_1162 ();
 b15zdnd11an1n64x5 FILLER_118_1226 ();
 b15zdnd11an1n64x5 FILLER_118_1290 ();
 b15zdnd11an1n64x5 FILLER_118_1354 ();
 b15zdnd11an1n32x5 FILLER_118_1418 ();
 b15zdnd11an1n16x5 FILLER_118_1450 ();
 b15zdnd11an1n08x5 FILLER_118_1466 ();
 b15zdnd11an1n04x5 FILLER_118_1474 ();
 b15zdnd11an1n08x5 FILLER_118_2265 ();
 b15zdnd00an1n02x5 FILLER_118_2273 ();
 b15zdnd00an1n01x5 FILLER_118_2275 ();
 b15zdnd11an1n64x5 FILLER_119_0 ();
 b15zdnd11an1n64x5 FILLER_119_64 ();
 b15zdnd11an1n64x5 FILLER_119_128 ();
 b15zdnd11an1n64x5 FILLER_119_192 ();
 b15zdnd11an1n64x5 FILLER_119_256 ();
 b15zdnd11an1n64x5 FILLER_119_320 ();
 b15zdnd11an1n64x5 FILLER_119_384 ();
 b15zdnd11an1n64x5 FILLER_119_448 ();
 b15zdnd11an1n64x5 FILLER_119_512 ();
 b15zdnd11an1n64x5 FILLER_119_576 ();
 b15zdnd11an1n64x5 FILLER_119_640 ();
 b15zdnd11an1n04x5 FILLER_119_704 ();
 b15zdnd00an1n02x5 FILLER_119_708 ();
 b15zdnd00an1n01x5 FILLER_119_710 ();
 b15zdnd11an1n64x5 FILLER_119_753 ();
 b15zdnd11an1n64x5 FILLER_119_817 ();
 b15zdnd11an1n64x5 FILLER_119_881 ();
 b15zdnd11an1n32x5 FILLER_119_945 ();
 b15zdnd11an1n16x5 FILLER_119_977 ();
 b15zdnd11an1n08x5 FILLER_119_993 ();
 b15zdnd11an1n04x5 FILLER_119_1001 ();
 b15zdnd00an1n02x5 FILLER_119_1005 ();
 b15zdnd11an1n64x5 FILLER_119_1010 ();
 b15zdnd11an1n64x5 FILLER_119_1074 ();
 b15zdnd11an1n64x5 FILLER_119_1138 ();
 b15zdnd11an1n64x5 FILLER_119_1202 ();
 b15zdnd11an1n64x5 FILLER_119_1266 ();
 b15zdnd11an1n64x5 FILLER_119_1330 ();
 b15zdnd11an1n64x5 FILLER_119_1394 ();
 b15zdnd11an1n16x5 FILLER_119_1458 ();
 b15zdnd11an1n08x5 FILLER_119_1474 ();
 b15zdnd11an1n04x5 FILLER_119_1482 ();
 b15zdnd11an1n16x5 FILLER_119_2257 ();
 b15zdnd11an1n08x5 FILLER_119_2273 ();
 b15zdnd00an1n02x5 FILLER_119_2281 ();
 b15zdnd00an1n01x5 FILLER_119_2283 ();
 b15zdnd11an1n64x5 FILLER_120_8 ();
 b15zdnd11an1n64x5 FILLER_120_72 ();
 b15zdnd11an1n64x5 FILLER_120_136 ();
 b15zdnd11an1n64x5 FILLER_120_200 ();
 b15zdnd11an1n64x5 FILLER_120_264 ();
 b15zdnd11an1n64x5 FILLER_120_328 ();
 b15zdnd11an1n64x5 FILLER_120_392 ();
 b15zdnd11an1n64x5 FILLER_120_456 ();
 b15zdnd11an1n64x5 FILLER_120_520 ();
 b15zdnd11an1n64x5 FILLER_120_584 ();
 b15zdnd11an1n64x5 FILLER_120_648 ();
 b15zdnd11an1n04x5 FILLER_120_712 ();
 b15zdnd00an1n02x5 FILLER_120_716 ();
 b15zdnd11an1n64x5 FILLER_120_726 ();
 b15zdnd11an1n64x5 FILLER_120_790 ();
 b15zdnd11an1n64x5 FILLER_120_854 ();
 b15zdnd11an1n64x5 FILLER_120_918 ();
 b15zdnd11an1n16x5 FILLER_120_982 ();
 b15zdnd11an1n64x5 FILLER_120_1042 ();
 b15zdnd11an1n64x5 FILLER_120_1106 ();
 b15zdnd11an1n64x5 FILLER_120_1170 ();
 b15zdnd11an1n16x5 FILLER_120_1234 ();
 b15zdnd11an1n08x5 FILLER_120_1250 ();
 b15zdnd11an1n04x5 FILLER_120_1258 ();
 b15zdnd00an1n01x5 FILLER_120_1262 ();
 b15zdnd11an1n64x5 FILLER_120_1305 ();
 b15zdnd11an1n64x5 FILLER_120_1369 ();
 b15zdnd11an1n32x5 FILLER_120_1433 ();
 b15zdnd11an1n08x5 FILLER_120_1465 ();
 b15zdnd11an1n04x5 FILLER_120_1473 ();
 b15zdnd00an1n01x5 FILLER_120_1477 ();
 b15zdnd11an1n08x5 FILLER_120_2265 ();
 b15zdnd00an1n02x5 FILLER_120_2273 ();
 b15zdnd00an1n01x5 FILLER_120_2275 ();
 b15zdnd11an1n64x5 FILLER_121_0 ();
 b15zdnd11an1n64x5 FILLER_121_64 ();
 b15zdnd11an1n64x5 FILLER_121_128 ();
 b15zdnd11an1n64x5 FILLER_121_192 ();
 b15zdnd11an1n64x5 FILLER_121_256 ();
 b15zdnd11an1n64x5 FILLER_121_320 ();
 b15zdnd11an1n64x5 FILLER_121_384 ();
 b15zdnd11an1n64x5 FILLER_121_448 ();
 b15zdnd11an1n64x5 FILLER_121_512 ();
 b15zdnd11an1n64x5 FILLER_121_576 ();
 b15zdnd11an1n64x5 FILLER_121_640 ();
 b15zdnd11an1n64x5 FILLER_121_704 ();
 b15zdnd11an1n64x5 FILLER_121_768 ();
 b15zdnd11an1n64x5 FILLER_121_832 ();
 b15zdnd11an1n64x5 FILLER_121_896 ();
 b15zdnd11an1n08x5 FILLER_121_960 ();
 b15zdnd11an1n04x5 FILLER_121_968 ();
 b15zdnd11an1n04x5 FILLER_121_1016 ();
 b15zdnd11an1n04x5 FILLER_121_1023 ();
 b15zdnd00an1n01x5 FILLER_121_1027 ();
 b15zdnd11an1n64x5 FILLER_121_1031 ();
 b15zdnd11an1n64x5 FILLER_121_1095 ();
 b15zdnd11an1n64x5 FILLER_121_1159 ();
 b15zdnd11an1n16x5 FILLER_121_1223 ();
 b15zdnd11an1n04x5 FILLER_121_1239 ();
 b15zdnd00an1n02x5 FILLER_121_1243 ();
 b15zdnd00an1n01x5 FILLER_121_1245 ();
 b15zdnd11an1n64x5 FILLER_121_1288 ();
 b15zdnd11an1n64x5 FILLER_121_1352 ();
 b15zdnd11an1n64x5 FILLER_121_1416 ();
 b15zdnd11an1n04x5 FILLER_121_1480 ();
 b15zdnd00an1n02x5 FILLER_121_1484 ();
 b15zdnd11an1n16x5 FILLER_121_2257 ();
 b15zdnd11an1n08x5 FILLER_121_2273 ();
 b15zdnd00an1n02x5 FILLER_121_2281 ();
 b15zdnd00an1n01x5 FILLER_121_2283 ();
 b15zdnd11an1n64x5 FILLER_122_8 ();
 b15zdnd11an1n64x5 FILLER_122_72 ();
 b15zdnd11an1n64x5 FILLER_122_136 ();
 b15zdnd11an1n64x5 FILLER_122_200 ();
 b15zdnd11an1n64x5 FILLER_122_264 ();
 b15zdnd11an1n64x5 FILLER_122_328 ();
 b15zdnd11an1n64x5 FILLER_122_392 ();
 b15zdnd11an1n64x5 FILLER_122_456 ();
 b15zdnd11an1n64x5 FILLER_122_520 ();
 b15zdnd11an1n16x5 FILLER_122_584 ();
 b15zdnd00an1n02x5 FILLER_122_600 ();
 b15zdnd11an1n64x5 FILLER_122_644 ();
 b15zdnd11an1n08x5 FILLER_122_708 ();
 b15zdnd00an1n02x5 FILLER_122_716 ();
 b15zdnd11an1n64x5 FILLER_122_726 ();
 b15zdnd11an1n64x5 FILLER_122_790 ();
 b15zdnd11an1n64x5 FILLER_122_854 ();
 b15zdnd11an1n64x5 FILLER_122_918 ();
 b15zdnd11an1n04x5 FILLER_122_982 ();
 b15zdnd00an1n02x5 FILLER_122_986 ();
 b15zdnd00an1n01x5 FILLER_122_988 ();
 b15zdnd11an1n04x5 FILLER_122_992 ();
 b15zdnd00an1n02x5 FILLER_122_996 ();
 b15zdnd00an1n01x5 FILLER_122_998 ();
 b15zdnd11an1n16x5 FILLER_122_1002 ();
 b15zdnd11an1n64x5 FILLER_122_1021 ();
 b15zdnd11an1n64x5 FILLER_122_1085 ();
 b15zdnd11an1n64x5 FILLER_122_1149 ();
 b15zdnd11an1n64x5 FILLER_122_1213 ();
 b15zdnd11an1n64x5 FILLER_122_1277 ();
 b15zdnd11an1n64x5 FILLER_122_1341 ();
 b15zdnd11an1n64x5 FILLER_122_1405 ();
 b15zdnd11an1n08x5 FILLER_122_1469 ();
 b15zdnd00an1n01x5 FILLER_122_1477 ();
 b15zdnd11an1n08x5 FILLER_122_2265 ();
 b15zdnd00an1n02x5 FILLER_122_2273 ();
 b15zdnd00an1n01x5 FILLER_122_2275 ();
 b15zdnd11an1n64x5 FILLER_123_0 ();
 b15zdnd11an1n64x5 FILLER_123_64 ();
 b15zdnd11an1n04x5 FILLER_123_128 ();
 b15zdnd00an1n02x5 FILLER_123_132 ();
 b15zdnd11an1n64x5 FILLER_123_138 ();
 b15zdnd11an1n64x5 FILLER_123_202 ();
 b15zdnd11an1n64x5 FILLER_123_266 ();
 b15zdnd11an1n64x5 FILLER_123_330 ();
 b15zdnd11an1n64x5 FILLER_123_394 ();
 b15zdnd11an1n64x5 FILLER_123_458 ();
 b15zdnd11an1n64x5 FILLER_123_522 ();
 b15zdnd11an1n04x5 FILLER_123_586 ();
 b15zdnd00an1n02x5 FILLER_123_590 ();
 b15zdnd00an1n01x5 FILLER_123_592 ();
 b15zdnd11an1n64x5 FILLER_123_635 ();
 b15zdnd11an1n64x5 FILLER_123_699 ();
 b15zdnd11an1n64x5 FILLER_123_763 ();
 b15zdnd11an1n64x5 FILLER_123_827 ();
 b15zdnd11an1n64x5 FILLER_123_891 ();
 b15zdnd11an1n32x5 FILLER_123_955 ();
 b15zdnd00an1n02x5 FILLER_123_987 ();
 b15zdnd00an1n01x5 FILLER_123_989 ();
 b15zdnd11an1n64x5 FILLER_123_993 ();
 b15zdnd11an1n64x5 FILLER_123_1057 ();
 b15zdnd11an1n64x5 FILLER_123_1121 ();
 b15zdnd11an1n64x5 FILLER_123_1185 ();
 b15zdnd11an1n64x5 FILLER_123_1249 ();
 b15zdnd11an1n64x5 FILLER_123_1313 ();
 b15zdnd11an1n64x5 FILLER_123_1377 ();
 b15zdnd11an1n32x5 FILLER_123_1441 ();
 b15zdnd11an1n08x5 FILLER_123_1473 ();
 b15zdnd11an1n04x5 FILLER_123_1481 ();
 b15zdnd00an1n01x5 FILLER_123_1485 ();
 b15zdnd11an1n16x5 FILLER_123_2257 ();
 b15zdnd11an1n08x5 FILLER_123_2273 ();
 b15zdnd00an1n02x5 FILLER_123_2281 ();
 b15zdnd00an1n01x5 FILLER_123_2283 ();
 b15zdnd11an1n64x5 FILLER_124_8 ();
 b15zdnd11an1n32x5 FILLER_124_72 ();
 b15zdnd11an1n16x5 FILLER_124_104 ();
 b15zdnd11an1n04x5 FILLER_124_120 ();
 b15zdnd00an1n01x5 FILLER_124_124 ();
 b15zdnd11an1n08x5 FILLER_124_138 ();
 b15zdnd00an1n02x5 FILLER_124_146 ();
 b15zdnd00an1n01x5 FILLER_124_148 ();
 b15zdnd11an1n64x5 FILLER_124_153 ();
 b15zdnd11an1n64x5 FILLER_124_217 ();
 b15zdnd11an1n64x5 FILLER_124_281 ();
 b15zdnd11an1n64x5 FILLER_124_345 ();
 b15zdnd11an1n64x5 FILLER_124_409 ();
 b15zdnd11an1n64x5 FILLER_124_473 ();
 b15zdnd11an1n64x5 FILLER_124_537 ();
 b15zdnd11an1n64x5 FILLER_124_601 ();
 b15zdnd11an1n32x5 FILLER_124_665 ();
 b15zdnd11an1n16x5 FILLER_124_697 ();
 b15zdnd11an1n04x5 FILLER_124_713 ();
 b15zdnd00an1n01x5 FILLER_124_717 ();
 b15zdnd11an1n64x5 FILLER_124_726 ();
 b15zdnd11an1n64x5 FILLER_124_790 ();
 b15zdnd11an1n64x5 FILLER_124_854 ();
 b15zdnd11an1n64x5 FILLER_124_918 ();
 b15zdnd11an1n64x5 FILLER_124_982 ();
 b15zdnd11an1n64x5 FILLER_124_1046 ();
 b15zdnd11an1n64x5 FILLER_124_1110 ();
 b15zdnd11an1n64x5 FILLER_124_1174 ();
 b15zdnd11an1n64x5 FILLER_124_1238 ();
 b15zdnd11an1n64x5 FILLER_124_1302 ();
 b15zdnd11an1n64x5 FILLER_124_1366 ();
 b15zdnd11an1n32x5 FILLER_124_1430 ();
 b15zdnd11an1n16x5 FILLER_124_1462 ();
 b15zdnd11an1n08x5 FILLER_124_2265 ();
 b15zdnd00an1n02x5 FILLER_124_2273 ();
 b15zdnd00an1n01x5 FILLER_124_2275 ();
 b15zdnd11an1n64x5 FILLER_125_0 ();
 b15zdnd11an1n64x5 FILLER_125_64 ();
 b15zdnd11an1n64x5 FILLER_125_128 ();
 b15zdnd11an1n64x5 FILLER_125_192 ();
 b15zdnd11an1n64x5 FILLER_125_256 ();
 b15zdnd11an1n64x5 FILLER_125_320 ();
 b15zdnd11an1n32x5 FILLER_125_384 ();
 b15zdnd11an1n08x5 FILLER_125_416 ();
 b15zdnd11an1n04x5 FILLER_125_424 ();
 b15zdnd00an1n01x5 FILLER_125_428 ();
 b15zdnd11an1n64x5 FILLER_125_439 ();
 b15zdnd11an1n64x5 FILLER_125_503 ();
 b15zdnd11an1n32x5 FILLER_125_567 ();
 b15zdnd11an1n04x5 FILLER_125_599 ();
 b15zdnd00an1n01x5 FILLER_125_603 ();
 b15zdnd11an1n64x5 FILLER_125_646 ();
 b15zdnd11an1n64x5 FILLER_125_710 ();
 b15zdnd11an1n64x5 FILLER_125_774 ();
 b15zdnd11an1n64x5 FILLER_125_838 ();
 b15zdnd11an1n64x5 FILLER_125_902 ();
 b15zdnd11an1n64x5 FILLER_125_966 ();
 b15zdnd11an1n64x5 FILLER_125_1030 ();
 b15zdnd11an1n64x5 FILLER_125_1094 ();
 b15zdnd11an1n64x5 FILLER_125_1158 ();
 b15zdnd11an1n64x5 FILLER_125_1222 ();
 b15zdnd11an1n64x5 FILLER_125_1286 ();
 b15zdnd11an1n64x5 FILLER_125_1350 ();
 b15zdnd11an1n64x5 FILLER_125_1414 ();
 b15zdnd11an1n08x5 FILLER_125_1478 ();
 b15zdnd11an1n16x5 FILLER_125_2257 ();
 b15zdnd11an1n08x5 FILLER_125_2273 ();
 b15zdnd00an1n02x5 FILLER_125_2281 ();
 b15zdnd00an1n01x5 FILLER_125_2283 ();
 b15zdnd11an1n64x5 FILLER_126_8 ();
 b15zdnd11an1n64x5 FILLER_126_72 ();
 b15zdnd11an1n32x5 FILLER_126_136 ();
 b15zdnd11an1n08x5 FILLER_126_168 ();
 b15zdnd11an1n04x5 FILLER_126_176 ();
 b15zdnd00an1n02x5 FILLER_126_180 ();
 b15zdnd11an1n64x5 FILLER_126_205 ();
 b15zdnd11an1n64x5 FILLER_126_269 ();
 b15zdnd11an1n64x5 FILLER_126_333 ();
 b15zdnd11an1n08x5 FILLER_126_397 ();
 b15zdnd00an1n02x5 FILLER_126_405 ();
 b15zdnd11an1n64x5 FILLER_126_414 ();
 b15zdnd11an1n64x5 FILLER_126_478 ();
 b15zdnd11an1n32x5 FILLER_126_542 ();
 b15zdnd11an1n08x5 FILLER_126_574 ();
 b15zdnd00an1n02x5 FILLER_126_582 ();
 b15zdnd00an1n01x5 FILLER_126_584 ();
 b15zdnd11an1n64x5 FILLER_126_627 ();
 b15zdnd11an1n16x5 FILLER_126_691 ();
 b15zdnd11an1n08x5 FILLER_126_707 ();
 b15zdnd00an1n02x5 FILLER_126_715 ();
 b15zdnd00an1n01x5 FILLER_126_717 ();
 b15zdnd11an1n64x5 FILLER_126_726 ();
 b15zdnd11an1n64x5 FILLER_126_790 ();
 b15zdnd11an1n64x5 FILLER_126_854 ();
 b15zdnd11an1n64x5 FILLER_126_918 ();
 b15zdnd11an1n64x5 FILLER_126_982 ();
 b15zdnd11an1n64x5 FILLER_126_1046 ();
 b15zdnd11an1n64x5 FILLER_126_1110 ();
 b15zdnd11an1n64x5 FILLER_126_1174 ();
 b15zdnd11an1n64x5 FILLER_126_1238 ();
 b15zdnd11an1n64x5 FILLER_126_1302 ();
 b15zdnd11an1n64x5 FILLER_126_1366 ();
 b15zdnd11an1n32x5 FILLER_126_1430 ();
 b15zdnd11an1n16x5 FILLER_126_1462 ();
 b15zdnd00an1n02x5 FILLER_126_2265 ();
 b15zdnd00an1n02x5 FILLER_126_2274 ();
 b15zdnd11an1n64x5 FILLER_127_0 ();
 b15zdnd11an1n32x5 FILLER_127_64 ();
 b15zdnd11an1n16x5 FILLER_127_96 ();
 b15zdnd11an1n08x5 FILLER_127_112 ();
 b15zdnd00an1n02x5 FILLER_127_120 ();
 b15zdnd11an1n64x5 FILLER_127_137 ();
 b15zdnd11an1n64x5 FILLER_127_201 ();
 b15zdnd11an1n64x5 FILLER_127_265 ();
 b15zdnd11an1n64x5 FILLER_127_329 ();
 b15zdnd11an1n64x5 FILLER_127_393 ();
 b15zdnd11an1n64x5 FILLER_127_457 ();
 b15zdnd11an1n64x5 FILLER_127_521 ();
 b15zdnd11an1n64x5 FILLER_127_585 ();
 b15zdnd11an1n64x5 FILLER_127_649 ();
 b15zdnd11an1n64x5 FILLER_127_713 ();
 b15zdnd11an1n64x5 FILLER_127_777 ();
 b15zdnd11an1n64x5 FILLER_127_841 ();
 b15zdnd11an1n64x5 FILLER_127_905 ();
 b15zdnd11an1n64x5 FILLER_127_969 ();
 b15zdnd11an1n64x5 FILLER_127_1033 ();
 b15zdnd11an1n64x5 FILLER_127_1097 ();
 b15zdnd11an1n64x5 FILLER_127_1161 ();
 b15zdnd11an1n64x5 FILLER_127_1225 ();
 b15zdnd11an1n64x5 FILLER_127_1289 ();
 b15zdnd11an1n64x5 FILLER_127_1353 ();
 b15zdnd11an1n64x5 FILLER_127_1417 ();
 b15zdnd11an1n04x5 FILLER_127_1481 ();
 b15zdnd00an1n01x5 FILLER_127_1485 ();
 b15zdnd11an1n16x5 FILLER_127_2257 ();
 b15zdnd00an1n02x5 FILLER_127_2273 ();
 b15zdnd00an1n01x5 FILLER_127_2275 ();
 b15zdnd00an1n02x5 FILLER_127_2282 ();
 b15zdnd11an1n64x5 FILLER_128_8 ();
 b15zdnd11an1n64x5 FILLER_128_72 ();
 b15zdnd11an1n64x5 FILLER_128_136 ();
 b15zdnd11an1n32x5 FILLER_128_200 ();
 b15zdnd00an1n02x5 FILLER_128_232 ();
 b15zdnd11an1n64x5 FILLER_128_276 ();
 b15zdnd11an1n64x5 FILLER_128_340 ();
 b15zdnd11an1n64x5 FILLER_128_404 ();
 b15zdnd11an1n64x5 FILLER_128_468 ();
 b15zdnd11an1n64x5 FILLER_128_532 ();
 b15zdnd11an1n64x5 FILLER_128_596 ();
 b15zdnd11an1n32x5 FILLER_128_660 ();
 b15zdnd11an1n16x5 FILLER_128_692 ();
 b15zdnd11an1n08x5 FILLER_128_708 ();
 b15zdnd00an1n02x5 FILLER_128_716 ();
 b15zdnd11an1n16x5 FILLER_128_726 ();
 b15zdnd11an1n08x5 FILLER_128_742 ();
 b15zdnd11an1n64x5 FILLER_128_761 ();
 b15zdnd11an1n64x5 FILLER_128_825 ();
 b15zdnd11an1n64x5 FILLER_128_889 ();
 b15zdnd11an1n64x5 FILLER_128_953 ();
 b15zdnd11an1n64x5 FILLER_128_1017 ();
 b15zdnd11an1n64x5 FILLER_128_1081 ();
 b15zdnd11an1n64x5 FILLER_128_1145 ();
 b15zdnd11an1n64x5 FILLER_128_1209 ();
 b15zdnd11an1n64x5 FILLER_128_1273 ();
 b15zdnd11an1n64x5 FILLER_128_1337 ();
 b15zdnd11an1n64x5 FILLER_128_1401 ();
 b15zdnd11an1n08x5 FILLER_128_1465 ();
 b15zdnd11an1n04x5 FILLER_128_1473 ();
 b15zdnd00an1n01x5 FILLER_128_1477 ();
 b15zdnd11an1n08x5 FILLER_128_2265 ();
 b15zdnd00an1n02x5 FILLER_128_2273 ();
 b15zdnd00an1n01x5 FILLER_128_2275 ();
 b15zdnd11an1n64x5 FILLER_129_0 ();
 b15zdnd11an1n64x5 FILLER_129_64 ();
 b15zdnd11an1n64x5 FILLER_129_128 ();
 b15zdnd11an1n64x5 FILLER_129_192 ();
 b15zdnd11an1n64x5 FILLER_129_256 ();
 b15zdnd11an1n64x5 FILLER_129_320 ();
 b15zdnd11an1n64x5 FILLER_129_384 ();
 b15zdnd11an1n64x5 FILLER_129_448 ();
 b15zdnd11an1n64x5 FILLER_129_512 ();
 b15zdnd11an1n64x5 FILLER_129_576 ();
 b15zdnd11an1n64x5 FILLER_129_640 ();
 b15zdnd11an1n64x5 FILLER_129_704 ();
 b15zdnd11an1n64x5 FILLER_129_768 ();
 b15zdnd11an1n64x5 FILLER_129_832 ();
 b15zdnd11an1n64x5 FILLER_129_896 ();
 b15zdnd11an1n64x5 FILLER_129_960 ();
 b15zdnd11an1n64x5 FILLER_129_1024 ();
 b15zdnd11an1n64x5 FILLER_129_1088 ();
 b15zdnd11an1n64x5 FILLER_129_1152 ();
 b15zdnd11an1n64x5 FILLER_129_1216 ();
 b15zdnd11an1n64x5 FILLER_129_1280 ();
 b15zdnd11an1n64x5 FILLER_129_1344 ();
 b15zdnd11an1n64x5 FILLER_129_1408 ();
 b15zdnd11an1n08x5 FILLER_129_1472 ();
 b15zdnd11an1n04x5 FILLER_129_1480 ();
 b15zdnd00an1n02x5 FILLER_129_1484 ();
 b15zdnd11an1n16x5 FILLER_129_2257 ();
 b15zdnd00an1n02x5 FILLER_129_2273 ();
 b15zdnd00an1n01x5 FILLER_129_2275 ();
 b15zdnd00an1n02x5 FILLER_129_2282 ();
 b15zdnd11an1n08x5 FILLER_130_8 ();
 b15zdnd11an1n04x5 FILLER_130_16 ();
 b15zdnd11an1n04x5 FILLER_130_25 ();
 b15zdnd11an1n04x5 FILLER_130_34 ();
 b15zdnd11an1n64x5 FILLER_130_42 ();
 b15zdnd11an1n32x5 FILLER_130_106 ();
 b15zdnd11an1n08x5 FILLER_130_138 ();
 b15zdnd11an1n64x5 FILLER_130_168 ();
 b15zdnd11an1n64x5 FILLER_130_232 ();
 b15zdnd11an1n64x5 FILLER_130_296 ();
 b15zdnd11an1n64x5 FILLER_130_360 ();
 b15zdnd11an1n64x5 FILLER_130_424 ();
 b15zdnd11an1n64x5 FILLER_130_488 ();
 b15zdnd11an1n64x5 FILLER_130_552 ();
 b15zdnd11an1n64x5 FILLER_130_616 ();
 b15zdnd11an1n32x5 FILLER_130_680 ();
 b15zdnd11an1n04x5 FILLER_130_712 ();
 b15zdnd00an1n02x5 FILLER_130_716 ();
 b15zdnd11an1n64x5 FILLER_130_726 ();
 b15zdnd11an1n64x5 FILLER_130_790 ();
 b15zdnd11an1n64x5 FILLER_130_854 ();
 b15zdnd11an1n64x5 FILLER_130_918 ();
 b15zdnd11an1n64x5 FILLER_130_982 ();
 b15zdnd11an1n64x5 FILLER_130_1046 ();
 b15zdnd11an1n64x5 FILLER_130_1110 ();
 b15zdnd11an1n64x5 FILLER_130_1174 ();
 b15zdnd11an1n64x5 FILLER_130_1238 ();
 b15zdnd11an1n64x5 FILLER_130_1302 ();
 b15zdnd11an1n64x5 FILLER_130_1366 ();
 b15zdnd11an1n32x5 FILLER_130_1430 ();
 b15zdnd11an1n16x5 FILLER_130_1462 ();
 b15zdnd11an1n08x5 FILLER_130_2265 ();
 b15zdnd00an1n02x5 FILLER_130_2273 ();
 b15zdnd00an1n01x5 FILLER_130_2275 ();
 b15zdnd11an1n08x5 FILLER_131_0 ();
 b15zdnd00an1n02x5 FILLER_131_8 ();
 b15zdnd00an1n01x5 FILLER_131_10 ();
 b15zdnd11an1n64x5 FILLER_131_53 ();
 b15zdnd11an1n64x5 FILLER_131_117 ();
 b15zdnd11an1n64x5 FILLER_131_181 ();
 b15zdnd11an1n64x5 FILLER_131_245 ();
 b15zdnd11an1n64x5 FILLER_131_309 ();
 b15zdnd11an1n32x5 FILLER_131_373 ();
 b15zdnd11an1n04x5 FILLER_131_405 ();
 b15zdnd00an1n02x5 FILLER_131_409 ();
 b15zdnd11an1n64x5 FILLER_131_419 ();
 b15zdnd11an1n64x5 FILLER_131_483 ();
 b15zdnd11an1n64x5 FILLER_131_547 ();
 b15zdnd11an1n64x5 FILLER_131_611 ();
 b15zdnd11an1n08x5 FILLER_131_675 ();
 b15zdnd11an1n04x5 FILLER_131_683 ();
 b15zdnd00an1n01x5 FILLER_131_687 ();
 b15zdnd11an1n64x5 FILLER_131_730 ();
 b15zdnd11an1n64x5 FILLER_131_794 ();
 b15zdnd11an1n64x5 FILLER_131_858 ();
 b15zdnd11an1n64x5 FILLER_131_922 ();
 b15zdnd11an1n64x5 FILLER_131_986 ();
 b15zdnd11an1n64x5 FILLER_131_1050 ();
 b15zdnd11an1n64x5 FILLER_131_1114 ();
 b15zdnd11an1n64x5 FILLER_131_1178 ();
 b15zdnd11an1n64x5 FILLER_131_1242 ();
 b15zdnd11an1n64x5 FILLER_131_1306 ();
 b15zdnd11an1n64x5 FILLER_131_1370 ();
 b15zdnd11an1n32x5 FILLER_131_1434 ();
 b15zdnd11an1n16x5 FILLER_131_1466 ();
 b15zdnd11an1n04x5 FILLER_131_1482 ();
 b15zdnd11an1n16x5 FILLER_131_2257 ();
 b15zdnd11an1n08x5 FILLER_131_2273 ();
 b15zdnd00an1n02x5 FILLER_131_2281 ();
 b15zdnd00an1n01x5 FILLER_131_2283 ();
 b15zdnd11an1n08x5 FILLER_132_8 ();
 b15zdnd11an1n04x5 FILLER_132_16 ();
 b15zdnd00an1n01x5 FILLER_132_20 ();
 b15zdnd11an1n64x5 FILLER_132_26 ();
 b15zdnd11an1n64x5 FILLER_132_90 ();
 b15zdnd11an1n64x5 FILLER_132_154 ();
 b15zdnd11an1n64x5 FILLER_132_218 ();
 b15zdnd11an1n64x5 FILLER_132_282 ();
 b15zdnd11an1n64x5 FILLER_132_346 ();
 b15zdnd11an1n64x5 FILLER_132_410 ();
 b15zdnd11an1n64x5 FILLER_132_474 ();
 b15zdnd11an1n64x5 FILLER_132_538 ();
 b15zdnd11an1n32x5 FILLER_132_602 ();
 b15zdnd11an1n16x5 FILLER_132_634 ();
 b15zdnd11an1n08x5 FILLER_132_650 ();
 b15zdnd11an1n04x5 FILLER_132_658 ();
 b15zdnd11an1n08x5 FILLER_132_704 ();
 b15zdnd11an1n04x5 FILLER_132_712 ();
 b15zdnd00an1n02x5 FILLER_132_716 ();
 b15zdnd11an1n64x5 FILLER_132_726 ();
 b15zdnd11an1n64x5 FILLER_132_790 ();
 b15zdnd11an1n64x5 FILLER_132_854 ();
 b15zdnd11an1n64x5 FILLER_132_918 ();
 b15zdnd11an1n64x5 FILLER_132_982 ();
 b15zdnd11an1n64x5 FILLER_132_1046 ();
 b15zdnd11an1n64x5 FILLER_132_1110 ();
 b15zdnd11an1n64x5 FILLER_132_1174 ();
 b15zdnd11an1n64x5 FILLER_132_1238 ();
 b15zdnd11an1n64x5 FILLER_132_1302 ();
 b15zdnd11an1n64x5 FILLER_132_1366 ();
 b15zdnd11an1n32x5 FILLER_132_1430 ();
 b15zdnd11an1n16x5 FILLER_132_1462 ();
 b15zdnd11an1n08x5 FILLER_132_2265 ();
 b15zdnd00an1n02x5 FILLER_132_2273 ();
 b15zdnd00an1n01x5 FILLER_132_2275 ();
 b15zdnd11an1n16x5 FILLER_133_0 ();
 b15zdnd00an1n02x5 FILLER_133_16 ();
 b15zdnd11an1n64x5 FILLER_133_23 ();
 b15zdnd11an1n64x5 FILLER_133_87 ();
 b15zdnd11an1n64x5 FILLER_133_151 ();
 b15zdnd11an1n64x5 FILLER_133_215 ();
 b15zdnd11an1n64x5 FILLER_133_279 ();
 b15zdnd11an1n64x5 FILLER_133_343 ();
 b15zdnd11an1n64x5 FILLER_133_407 ();
 b15zdnd11an1n64x5 FILLER_133_471 ();
 b15zdnd11an1n64x5 FILLER_133_535 ();
 b15zdnd11an1n64x5 FILLER_133_599 ();
 b15zdnd11an1n16x5 FILLER_133_663 ();
 b15zdnd11an1n04x5 FILLER_133_679 ();
 b15zdnd00an1n02x5 FILLER_133_683 ();
 b15zdnd11an1n64x5 FILLER_133_727 ();
 b15zdnd11an1n64x5 FILLER_133_791 ();
 b15zdnd11an1n64x5 FILLER_133_855 ();
 b15zdnd11an1n64x5 FILLER_133_919 ();
 b15zdnd11an1n64x5 FILLER_133_983 ();
 b15zdnd11an1n64x5 FILLER_133_1047 ();
 b15zdnd11an1n64x5 FILLER_133_1111 ();
 b15zdnd11an1n64x5 FILLER_133_1175 ();
 b15zdnd11an1n64x5 FILLER_133_1239 ();
 b15zdnd11an1n64x5 FILLER_133_1303 ();
 b15zdnd11an1n64x5 FILLER_133_1367 ();
 b15zdnd11an1n32x5 FILLER_133_1431 ();
 b15zdnd11an1n16x5 FILLER_133_1463 ();
 b15zdnd11an1n04x5 FILLER_133_1479 ();
 b15zdnd00an1n02x5 FILLER_133_1483 ();
 b15zdnd00an1n01x5 FILLER_133_1485 ();
 b15zdnd11an1n16x5 FILLER_133_2257 ();
 b15zdnd11an1n08x5 FILLER_133_2273 ();
 b15zdnd00an1n02x5 FILLER_133_2281 ();
 b15zdnd00an1n01x5 FILLER_133_2283 ();
 b15zdnd00an1n02x5 FILLER_134_8 ();
 b15zdnd11an1n64x5 FILLER_134_18 ();
 b15zdnd11an1n64x5 FILLER_134_82 ();
 b15zdnd11an1n64x5 FILLER_134_146 ();
 b15zdnd11an1n64x5 FILLER_134_210 ();
 b15zdnd11an1n64x5 FILLER_134_274 ();
 b15zdnd11an1n64x5 FILLER_134_338 ();
 b15zdnd11an1n64x5 FILLER_134_402 ();
 b15zdnd11an1n64x5 FILLER_134_466 ();
 b15zdnd11an1n64x5 FILLER_134_530 ();
 b15zdnd11an1n64x5 FILLER_134_594 ();
 b15zdnd11an1n32x5 FILLER_134_658 ();
 b15zdnd11an1n16x5 FILLER_134_690 ();
 b15zdnd11an1n08x5 FILLER_134_706 ();
 b15zdnd11an1n04x5 FILLER_134_714 ();
 b15zdnd11an1n64x5 FILLER_134_726 ();
 b15zdnd11an1n64x5 FILLER_134_790 ();
 b15zdnd11an1n64x5 FILLER_134_854 ();
 b15zdnd11an1n64x5 FILLER_134_918 ();
 b15zdnd11an1n64x5 FILLER_134_982 ();
 b15zdnd11an1n64x5 FILLER_134_1046 ();
 b15zdnd11an1n64x5 FILLER_134_1110 ();
 b15zdnd11an1n64x5 FILLER_134_1174 ();
 b15zdnd11an1n64x5 FILLER_134_1238 ();
 b15zdnd11an1n64x5 FILLER_134_1302 ();
 b15zdnd11an1n64x5 FILLER_134_1366 ();
 b15zdnd11an1n16x5 FILLER_134_1430 ();
 b15zdnd11an1n08x5 FILLER_134_1446 ();
 b15zdnd11an1n04x5 FILLER_134_1454 ();
 b15zdnd00an1n02x5 FILLER_134_1458 ();
 b15zdnd11an1n04x5 FILLER_134_1471 ();
 b15zdnd00an1n02x5 FILLER_134_1475 ();
 b15zdnd00an1n01x5 FILLER_134_1477 ();
 b15zdnd11an1n08x5 FILLER_134_2265 ();
 b15zdnd00an1n02x5 FILLER_134_2273 ();
 b15zdnd00an1n01x5 FILLER_134_2275 ();
 b15zdnd00an1n02x5 FILLER_135_0 ();
 b15zdnd11an1n04x5 FILLER_135_13 ();
 b15zdnd11an1n64x5 FILLER_135_28 ();
 b15zdnd11an1n64x5 FILLER_135_92 ();
 b15zdnd11an1n64x5 FILLER_135_156 ();
 b15zdnd11an1n64x5 FILLER_135_220 ();
 b15zdnd11an1n64x5 FILLER_135_284 ();
 b15zdnd11an1n64x5 FILLER_135_348 ();
 b15zdnd11an1n08x5 FILLER_135_412 ();
 b15zdnd11an1n04x5 FILLER_135_420 ();
 b15zdnd11an1n08x5 FILLER_135_438 ();
 b15zdnd11an1n04x5 FILLER_135_446 ();
 b15zdnd00an1n02x5 FILLER_135_450 ();
 b15zdnd00an1n01x5 FILLER_135_452 ();
 b15zdnd11an1n64x5 FILLER_135_471 ();
 b15zdnd11an1n64x5 FILLER_135_535 ();
 b15zdnd11an1n32x5 FILLER_135_599 ();
 b15zdnd11an1n16x5 FILLER_135_631 ();
 b15zdnd11an1n08x5 FILLER_135_647 ();
 b15zdnd11an1n08x5 FILLER_135_697 ();
 b15zdnd11an1n04x5 FILLER_135_705 ();
 b15zdnd00an1n01x5 FILLER_135_709 ();
 b15zdnd11an1n64x5 FILLER_135_719 ();
 b15zdnd11an1n64x5 FILLER_135_783 ();
 b15zdnd11an1n64x5 FILLER_135_847 ();
 b15zdnd11an1n64x5 FILLER_135_911 ();
 b15zdnd11an1n64x5 FILLER_135_975 ();
 b15zdnd11an1n64x5 FILLER_135_1039 ();
 b15zdnd11an1n64x5 FILLER_135_1103 ();
 b15zdnd11an1n64x5 FILLER_135_1167 ();
 b15zdnd11an1n64x5 FILLER_135_1231 ();
 b15zdnd11an1n64x5 FILLER_135_1295 ();
 b15zdnd11an1n64x5 FILLER_135_1359 ();
 b15zdnd11an1n32x5 FILLER_135_1423 ();
 b15zdnd11an1n16x5 FILLER_135_1455 ();
 b15zdnd11an1n08x5 FILLER_135_1471 ();
 b15zdnd11an1n04x5 FILLER_135_1479 ();
 b15zdnd00an1n02x5 FILLER_135_1483 ();
 b15zdnd00an1n01x5 FILLER_135_1485 ();
 b15zdnd11an1n16x5 FILLER_135_2257 ();
 b15zdnd11an1n08x5 FILLER_135_2273 ();
 b15zdnd00an1n02x5 FILLER_135_2281 ();
 b15zdnd00an1n01x5 FILLER_135_2283 ();
 b15zdnd11an1n16x5 FILLER_136_8 ();
 b15zdnd00an1n02x5 FILLER_136_24 ();
 b15zdnd00an1n01x5 FILLER_136_26 ();
 b15zdnd11an1n64x5 FILLER_136_34 ();
 b15zdnd11an1n64x5 FILLER_136_98 ();
 b15zdnd11an1n64x5 FILLER_136_162 ();
 b15zdnd11an1n64x5 FILLER_136_226 ();
 b15zdnd11an1n64x5 FILLER_136_290 ();
 b15zdnd11an1n32x5 FILLER_136_354 ();
 b15zdnd11an1n16x5 FILLER_136_386 ();
 b15zdnd11an1n08x5 FILLER_136_402 ();
 b15zdnd00an1n02x5 FILLER_136_410 ();
 b15zdnd11an1n64x5 FILLER_136_434 ();
 b15zdnd11an1n64x5 FILLER_136_498 ();
 b15zdnd11an1n64x5 FILLER_136_562 ();
 b15zdnd11an1n64x5 FILLER_136_626 ();
 b15zdnd11an1n16x5 FILLER_136_690 ();
 b15zdnd11an1n08x5 FILLER_136_706 ();
 b15zdnd11an1n04x5 FILLER_136_714 ();
 b15zdnd11an1n64x5 FILLER_136_726 ();
 b15zdnd11an1n64x5 FILLER_136_790 ();
 b15zdnd11an1n64x5 FILLER_136_854 ();
 b15zdnd11an1n64x5 FILLER_136_918 ();
 b15zdnd11an1n64x5 FILLER_136_982 ();
 b15zdnd11an1n64x5 FILLER_136_1046 ();
 b15zdnd11an1n64x5 FILLER_136_1110 ();
 b15zdnd11an1n64x5 FILLER_136_1174 ();
 b15zdnd11an1n64x5 FILLER_136_1238 ();
 b15zdnd11an1n64x5 FILLER_136_1302 ();
 b15zdnd11an1n64x5 FILLER_136_1366 ();
 b15zdnd11an1n32x5 FILLER_136_1430 ();
 b15zdnd11an1n16x5 FILLER_136_1462 ();
 b15zdnd11an1n08x5 FILLER_136_2265 ();
 b15zdnd00an1n02x5 FILLER_136_2273 ();
 b15zdnd00an1n01x5 FILLER_136_2275 ();
 b15zdnd11an1n08x5 FILLER_137_0 ();
 b15zdnd11an1n04x5 FILLER_137_8 ();
 b15zdnd00an1n02x5 FILLER_137_12 ();
 b15zdnd11an1n64x5 FILLER_137_22 ();
 b15zdnd11an1n64x5 FILLER_137_86 ();
 b15zdnd11an1n64x5 FILLER_137_150 ();
 b15zdnd11an1n64x5 FILLER_137_214 ();
 b15zdnd11an1n64x5 FILLER_137_278 ();
 b15zdnd11an1n64x5 FILLER_137_342 ();
 b15zdnd11an1n04x5 FILLER_137_406 ();
 b15zdnd00an1n02x5 FILLER_137_410 ();
 b15zdnd11an1n64x5 FILLER_137_422 ();
 b15zdnd11an1n64x5 FILLER_137_486 ();
 b15zdnd11an1n64x5 FILLER_137_550 ();
 b15zdnd11an1n64x5 FILLER_137_614 ();
 b15zdnd11an1n64x5 FILLER_137_678 ();
 b15zdnd11an1n64x5 FILLER_137_742 ();
 b15zdnd11an1n64x5 FILLER_137_806 ();
 b15zdnd11an1n64x5 FILLER_137_870 ();
 b15zdnd11an1n64x5 FILLER_137_934 ();
 b15zdnd11an1n64x5 FILLER_137_998 ();
 b15zdnd11an1n64x5 FILLER_137_1062 ();
 b15zdnd11an1n64x5 FILLER_137_1126 ();
 b15zdnd11an1n16x5 FILLER_137_1190 ();
 b15zdnd11an1n08x5 FILLER_137_1206 ();
 b15zdnd11an1n04x5 FILLER_137_1214 ();
 b15zdnd11an1n64x5 FILLER_137_1221 ();
 b15zdnd11an1n64x5 FILLER_137_1285 ();
 b15zdnd11an1n64x5 FILLER_137_1349 ();
 b15zdnd11an1n64x5 FILLER_137_1413 ();
 b15zdnd11an1n08x5 FILLER_137_1477 ();
 b15zdnd00an1n01x5 FILLER_137_1485 ();
 b15zdnd11an1n16x5 FILLER_137_2257 ();
 b15zdnd11an1n08x5 FILLER_137_2273 ();
 b15zdnd00an1n02x5 FILLER_137_2281 ();
 b15zdnd00an1n01x5 FILLER_137_2283 ();
 b15zdnd11an1n64x5 FILLER_138_8 ();
 b15zdnd11an1n64x5 FILLER_138_72 ();
 b15zdnd11an1n64x5 FILLER_138_136 ();
 b15zdnd11an1n64x5 FILLER_138_200 ();
 b15zdnd11an1n64x5 FILLER_138_264 ();
 b15zdnd11an1n64x5 FILLER_138_328 ();
 b15zdnd11an1n64x5 FILLER_138_392 ();
 b15zdnd11an1n08x5 FILLER_138_456 ();
 b15zdnd11an1n64x5 FILLER_138_476 ();
 b15zdnd11an1n64x5 FILLER_138_540 ();
 b15zdnd11an1n64x5 FILLER_138_604 ();
 b15zdnd11an1n32x5 FILLER_138_668 ();
 b15zdnd11an1n16x5 FILLER_138_700 ();
 b15zdnd00an1n02x5 FILLER_138_716 ();
 b15zdnd11an1n64x5 FILLER_138_726 ();
 b15zdnd11an1n64x5 FILLER_138_790 ();
 b15zdnd11an1n64x5 FILLER_138_854 ();
 b15zdnd11an1n64x5 FILLER_138_918 ();
 b15zdnd11an1n64x5 FILLER_138_982 ();
 b15zdnd11an1n64x5 FILLER_138_1046 ();
 b15zdnd11an1n64x5 FILLER_138_1110 ();
 b15zdnd11an1n32x5 FILLER_138_1174 ();
 b15zdnd11an1n08x5 FILLER_138_1206 ();
 b15zdnd11an1n04x5 FILLER_138_1214 ();
 b15zdnd11an1n08x5 FILLER_138_1221 ();
 b15zdnd00an1n01x5 FILLER_138_1229 ();
 b15zdnd11an1n64x5 FILLER_138_1233 ();
 b15zdnd11an1n64x5 FILLER_138_1297 ();
 b15zdnd11an1n64x5 FILLER_138_1361 ();
 b15zdnd11an1n32x5 FILLER_138_1425 ();
 b15zdnd11an1n16x5 FILLER_138_1457 ();
 b15zdnd11an1n04x5 FILLER_138_1473 ();
 b15zdnd00an1n01x5 FILLER_138_1477 ();
 b15zdnd00an1n02x5 FILLER_138_2265 ();
 b15zdnd00an1n01x5 FILLER_138_2267 ();
 b15zdnd00an1n02x5 FILLER_138_2274 ();
 b15zdnd11an1n16x5 FILLER_139_0 ();
 b15zdnd00an1n01x5 FILLER_139_16 ();
 b15zdnd11an1n64x5 FILLER_139_28 ();
 b15zdnd11an1n64x5 FILLER_139_92 ();
 b15zdnd11an1n64x5 FILLER_139_156 ();
 b15zdnd11an1n64x5 FILLER_139_220 ();
 b15zdnd11an1n64x5 FILLER_139_284 ();
 b15zdnd11an1n64x5 FILLER_139_348 ();
 b15zdnd11an1n64x5 FILLER_139_412 ();
 b15zdnd11an1n64x5 FILLER_139_476 ();
 b15zdnd11an1n64x5 FILLER_139_540 ();
 b15zdnd11an1n64x5 FILLER_139_604 ();
 b15zdnd11an1n64x5 FILLER_139_668 ();
 b15zdnd11an1n04x5 FILLER_139_732 ();
 b15zdnd00an1n02x5 FILLER_139_736 ();
 b15zdnd11an1n64x5 FILLER_139_747 ();
 b15zdnd11an1n64x5 FILLER_139_811 ();
 b15zdnd11an1n64x5 FILLER_139_875 ();
 b15zdnd11an1n64x5 FILLER_139_939 ();
 b15zdnd11an1n64x5 FILLER_139_1003 ();
 b15zdnd11an1n64x5 FILLER_139_1067 ();
 b15zdnd11an1n64x5 FILLER_139_1131 ();
 b15zdnd11an1n64x5 FILLER_139_1247 ();
 b15zdnd11an1n64x5 FILLER_139_1311 ();
 b15zdnd11an1n64x5 FILLER_139_1375 ();
 b15zdnd11an1n32x5 FILLER_139_1439 ();
 b15zdnd11an1n08x5 FILLER_139_1471 ();
 b15zdnd11an1n04x5 FILLER_139_1479 ();
 b15zdnd00an1n02x5 FILLER_139_1483 ();
 b15zdnd00an1n01x5 FILLER_139_1485 ();
 b15zdnd11an1n16x5 FILLER_139_2257 ();
 b15zdnd11an1n08x5 FILLER_139_2273 ();
 b15zdnd00an1n02x5 FILLER_139_2281 ();
 b15zdnd00an1n01x5 FILLER_139_2283 ();
 b15zdnd11an1n08x5 FILLER_140_8 ();
 b15zdnd11an1n04x5 FILLER_140_16 ();
 b15zdnd00an1n02x5 FILLER_140_20 ();
 b15zdnd00an1n01x5 FILLER_140_22 ();
 b15zdnd11an1n04x5 FILLER_140_30 ();
 b15zdnd11an1n64x5 FILLER_140_45 ();
 b15zdnd11an1n64x5 FILLER_140_109 ();
 b15zdnd11an1n64x5 FILLER_140_173 ();
 b15zdnd11an1n64x5 FILLER_140_237 ();
 b15zdnd11an1n64x5 FILLER_140_301 ();
 b15zdnd11an1n32x5 FILLER_140_365 ();
 b15zdnd11an1n16x5 FILLER_140_397 ();
 b15zdnd00an1n02x5 FILLER_140_413 ();
 b15zdnd00an1n01x5 FILLER_140_415 ();
 b15zdnd11an1n64x5 FILLER_140_437 ();
 b15zdnd11an1n64x5 FILLER_140_501 ();
 b15zdnd11an1n64x5 FILLER_140_565 ();
 b15zdnd11an1n32x5 FILLER_140_629 ();
 b15zdnd11an1n16x5 FILLER_140_661 ();
 b15zdnd11an1n08x5 FILLER_140_677 ();
 b15zdnd11an1n04x5 FILLER_140_685 ();
 b15zdnd00an1n02x5 FILLER_140_689 ();
 b15zdnd00an1n02x5 FILLER_140_716 ();
 b15zdnd00an1n02x5 FILLER_140_726 ();
 b15zdnd11an1n64x5 FILLER_140_772 ();
 b15zdnd11an1n64x5 FILLER_140_836 ();
 b15zdnd11an1n64x5 FILLER_140_900 ();
 b15zdnd11an1n64x5 FILLER_140_964 ();
 b15zdnd11an1n32x5 FILLER_140_1028 ();
 b15zdnd11an1n16x5 FILLER_140_1060 ();
 b15zdnd11an1n08x5 FILLER_140_1076 ();
 b15zdnd00an1n02x5 FILLER_140_1084 ();
 b15zdnd00an1n01x5 FILLER_140_1086 ();
 b15zdnd11an1n64x5 FILLER_140_1129 ();
 b15zdnd11an1n32x5 FILLER_140_1193 ();
 b15zdnd11an1n16x5 FILLER_140_1225 ();
 b15zdnd11an1n64x5 FILLER_140_1248 ();
 b15zdnd11an1n64x5 FILLER_140_1312 ();
 b15zdnd11an1n64x5 FILLER_140_1376 ();
 b15zdnd11an1n32x5 FILLER_140_1440 ();
 b15zdnd11an1n04x5 FILLER_140_1472 ();
 b15zdnd00an1n02x5 FILLER_140_1476 ();
 b15zdnd11an1n08x5 FILLER_140_2265 ();
 b15zdnd00an1n02x5 FILLER_140_2273 ();
 b15zdnd00an1n01x5 FILLER_140_2275 ();
 b15zdnd11an1n64x5 FILLER_141_0 ();
 b15zdnd11an1n64x5 FILLER_141_64 ();
 b15zdnd11an1n64x5 FILLER_141_128 ();
 b15zdnd11an1n64x5 FILLER_141_192 ();
 b15zdnd11an1n64x5 FILLER_141_256 ();
 b15zdnd11an1n64x5 FILLER_141_320 ();
 b15zdnd11an1n64x5 FILLER_141_384 ();
 b15zdnd11an1n64x5 FILLER_141_448 ();
 b15zdnd11an1n64x5 FILLER_141_512 ();
 b15zdnd11an1n64x5 FILLER_141_576 ();
 b15zdnd11an1n64x5 FILLER_141_640 ();
 b15zdnd11an1n16x5 FILLER_141_704 ();
 b15zdnd00an1n02x5 FILLER_141_720 ();
 b15zdnd11an1n64x5 FILLER_141_766 ();
 b15zdnd11an1n64x5 FILLER_141_830 ();
 b15zdnd11an1n64x5 FILLER_141_894 ();
 b15zdnd11an1n64x5 FILLER_141_958 ();
 b15zdnd11an1n64x5 FILLER_141_1022 ();
 b15zdnd11an1n64x5 FILLER_141_1086 ();
 b15zdnd11an1n64x5 FILLER_141_1150 ();
 b15zdnd11an1n64x5 FILLER_141_1214 ();
 b15zdnd11an1n64x5 FILLER_141_1278 ();
 b15zdnd11an1n64x5 FILLER_141_1342 ();
 b15zdnd11an1n64x5 FILLER_141_1406 ();
 b15zdnd11an1n16x5 FILLER_141_1470 ();
 b15zdnd11an1n16x5 FILLER_141_2257 ();
 b15zdnd11an1n08x5 FILLER_141_2273 ();
 b15zdnd00an1n02x5 FILLER_141_2281 ();
 b15zdnd00an1n01x5 FILLER_141_2283 ();
 b15zdnd11an1n64x5 FILLER_142_8 ();
 b15zdnd11an1n64x5 FILLER_142_72 ();
 b15zdnd11an1n64x5 FILLER_142_136 ();
 b15zdnd11an1n64x5 FILLER_142_200 ();
 b15zdnd11an1n64x5 FILLER_142_264 ();
 b15zdnd11an1n64x5 FILLER_142_328 ();
 b15zdnd11an1n64x5 FILLER_142_392 ();
 b15zdnd11an1n64x5 FILLER_142_456 ();
 b15zdnd11an1n64x5 FILLER_142_520 ();
 b15zdnd11an1n64x5 FILLER_142_584 ();
 b15zdnd11an1n32x5 FILLER_142_648 ();
 b15zdnd00an1n02x5 FILLER_142_680 ();
 b15zdnd11an1n04x5 FILLER_142_685 ();
 b15zdnd00an1n02x5 FILLER_142_716 ();
 b15zdnd00an1n02x5 FILLER_142_726 ();
 b15zdnd11an1n32x5 FILLER_142_772 ();
 b15zdnd11an1n04x5 FILLER_142_804 ();
 b15zdnd00an1n01x5 FILLER_142_808 ();
 b15zdnd11an1n64x5 FILLER_142_851 ();
 b15zdnd11an1n64x5 FILLER_142_915 ();
 b15zdnd11an1n32x5 FILLER_142_979 ();
 b15zdnd11an1n08x5 FILLER_142_1011 ();
 b15zdnd11an1n64x5 FILLER_142_1061 ();
 b15zdnd11an1n64x5 FILLER_142_1125 ();
 b15zdnd11an1n64x5 FILLER_142_1189 ();
 b15zdnd11an1n64x5 FILLER_142_1253 ();
 b15zdnd11an1n64x5 FILLER_142_1317 ();
 b15zdnd11an1n64x5 FILLER_142_1381 ();
 b15zdnd11an1n32x5 FILLER_142_1445 ();
 b15zdnd00an1n01x5 FILLER_142_1477 ();
 b15zdnd11an1n08x5 FILLER_142_2265 ();
 b15zdnd00an1n02x5 FILLER_142_2273 ();
 b15zdnd00an1n01x5 FILLER_142_2275 ();
 b15zdnd11an1n64x5 FILLER_143_0 ();
 b15zdnd11an1n64x5 FILLER_143_64 ();
 b15zdnd11an1n64x5 FILLER_143_128 ();
 b15zdnd11an1n64x5 FILLER_143_192 ();
 b15zdnd11an1n64x5 FILLER_143_256 ();
 b15zdnd11an1n64x5 FILLER_143_320 ();
 b15zdnd11an1n32x5 FILLER_143_384 ();
 b15zdnd00an1n01x5 FILLER_143_416 ();
 b15zdnd11an1n64x5 FILLER_143_437 ();
 b15zdnd11an1n64x5 FILLER_143_501 ();
 b15zdnd11an1n64x5 FILLER_143_565 ();
 b15zdnd11an1n32x5 FILLER_143_629 ();
 b15zdnd11an1n16x5 FILLER_143_661 ();
 b15zdnd11an1n08x5 FILLER_143_677 ();
 b15zdnd11an1n04x5 FILLER_143_685 ();
 b15zdnd11an1n04x5 FILLER_143_692 ();
 b15zdnd11an1n16x5 FILLER_143_699 ();
 b15zdnd11an1n04x5 FILLER_143_715 ();
 b15zdnd00an1n02x5 FILLER_143_719 ();
 b15zdnd00an1n01x5 FILLER_143_721 ();
 b15zdnd11an1n04x5 FILLER_143_766 ();
 b15zdnd11an1n64x5 FILLER_143_773 ();
 b15zdnd11an1n64x5 FILLER_143_837 ();
 b15zdnd11an1n64x5 FILLER_143_901 ();
 b15zdnd11an1n64x5 FILLER_143_965 ();
 b15zdnd11an1n64x5 FILLER_143_1029 ();
 b15zdnd11an1n64x5 FILLER_143_1093 ();
 b15zdnd11an1n64x5 FILLER_143_1157 ();
 b15zdnd11an1n64x5 FILLER_143_1221 ();
 b15zdnd11an1n64x5 FILLER_143_1285 ();
 b15zdnd11an1n64x5 FILLER_143_1349 ();
 b15zdnd11an1n64x5 FILLER_143_1413 ();
 b15zdnd11an1n08x5 FILLER_143_1477 ();
 b15zdnd00an1n01x5 FILLER_143_1485 ();
 b15zdnd11an1n16x5 FILLER_143_2257 ();
 b15zdnd11an1n08x5 FILLER_143_2273 ();
 b15zdnd00an1n02x5 FILLER_143_2281 ();
 b15zdnd00an1n01x5 FILLER_143_2283 ();
 b15zdnd11an1n64x5 FILLER_144_8 ();
 b15zdnd11an1n64x5 FILLER_144_72 ();
 b15zdnd11an1n64x5 FILLER_144_136 ();
 b15zdnd11an1n64x5 FILLER_144_200 ();
 b15zdnd11an1n64x5 FILLER_144_264 ();
 b15zdnd11an1n64x5 FILLER_144_328 ();
 b15zdnd11an1n64x5 FILLER_144_392 ();
 b15zdnd11an1n08x5 FILLER_144_456 ();
 b15zdnd11an1n04x5 FILLER_144_464 ();
 b15zdnd11an1n64x5 FILLER_144_480 ();
 b15zdnd11an1n64x5 FILLER_144_544 ();
 b15zdnd11an1n64x5 FILLER_144_608 ();
 b15zdnd11an1n32x5 FILLER_144_672 ();
 b15zdnd11an1n08x5 FILLER_144_704 ();
 b15zdnd11an1n04x5 FILLER_144_712 ();
 b15zdnd00an1n02x5 FILLER_144_716 ();
 b15zdnd00an1n02x5 FILLER_144_726 ();
 b15zdnd11an1n08x5 FILLER_144_737 ();
 b15zdnd00an1n01x5 FILLER_144_745 ();
 b15zdnd11an1n04x5 FILLER_144_749 ();
 b15zdnd11an1n04x5 FILLER_144_756 ();
 b15zdnd11an1n64x5 FILLER_144_763 ();
 b15zdnd11an1n64x5 FILLER_144_827 ();
 b15zdnd11an1n64x5 FILLER_144_891 ();
 b15zdnd11an1n64x5 FILLER_144_955 ();
 b15zdnd11an1n64x5 FILLER_144_1019 ();
 b15zdnd11an1n64x5 FILLER_144_1083 ();
 b15zdnd11an1n64x5 FILLER_144_1147 ();
 b15zdnd11an1n64x5 FILLER_144_1211 ();
 b15zdnd11an1n32x5 FILLER_144_1275 ();
 b15zdnd11an1n04x5 FILLER_144_1307 ();
 b15zdnd00an1n01x5 FILLER_144_1311 ();
 b15zdnd11an1n04x5 FILLER_144_1315 ();
 b15zdnd11an1n64x5 FILLER_144_1322 ();
 b15zdnd11an1n64x5 FILLER_144_1386 ();
 b15zdnd11an1n16x5 FILLER_144_1450 ();
 b15zdnd11an1n08x5 FILLER_144_1466 ();
 b15zdnd11an1n04x5 FILLER_144_1474 ();
 b15zdnd11an1n08x5 FILLER_144_2265 ();
 b15zdnd00an1n02x5 FILLER_144_2273 ();
 b15zdnd00an1n01x5 FILLER_144_2275 ();
 b15zdnd11an1n64x5 FILLER_145_0 ();
 b15zdnd11an1n64x5 FILLER_145_64 ();
 b15zdnd11an1n64x5 FILLER_145_128 ();
 b15zdnd11an1n64x5 FILLER_145_192 ();
 b15zdnd11an1n64x5 FILLER_145_256 ();
 b15zdnd11an1n64x5 FILLER_145_320 ();
 b15zdnd11an1n64x5 FILLER_145_384 ();
 b15zdnd11an1n64x5 FILLER_145_448 ();
 b15zdnd11an1n64x5 FILLER_145_512 ();
 b15zdnd11an1n64x5 FILLER_145_576 ();
 b15zdnd11an1n64x5 FILLER_145_640 ();
 b15zdnd11an1n16x5 FILLER_145_704 ();
 b15zdnd11an1n08x5 FILLER_145_720 ();
 b15zdnd11an1n04x5 FILLER_145_728 ();
 b15zdnd11an1n04x5 FILLER_145_735 ();
 b15zdnd11an1n04x5 FILLER_145_742 ();
 b15zdnd11an1n04x5 FILLER_145_749 ();
 b15zdnd11an1n04x5 FILLER_145_756 ();
 b15zdnd11an1n64x5 FILLER_145_763 ();
 b15zdnd11an1n64x5 FILLER_145_827 ();
 b15zdnd11an1n64x5 FILLER_145_891 ();
 b15zdnd11an1n64x5 FILLER_145_955 ();
 b15zdnd00an1n01x5 FILLER_145_1019 ();
 b15zdnd11an1n64x5 FILLER_145_1062 ();
 b15zdnd11an1n64x5 FILLER_145_1126 ();
 b15zdnd11an1n64x5 FILLER_145_1190 ();
 b15zdnd11an1n32x5 FILLER_145_1254 ();
 b15zdnd11an1n16x5 FILLER_145_1286 ();
 b15zdnd11an1n08x5 FILLER_145_1302 ();
 b15zdnd11an1n04x5 FILLER_145_1310 ();
 b15zdnd00an1n02x5 FILLER_145_1314 ();
 b15zdnd00an1n01x5 FILLER_145_1316 ();
 b15zdnd11an1n64x5 FILLER_145_1342 ();
 b15zdnd11an1n64x5 FILLER_145_1406 ();
 b15zdnd11an1n16x5 FILLER_145_1470 ();
 b15zdnd11an1n16x5 FILLER_145_2257 ();
 b15zdnd11an1n08x5 FILLER_145_2273 ();
 b15zdnd00an1n02x5 FILLER_145_2281 ();
 b15zdnd00an1n01x5 FILLER_145_2283 ();
 b15zdnd11an1n64x5 FILLER_146_8 ();
 b15zdnd11an1n64x5 FILLER_146_72 ();
 b15zdnd11an1n64x5 FILLER_146_136 ();
 b15zdnd11an1n64x5 FILLER_146_200 ();
 b15zdnd11an1n64x5 FILLER_146_264 ();
 b15zdnd11an1n64x5 FILLER_146_328 ();
 b15zdnd11an1n64x5 FILLER_146_392 ();
 b15zdnd11an1n64x5 FILLER_146_456 ();
 b15zdnd11an1n64x5 FILLER_146_520 ();
 b15zdnd11an1n64x5 FILLER_146_584 ();
 b15zdnd11an1n64x5 FILLER_146_648 ();
 b15zdnd11an1n04x5 FILLER_146_712 ();
 b15zdnd00an1n02x5 FILLER_146_716 ();
 b15zdnd11an1n04x5 FILLER_146_726 ();
 b15zdnd00an1n02x5 FILLER_146_730 ();
 b15zdnd11an1n08x5 FILLER_146_735 ();
 b15zdnd00an1n02x5 FILLER_146_743 ();
 b15zdnd11an1n04x5 FILLER_146_748 ();
 b15zdnd11an1n64x5 FILLER_146_755 ();
 b15zdnd11an1n64x5 FILLER_146_819 ();
 b15zdnd11an1n64x5 FILLER_146_883 ();
 b15zdnd11an1n64x5 FILLER_146_947 ();
 b15zdnd11an1n64x5 FILLER_146_1011 ();
 b15zdnd11an1n64x5 FILLER_146_1075 ();
 b15zdnd11an1n64x5 FILLER_146_1139 ();
 b15zdnd11an1n64x5 FILLER_146_1203 ();
 b15zdnd11an1n32x5 FILLER_146_1267 ();
 b15zdnd11an1n16x5 FILLER_146_1299 ();
 b15zdnd11an1n08x5 FILLER_146_1315 ();
 b15zdnd11an1n04x5 FILLER_146_1323 ();
 b15zdnd00an1n01x5 FILLER_146_1327 ();
 b15zdnd11an1n04x5 FILLER_146_1331 ();
 b15zdnd11an1n64x5 FILLER_146_1338 ();
 b15zdnd11an1n64x5 FILLER_146_1402 ();
 b15zdnd11an1n08x5 FILLER_146_1466 ();
 b15zdnd11an1n04x5 FILLER_146_1474 ();
 b15zdnd11an1n08x5 FILLER_146_2265 ();
 b15zdnd00an1n02x5 FILLER_146_2273 ();
 b15zdnd00an1n01x5 FILLER_146_2275 ();
 b15zdnd11an1n64x5 FILLER_147_0 ();
 b15zdnd11an1n64x5 FILLER_147_64 ();
 b15zdnd11an1n64x5 FILLER_147_128 ();
 b15zdnd11an1n64x5 FILLER_147_192 ();
 b15zdnd11an1n64x5 FILLER_147_256 ();
 b15zdnd11an1n64x5 FILLER_147_320 ();
 b15zdnd11an1n64x5 FILLER_147_384 ();
 b15zdnd11an1n64x5 FILLER_147_448 ();
 b15zdnd11an1n64x5 FILLER_147_512 ();
 b15zdnd11an1n64x5 FILLER_147_576 ();
 b15zdnd11an1n64x5 FILLER_147_640 ();
 b15zdnd11an1n64x5 FILLER_147_704 ();
 b15zdnd11an1n64x5 FILLER_147_768 ();
 b15zdnd11an1n64x5 FILLER_147_832 ();
 b15zdnd11an1n64x5 FILLER_147_896 ();
 b15zdnd11an1n64x5 FILLER_147_960 ();
 b15zdnd11an1n64x5 FILLER_147_1024 ();
 b15zdnd11an1n32x5 FILLER_147_1088 ();
 b15zdnd11an1n16x5 FILLER_147_1120 ();
 b15zdnd11an1n04x5 FILLER_147_1136 ();
 b15zdnd00an1n02x5 FILLER_147_1140 ();
 b15zdnd11an1n08x5 FILLER_147_1145 ();
 b15zdnd11an1n04x5 FILLER_147_1153 ();
 b15zdnd00an1n01x5 FILLER_147_1157 ();
 b15zdnd11an1n32x5 FILLER_147_1166 ();
 b15zdnd11an1n08x5 FILLER_147_1198 ();
 b15zdnd11an1n04x5 FILLER_147_1206 ();
 b15zdnd00an1n01x5 FILLER_147_1210 ();
 b15zdnd11an1n16x5 FILLER_147_1221 ();
 b15zdnd11an1n04x5 FILLER_147_1237 ();
 b15zdnd00an1n02x5 FILLER_147_1241 ();
 b15zdnd00an1n01x5 FILLER_147_1243 ();
 b15zdnd11an1n64x5 FILLER_147_1254 ();
 b15zdnd11an1n08x5 FILLER_147_1318 ();
 b15zdnd00an1n02x5 FILLER_147_1326 ();
 b15zdnd00an1n01x5 FILLER_147_1328 ();
 b15zdnd11an1n64x5 FILLER_147_1364 ();
 b15zdnd11an1n32x5 FILLER_147_1428 ();
 b15zdnd11an1n16x5 FILLER_147_1460 ();
 b15zdnd11an1n08x5 FILLER_147_1476 ();
 b15zdnd00an1n02x5 FILLER_147_1484 ();
 b15zdnd11an1n16x5 FILLER_147_2257 ();
 b15zdnd11an1n08x5 FILLER_147_2273 ();
 b15zdnd00an1n02x5 FILLER_147_2281 ();
 b15zdnd00an1n01x5 FILLER_147_2283 ();
 b15zdnd11an1n64x5 FILLER_148_8 ();
 b15zdnd11an1n64x5 FILLER_148_72 ();
 b15zdnd11an1n64x5 FILLER_148_136 ();
 b15zdnd11an1n64x5 FILLER_148_200 ();
 b15zdnd11an1n64x5 FILLER_148_264 ();
 b15zdnd11an1n64x5 FILLER_148_328 ();
 b15zdnd11an1n64x5 FILLER_148_392 ();
 b15zdnd11an1n04x5 FILLER_148_456 ();
 b15zdnd00an1n01x5 FILLER_148_460 ();
 b15zdnd11an1n64x5 FILLER_148_470 ();
 b15zdnd11an1n64x5 FILLER_148_534 ();
 b15zdnd11an1n64x5 FILLER_148_598 ();
 b15zdnd11an1n32x5 FILLER_148_662 ();
 b15zdnd11an1n16x5 FILLER_148_694 ();
 b15zdnd11an1n08x5 FILLER_148_710 ();
 b15zdnd11an1n64x5 FILLER_148_726 ();
 b15zdnd11an1n64x5 FILLER_148_790 ();
 b15zdnd11an1n64x5 FILLER_148_854 ();
 b15zdnd11an1n64x5 FILLER_148_918 ();
 b15zdnd11an1n64x5 FILLER_148_982 ();
 b15zdnd11an1n64x5 FILLER_148_1046 ();
 b15zdnd11an1n16x5 FILLER_148_1110 ();
 b15zdnd11an1n08x5 FILLER_148_1126 ();
 b15zdnd11an1n04x5 FILLER_148_1134 ();
 b15zdnd00an1n02x5 FILLER_148_1138 ();
 b15zdnd00an1n01x5 FILLER_148_1140 ();
 b15zdnd11an1n04x5 FILLER_148_1144 ();
 b15zdnd11an1n08x5 FILLER_148_1151 ();
 b15zdnd11an1n04x5 FILLER_148_1159 ();
 b15zdnd00an1n01x5 FILLER_148_1163 ();
 b15zdnd11an1n64x5 FILLER_148_1206 ();
 b15zdnd11an1n64x5 FILLER_148_1270 ();
 b15zdnd11an1n64x5 FILLER_148_1334 ();
 b15zdnd11an1n64x5 FILLER_148_1398 ();
 b15zdnd11an1n16x5 FILLER_148_1462 ();
 b15zdnd00an1n02x5 FILLER_148_2265 ();
 b15zdnd00an1n01x5 FILLER_148_2267 ();
 b15zdnd00an1n02x5 FILLER_148_2274 ();
 b15zdnd11an1n64x5 FILLER_149_0 ();
 b15zdnd11an1n64x5 FILLER_149_64 ();
 b15zdnd11an1n64x5 FILLER_149_128 ();
 b15zdnd11an1n64x5 FILLER_149_192 ();
 b15zdnd11an1n64x5 FILLER_149_256 ();
 b15zdnd11an1n64x5 FILLER_149_320 ();
 b15zdnd11an1n64x5 FILLER_149_384 ();
 b15zdnd00an1n02x5 FILLER_149_448 ();
 b15zdnd00an1n01x5 FILLER_149_450 ();
 b15zdnd11an1n64x5 FILLER_149_493 ();
 b15zdnd11an1n64x5 FILLER_149_557 ();
 b15zdnd11an1n64x5 FILLER_149_621 ();
 b15zdnd11an1n64x5 FILLER_149_685 ();
 b15zdnd11an1n64x5 FILLER_149_749 ();
 b15zdnd11an1n64x5 FILLER_149_813 ();
 b15zdnd11an1n64x5 FILLER_149_877 ();
 b15zdnd11an1n64x5 FILLER_149_941 ();
 b15zdnd11an1n64x5 FILLER_149_1005 ();
 b15zdnd11an1n32x5 FILLER_149_1069 ();
 b15zdnd11an1n16x5 FILLER_149_1101 ();
 b15zdnd00an1n01x5 FILLER_149_1117 ();
 b15zdnd11an1n64x5 FILLER_149_1170 ();
 b15zdnd11an1n64x5 FILLER_149_1234 ();
 b15zdnd11an1n64x5 FILLER_149_1298 ();
 b15zdnd11an1n64x5 FILLER_149_1362 ();
 b15zdnd11an1n32x5 FILLER_149_1426 ();
 b15zdnd11an1n16x5 FILLER_149_1458 ();
 b15zdnd11an1n08x5 FILLER_149_1474 ();
 b15zdnd11an1n04x5 FILLER_149_1482 ();
 b15zdnd11an1n16x5 FILLER_149_2257 ();
 b15zdnd11an1n08x5 FILLER_149_2273 ();
 b15zdnd00an1n02x5 FILLER_149_2281 ();
 b15zdnd00an1n01x5 FILLER_149_2283 ();
 b15zdnd11an1n64x5 FILLER_150_8 ();
 b15zdnd11an1n64x5 FILLER_150_72 ();
 b15zdnd11an1n64x5 FILLER_150_136 ();
 b15zdnd11an1n64x5 FILLER_150_200 ();
 b15zdnd11an1n64x5 FILLER_150_264 ();
 b15zdnd11an1n64x5 FILLER_150_328 ();
 b15zdnd11an1n64x5 FILLER_150_392 ();
 b15zdnd11an1n64x5 FILLER_150_456 ();
 b15zdnd11an1n64x5 FILLER_150_520 ();
 b15zdnd11an1n64x5 FILLER_150_584 ();
 b15zdnd11an1n64x5 FILLER_150_648 ();
 b15zdnd11an1n04x5 FILLER_150_712 ();
 b15zdnd00an1n02x5 FILLER_150_716 ();
 b15zdnd11an1n64x5 FILLER_150_726 ();
 b15zdnd11an1n64x5 FILLER_150_790 ();
 b15zdnd11an1n64x5 FILLER_150_854 ();
 b15zdnd11an1n64x5 FILLER_150_918 ();
 b15zdnd11an1n64x5 FILLER_150_982 ();
 b15zdnd11an1n64x5 FILLER_150_1046 ();
 b15zdnd11an1n64x5 FILLER_150_1110 ();
 b15zdnd11an1n64x5 FILLER_150_1174 ();
 b15zdnd11an1n16x5 FILLER_150_1238 ();
 b15zdnd11an1n04x5 FILLER_150_1254 ();
 b15zdnd11an1n64x5 FILLER_150_1267 ();
 b15zdnd11an1n64x5 FILLER_150_1331 ();
 b15zdnd11an1n64x5 FILLER_150_1395 ();
 b15zdnd11an1n16x5 FILLER_150_1459 ();
 b15zdnd00an1n02x5 FILLER_150_1475 ();
 b15zdnd00an1n01x5 FILLER_150_1477 ();
 b15zdnd11an1n08x5 FILLER_150_2265 ();
 b15zdnd00an1n02x5 FILLER_150_2273 ();
 b15zdnd00an1n01x5 FILLER_150_2275 ();
 b15zdnd11an1n64x5 FILLER_151_0 ();
 b15zdnd11an1n64x5 FILLER_151_64 ();
 b15zdnd11an1n64x5 FILLER_151_128 ();
 b15zdnd11an1n64x5 FILLER_151_192 ();
 b15zdnd11an1n64x5 FILLER_151_256 ();
 b15zdnd11an1n64x5 FILLER_151_320 ();
 b15zdnd11an1n64x5 FILLER_151_384 ();
 b15zdnd11an1n64x5 FILLER_151_448 ();
 b15zdnd11an1n64x5 FILLER_151_512 ();
 b15zdnd11an1n64x5 FILLER_151_576 ();
 b15zdnd11an1n64x5 FILLER_151_640 ();
 b15zdnd11an1n16x5 FILLER_151_704 ();
 b15zdnd00an1n02x5 FILLER_151_720 ();
 b15zdnd00an1n01x5 FILLER_151_722 ();
 b15zdnd11an1n64x5 FILLER_151_765 ();
 b15zdnd11an1n64x5 FILLER_151_829 ();
 b15zdnd11an1n64x5 FILLER_151_893 ();
 b15zdnd11an1n64x5 FILLER_151_957 ();
 b15zdnd11an1n64x5 FILLER_151_1021 ();
 b15zdnd11an1n64x5 FILLER_151_1085 ();
 b15zdnd11an1n64x5 FILLER_151_1149 ();
 b15zdnd11an1n64x5 FILLER_151_1213 ();
 b15zdnd11an1n64x5 FILLER_151_1277 ();
 b15zdnd11an1n64x5 FILLER_151_1341 ();
 b15zdnd11an1n64x5 FILLER_151_1405 ();
 b15zdnd11an1n16x5 FILLER_151_1469 ();
 b15zdnd00an1n01x5 FILLER_151_1485 ();
 b15zdnd11an1n16x5 FILLER_151_2257 ();
 b15zdnd11an1n08x5 FILLER_151_2273 ();
 b15zdnd00an1n02x5 FILLER_151_2281 ();
 b15zdnd00an1n01x5 FILLER_151_2283 ();
 b15zdnd11an1n64x5 FILLER_152_8 ();
 b15zdnd11an1n64x5 FILLER_152_72 ();
 b15zdnd11an1n64x5 FILLER_152_136 ();
 b15zdnd11an1n64x5 FILLER_152_200 ();
 b15zdnd11an1n64x5 FILLER_152_264 ();
 b15zdnd11an1n64x5 FILLER_152_328 ();
 b15zdnd11an1n64x5 FILLER_152_392 ();
 b15zdnd11an1n32x5 FILLER_152_456 ();
 b15zdnd11an1n16x5 FILLER_152_488 ();
 b15zdnd11an1n08x5 FILLER_152_504 ();
 b15zdnd11an1n04x5 FILLER_152_512 ();
 b15zdnd00an1n02x5 FILLER_152_516 ();
 b15zdnd11an1n64x5 FILLER_152_534 ();
 b15zdnd11an1n64x5 FILLER_152_598 ();
 b15zdnd11an1n32x5 FILLER_152_662 ();
 b15zdnd11an1n16x5 FILLER_152_694 ();
 b15zdnd11an1n08x5 FILLER_152_710 ();
 b15zdnd11an1n64x5 FILLER_152_726 ();
 b15zdnd11an1n64x5 FILLER_152_790 ();
 b15zdnd11an1n64x5 FILLER_152_854 ();
 b15zdnd11an1n64x5 FILLER_152_918 ();
 b15zdnd11an1n64x5 FILLER_152_982 ();
 b15zdnd11an1n64x5 FILLER_152_1046 ();
 b15zdnd11an1n64x5 FILLER_152_1110 ();
 b15zdnd11an1n64x5 FILLER_152_1174 ();
 b15zdnd11an1n64x5 FILLER_152_1238 ();
 b15zdnd11an1n64x5 FILLER_152_1302 ();
 b15zdnd11an1n64x5 FILLER_152_1366 ();
 b15zdnd11an1n32x5 FILLER_152_1430 ();
 b15zdnd11an1n16x5 FILLER_152_1462 ();
 b15zdnd11an1n08x5 FILLER_152_2265 ();
 b15zdnd00an1n02x5 FILLER_152_2273 ();
 b15zdnd00an1n01x5 FILLER_152_2275 ();
 b15zdnd11an1n64x5 FILLER_153_0 ();
 b15zdnd11an1n64x5 FILLER_153_64 ();
 b15zdnd11an1n64x5 FILLER_153_128 ();
 b15zdnd11an1n64x5 FILLER_153_192 ();
 b15zdnd11an1n64x5 FILLER_153_256 ();
 b15zdnd11an1n64x5 FILLER_153_320 ();
 b15zdnd11an1n16x5 FILLER_153_384 ();
 b15zdnd11an1n08x5 FILLER_153_400 ();
 b15zdnd11an1n04x5 FILLER_153_408 ();
 b15zdnd00an1n02x5 FILLER_153_412 ();
 b15zdnd00an1n01x5 FILLER_153_414 ();
 b15zdnd11an1n64x5 FILLER_153_437 ();
 b15zdnd11an1n64x5 FILLER_153_501 ();
 b15zdnd11an1n64x5 FILLER_153_565 ();
 b15zdnd11an1n64x5 FILLER_153_629 ();
 b15zdnd11an1n64x5 FILLER_153_693 ();
 b15zdnd11an1n64x5 FILLER_153_757 ();
 b15zdnd11an1n64x5 FILLER_153_821 ();
 b15zdnd11an1n64x5 FILLER_153_885 ();
 b15zdnd11an1n64x5 FILLER_153_949 ();
 b15zdnd11an1n64x5 FILLER_153_1013 ();
 b15zdnd11an1n64x5 FILLER_153_1077 ();
 b15zdnd11an1n64x5 FILLER_153_1141 ();
 b15zdnd11an1n64x5 FILLER_153_1205 ();
 b15zdnd11an1n16x5 FILLER_153_1269 ();
 b15zdnd11an1n08x5 FILLER_153_1285 ();
 b15zdnd11an1n04x5 FILLER_153_1293 ();
 b15zdnd11an1n64x5 FILLER_153_1339 ();
 b15zdnd11an1n64x5 FILLER_153_1403 ();
 b15zdnd11an1n16x5 FILLER_153_1467 ();
 b15zdnd00an1n02x5 FILLER_153_1483 ();
 b15zdnd00an1n01x5 FILLER_153_1485 ();
 b15zdnd11an1n16x5 FILLER_153_2257 ();
 b15zdnd11an1n08x5 FILLER_153_2273 ();
 b15zdnd00an1n02x5 FILLER_153_2281 ();
 b15zdnd00an1n01x5 FILLER_153_2283 ();
 b15zdnd11an1n64x5 FILLER_154_8 ();
 b15zdnd11an1n64x5 FILLER_154_72 ();
 b15zdnd11an1n64x5 FILLER_154_136 ();
 b15zdnd11an1n64x5 FILLER_154_200 ();
 b15zdnd11an1n64x5 FILLER_154_264 ();
 b15zdnd11an1n64x5 FILLER_154_328 ();
 b15zdnd11an1n64x5 FILLER_154_392 ();
 b15zdnd11an1n64x5 FILLER_154_456 ();
 b15zdnd11an1n64x5 FILLER_154_520 ();
 b15zdnd11an1n64x5 FILLER_154_584 ();
 b15zdnd11an1n64x5 FILLER_154_648 ();
 b15zdnd11an1n04x5 FILLER_154_712 ();
 b15zdnd00an1n02x5 FILLER_154_716 ();
 b15zdnd11an1n64x5 FILLER_154_726 ();
 b15zdnd11an1n64x5 FILLER_154_790 ();
 b15zdnd11an1n64x5 FILLER_154_854 ();
 b15zdnd11an1n64x5 FILLER_154_918 ();
 b15zdnd11an1n64x5 FILLER_154_982 ();
 b15zdnd11an1n16x5 FILLER_154_1046 ();
 b15zdnd11an1n08x5 FILLER_154_1062 ();
 b15zdnd11an1n04x5 FILLER_154_1070 ();
 b15zdnd00an1n02x5 FILLER_154_1074 ();
 b15zdnd11an1n32x5 FILLER_154_1084 ();
 b15zdnd11an1n16x5 FILLER_154_1116 ();
 b15zdnd11an1n08x5 FILLER_154_1132 ();
 b15zdnd11an1n64x5 FILLER_154_1182 ();
 b15zdnd11an1n64x5 FILLER_154_1246 ();
 b15zdnd11an1n64x5 FILLER_154_1310 ();
 b15zdnd11an1n64x5 FILLER_154_1374 ();
 b15zdnd11an1n32x5 FILLER_154_1438 ();
 b15zdnd11an1n08x5 FILLER_154_1470 ();
 b15zdnd11an1n08x5 FILLER_154_2265 ();
 b15zdnd00an1n02x5 FILLER_154_2273 ();
 b15zdnd00an1n01x5 FILLER_154_2275 ();
 b15zdnd11an1n64x5 FILLER_155_0 ();
 b15zdnd11an1n64x5 FILLER_155_64 ();
 b15zdnd11an1n64x5 FILLER_155_128 ();
 b15zdnd11an1n64x5 FILLER_155_192 ();
 b15zdnd11an1n64x5 FILLER_155_256 ();
 b15zdnd11an1n64x5 FILLER_155_320 ();
 b15zdnd11an1n32x5 FILLER_155_384 ();
 b15zdnd11an1n04x5 FILLER_155_416 ();
 b15zdnd00an1n02x5 FILLER_155_420 ();
 b15zdnd11an1n64x5 FILLER_155_432 ();
 b15zdnd11an1n64x5 FILLER_155_496 ();
 b15zdnd11an1n64x5 FILLER_155_560 ();
 b15zdnd11an1n64x5 FILLER_155_624 ();
 b15zdnd11an1n64x5 FILLER_155_688 ();
 b15zdnd11an1n64x5 FILLER_155_752 ();
 b15zdnd11an1n64x5 FILLER_155_816 ();
 b15zdnd11an1n64x5 FILLER_155_880 ();
 b15zdnd11an1n64x5 FILLER_155_944 ();
 b15zdnd11an1n64x5 FILLER_155_1008 ();
 b15zdnd11an1n64x5 FILLER_155_1072 ();
 b15zdnd11an1n04x5 FILLER_155_1136 ();
 b15zdnd00an1n02x5 FILLER_155_1140 ();
 b15zdnd11an1n64x5 FILLER_155_1184 ();
 b15zdnd11an1n64x5 FILLER_155_1248 ();
 b15zdnd11an1n64x5 FILLER_155_1312 ();
 b15zdnd11an1n64x5 FILLER_155_1376 ();
 b15zdnd11an1n32x5 FILLER_155_1440 ();
 b15zdnd11an1n08x5 FILLER_155_1472 ();
 b15zdnd11an1n04x5 FILLER_155_1480 ();
 b15zdnd00an1n02x5 FILLER_155_1484 ();
 b15zdnd11an1n16x5 FILLER_155_2257 ();
 b15zdnd11an1n08x5 FILLER_155_2273 ();
 b15zdnd00an1n02x5 FILLER_155_2281 ();
 b15zdnd00an1n01x5 FILLER_155_2283 ();
 b15zdnd11an1n16x5 FILLER_156_8 ();
 b15zdnd00an1n01x5 FILLER_156_24 ();
 b15zdnd11an1n64x5 FILLER_156_36 ();
 b15zdnd11an1n64x5 FILLER_156_100 ();
 b15zdnd11an1n64x5 FILLER_156_164 ();
 b15zdnd11an1n64x5 FILLER_156_228 ();
 b15zdnd11an1n64x5 FILLER_156_292 ();
 b15zdnd11an1n64x5 FILLER_156_356 ();
 b15zdnd11an1n64x5 FILLER_156_420 ();
 b15zdnd11an1n64x5 FILLER_156_484 ();
 b15zdnd11an1n64x5 FILLER_156_548 ();
 b15zdnd11an1n64x5 FILLER_156_612 ();
 b15zdnd11an1n32x5 FILLER_156_676 ();
 b15zdnd11an1n08x5 FILLER_156_708 ();
 b15zdnd00an1n02x5 FILLER_156_716 ();
 b15zdnd11an1n64x5 FILLER_156_726 ();
 b15zdnd11an1n64x5 FILLER_156_790 ();
 b15zdnd11an1n64x5 FILLER_156_854 ();
 b15zdnd11an1n64x5 FILLER_156_918 ();
 b15zdnd11an1n64x5 FILLER_156_982 ();
 b15zdnd11an1n64x5 FILLER_156_1046 ();
 b15zdnd11an1n64x5 FILLER_156_1110 ();
 b15zdnd11an1n64x5 FILLER_156_1174 ();
 b15zdnd11an1n64x5 FILLER_156_1238 ();
 b15zdnd11an1n64x5 FILLER_156_1302 ();
 b15zdnd11an1n64x5 FILLER_156_1366 ();
 b15zdnd11an1n32x5 FILLER_156_1430 ();
 b15zdnd11an1n16x5 FILLER_156_1462 ();
 b15zdnd11an1n08x5 FILLER_156_2265 ();
 b15zdnd00an1n02x5 FILLER_156_2273 ();
 b15zdnd00an1n01x5 FILLER_156_2275 ();
 b15zdnd11an1n64x5 FILLER_157_0 ();
 b15zdnd11an1n64x5 FILLER_157_64 ();
 b15zdnd11an1n64x5 FILLER_157_128 ();
 b15zdnd11an1n64x5 FILLER_157_192 ();
 b15zdnd11an1n64x5 FILLER_157_256 ();
 b15zdnd11an1n64x5 FILLER_157_320 ();
 b15zdnd11an1n64x5 FILLER_157_384 ();
 b15zdnd11an1n64x5 FILLER_157_448 ();
 b15zdnd11an1n64x5 FILLER_157_512 ();
 b15zdnd11an1n64x5 FILLER_157_576 ();
 b15zdnd11an1n64x5 FILLER_157_640 ();
 b15zdnd11an1n64x5 FILLER_157_704 ();
 b15zdnd11an1n64x5 FILLER_157_768 ();
 b15zdnd11an1n64x5 FILLER_157_832 ();
 b15zdnd11an1n64x5 FILLER_157_896 ();
 b15zdnd11an1n64x5 FILLER_157_960 ();
 b15zdnd11an1n04x5 FILLER_157_1024 ();
 b15zdnd00an1n01x5 FILLER_157_1028 ();
 b15zdnd11an1n64x5 FILLER_157_1071 ();
 b15zdnd11an1n64x5 FILLER_157_1135 ();
 b15zdnd11an1n64x5 FILLER_157_1199 ();
 b15zdnd11an1n16x5 FILLER_157_1263 ();
 b15zdnd11an1n08x5 FILLER_157_1279 ();
 b15zdnd00an1n02x5 FILLER_157_1287 ();
 b15zdnd11an1n08x5 FILLER_157_1292 ();
 b15zdnd00an1n02x5 FILLER_157_1300 ();
 b15zdnd00an1n01x5 FILLER_157_1302 ();
 b15zdnd11an1n64x5 FILLER_157_1345 ();
 b15zdnd11an1n64x5 FILLER_157_1409 ();
 b15zdnd11an1n08x5 FILLER_157_1473 ();
 b15zdnd11an1n04x5 FILLER_157_1481 ();
 b15zdnd00an1n01x5 FILLER_157_1485 ();
 b15zdnd11an1n16x5 FILLER_157_2257 ();
 b15zdnd11an1n08x5 FILLER_157_2273 ();
 b15zdnd00an1n02x5 FILLER_157_2281 ();
 b15zdnd00an1n01x5 FILLER_157_2283 ();
 b15zdnd11an1n64x5 FILLER_158_8 ();
 b15zdnd11an1n64x5 FILLER_158_72 ();
 b15zdnd11an1n64x5 FILLER_158_136 ();
 b15zdnd11an1n64x5 FILLER_158_200 ();
 b15zdnd11an1n64x5 FILLER_158_264 ();
 b15zdnd11an1n64x5 FILLER_158_328 ();
 b15zdnd11an1n32x5 FILLER_158_392 ();
 b15zdnd11an1n16x5 FILLER_158_424 ();
 b15zdnd11an1n04x5 FILLER_158_440 ();
 b15zdnd00an1n02x5 FILLER_158_444 ();
 b15zdnd11an1n64x5 FILLER_158_468 ();
 b15zdnd11an1n64x5 FILLER_158_532 ();
 b15zdnd11an1n64x5 FILLER_158_596 ();
 b15zdnd11an1n32x5 FILLER_158_660 ();
 b15zdnd11an1n16x5 FILLER_158_692 ();
 b15zdnd11an1n08x5 FILLER_158_708 ();
 b15zdnd00an1n02x5 FILLER_158_716 ();
 b15zdnd11an1n64x5 FILLER_158_726 ();
 b15zdnd11an1n64x5 FILLER_158_790 ();
 b15zdnd11an1n64x5 FILLER_158_854 ();
 b15zdnd11an1n64x5 FILLER_158_918 ();
 b15zdnd11an1n64x5 FILLER_158_982 ();
 b15zdnd11an1n64x5 FILLER_158_1046 ();
 b15zdnd11an1n64x5 FILLER_158_1110 ();
 b15zdnd11an1n64x5 FILLER_158_1174 ();
 b15zdnd11an1n16x5 FILLER_158_1238 ();
 b15zdnd11an1n08x5 FILLER_158_1254 ();
 b15zdnd00an1n01x5 FILLER_158_1262 ();
 b15zdnd11an1n04x5 FILLER_158_1315 ();
 b15zdnd11an1n64x5 FILLER_158_1361 ();
 b15zdnd11an1n32x5 FILLER_158_1425 ();
 b15zdnd11an1n16x5 FILLER_158_1457 ();
 b15zdnd11an1n04x5 FILLER_158_1473 ();
 b15zdnd00an1n01x5 FILLER_158_1477 ();
 b15zdnd00an1n02x5 FILLER_158_2265 ();
 b15zdnd00an1n01x5 FILLER_158_2267 ();
 b15zdnd00an1n02x5 FILLER_158_2274 ();
 b15zdnd11an1n64x5 FILLER_159_0 ();
 b15zdnd11an1n64x5 FILLER_159_64 ();
 b15zdnd11an1n64x5 FILLER_159_128 ();
 b15zdnd11an1n64x5 FILLER_159_192 ();
 b15zdnd11an1n64x5 FILLER_159_256 ();
 b15zdnd11an1n64x5 FILLER_159_320 ();
 b15zdnd11an1n64x5 FILLER_159_384 ();
 b15zdnd11an1n64x5 FILLER_159_448 ();
 b15zdnd11an1n64x5 FILLER_159_512 ();
 b15zdnd11an1n64x5 FILLER_159_576 ();
 b15zdnd11an1n64x5 FILLER_159_640 ();
 b15zdnd11an1n64x5 FILLER_159_704 ();
 b15zdnd11an1n64x5 FILLER_159_768 ();
 b15zdnd11an1n64x5 FILLER_159_832 ();
 b15zdnd11an1n64x5 FILLER_159_896 ();
 b15zdnd11an1n64x5 FILLER_159_969 ();
 b15zdnd11an1n64x5 FILLER_159_1033 ();
 b15zdnd11an1n16x5 FILLER_159_1097 ();
 b15zdnd11an1n04x5 FILLER_159_1113 ();
 b15zdnd00an1n02x5 FILLER_159_1117 ();
 b15zdnd00an1n01x5 FILLER_159_1119 ();
 b15zdnd11an1n04x5 FILLER_159_1128 ();
 b15zdnd11an1n64x5 FILLER_159_1140 ();
 b15zdnd11an1n64x5 FILLER_159_1204 ();
 b15zdnd11an1n08x5 FILLER_159_1268 ();
 b15zdnd11an1n04x5 FILLER_159_1276 ();
 b15zdnd00an1n01x5 FILLER_159_1280 ();
 b15zdnd11an1n04x5 FILLER_159_1284 ();
 b15zdnd00an1n02x5 FILLER_159_1288 ();
 b15zdnd11an1n64x5 FILLER_159_1332 ();
 b15zdnd11an1n64x5 FILLER_159_1396 ();
 b15zdnd11an1n16x5 FILLER_159_1460 ();
 b15zdnd11an1n08x5 FILLER_159_1476 ();
 b15zdnd00an1n02x5 FILLER_159_1484 ();
 b15zdnd11an1n16x5 FILLER_159_2257 ();
 b15zdnd11an1n08x5 FILLER_159_2273 ();
 b15zdnd00an1n02x5 FILLER_159_2281 ();
 b15zdnd00an1n01x5 FILLER_159_2283 ();
 b15zdnd11an1n64x5 FILLER_160_8 ();
 b15zdnd11an1n64x5 FILLER_160_72 ();
 b15zdnd11an1n64x5 FILLER_160_136 ();
 b15zdnd11an1n64x5 FILLER_160_200 ();
 b15zdnd11an1n64x5 FILLER_160_264 ();
 b15zdnd11an1n64x5 FILLER_160_328 ();
 b15zdnd11an1n32x5 FILLER_160_392 ();
 b15zdnd11an1n08x5 FILLER_160_424 ();
 b15zdnd11an1n04x5 FILLER_160_432 ();
 b15zdnd00an1n02x5 FILLER_160_436 ();
 b15zdnd00an1n01x5 FILLER_160_438 ();
 b15zdnd11an1n64x5 FILLER_160_453 ();
 b15zdnd11an1n64x5 FILLER_160_517 ();
 b15zdnd11an1n64x5 FILLER_160_581 ();
 b15zdnd11an1n64x5 FILLER_160_645 ();
 b15zdnd11an1n08x5 FILLER_160_709 ();
 b15zdnd00an1n01x5 FILLER_160_717 ();
 b15zdnd11an1n64x5 FILLER_160_726 ();
 b15zdnd11an1n64x5 FILLER_160_790 ();
 b15zdnd11an1n64x5 FILLER_160_854 ();
 b15zdnd11an1n64x5 FILLER_160_918 ();
 b15zdnd11an1n64x5 FILLER_160_982 ();
 b15zdnd11an1n64x5 FILLER_160_1046 ();
 b15zdnd11an1n64x5 FILLER_160_1110 ();
 b15zdnd11an1n64x5 FILLER_160_1174 ();
 b15zdnd11an1n32x5 FILLER_160_1238 ();
 b15zdnd11an1n16x5 FILLER_160_1270 ();
 b15zdnd00an1n02x5 FILLER_160_1286 ();
 b15zdnd11an1n64x5 FILLER_160_1291 ();
 b15zdnd11an1n64x5 FILLER_160_1355 ();
 b15zdnd11an1n32x5 FILLER_160_1419 ();
 b15zdnd11an1n16x5 FILLER_160_1451 ();
 b15zdnd11an1n08x5 FILLER_160_1467 ();
 b15zdnd00an1n02x5 FILLER_160_1475 ();
 b15zdnd00an1n01x5 FILLER_160_1477 ();
 b15zdnd11an1n08x5 FILLER_160_2265 ();
 b15zdnd00an1n02x5 FILLER_160_2273 ();
 b15zdnd00an1n01x5 FILLER_160_2275 ();
 b15zdnd11an1n64x5 FILLER_161_0 ();
 b15zdnd11an1n64x5 FILLER_161_64 ();
 b15zdnd11an1n64x5 FILLER_161_128 ();
 b15zdnd11an1n64x5 FILLER_161_192 ();
 b15zdnd11an1n64x5 FILLER_161_256 ();
 b15zdnd11an1n64x5 FILLER_161_320 ();
 b15zdnd11an1n32x5 FILLER_161_384 ();
 b15zdnd11an1n08x5 FILLER_161_416 ();
 b15zdnd00an1n02x5 FILLER_161_424 ();
 b15zdnd00an1n01x5 FILLER_161_426 ();
 b15zdnd11an1n64x5 FILLER_161_442 ();
 b15zdnd11an1n64x5 FILLER_161_506 ();
 b15zdnd11an1n64x5 FILLER_161_570 ();
 b15zdnd11an1n64x5 FILLER_161_634 ();
 b15zdnd11an1n64x5 FILLER_161_698 ();
 b15zdnd11an1n64x5 FILLER_161_762 ();
 b15zdnd11an1n64x5 FILLER_161_826 ();
 b15zdnd11an1n64x5 FILLER_161_890 ();
 b15zdnd11an1n64x5 FILLER_161_954 ();
 b15zdnd11an1n64x5 FILLER_161_1018 ();
 b15zdnd11an1n64x5 FILLER_161_1082 ();
 b15zdnd11an1n64x5 FILLER_161_1146 ();
 b15zdnd11an1n64x5 FILLER_161_1210 ();
 b15zdnd11an1n64x5 FILLER_161_1274 ();
 b15zdnd11an1n64x5 FILLER_161_1338 ();
 b15zdnd11an1n64x5 FILLER_161_1402 ();
 b15zdnd11an1n16x5 FILLER_161_1466 ();
 b15zdnd11an1n04x5 FILLER_161_1482 ();
 b15zdnd11an1n16x5 FILLER_161_2257 ();
 b15zdnd11an1n08x5 FILLER_161_2273 ();
 b15zdnd00an1n02x5 FILLER_161_2281 ();
 b15zdnd00an1n01x5 FILLER_161_2283 ();
 b15zdnd11an1n64x5 FILLER_162_8 ();
 b15zdnd11an1n64x5 FILLER_162_72 ();
 b15zdnd11an1n64x5 FILLER_162_136 ();
 b15zdnd11an1n64x5 FILLER_162_200 ();
 b15zdnd11an1n64x5 FILLER_162_264 ();
 b15zdnd11an1n64x5 FILLER_162_328 ();
 b15zdnd11an1n64x5 FILLER_162_392 ();
 b15zdnd11an1n64x5 FILLER_162_456 ();
 b15zdnd11an1n64x5 FILLER_162_520 ();
 b15zdnd11an1n64x5 FILLER_162_584 ();
 b15zdnd11an1n64x5 FILLER_162_648 ();
 b15zdnd11an1n04x5 FILLER_162_712 ();
 b15zdnd00an1n02x5 FILLER_162_716 ();
 b15zdnd11an1n64x5 FILLER_162_726 ();
 b15zdnd11an1n64x5 FILLER_162_790 ();
 b15zdnd11an1n64x5 FILLER_162_854 ();
 b15zdnd11an1n64x5 FILLER_162_918 ();
 b15zdnd11an1n64x5 FILLER_162_982 ();
 b15zdnd11an1n16x5 FILLER_162_1046 ();
 b15zdnd00an1n02x5 FILLER_162_1062 ();
 b15zdnd11an1n64x5 FILLER_162_1072 ();
 b15zdnd11an1n64x5 FILLER_162_1136 ();
 b15zdnd11an1n64x5 FILLER_162_1200 ();
 b15zdnd11an1n64x5 FILLER_162_1264 ();
 b15zdnd11an1n64x5 FILLER_162_1328 ();
 b15zdnd11an1n64x5 FILLER_162_1392 ();
 b15zdnd11an1n16x5 FILLER_162_1456 ();
 b15zdnd11an1n04x5 FILLER_162_1472 ();
 b15zdnd00an1n02x5 FILLER_162_1476 ();
 b15zdnd11an1n08x5 FILLER_162_2265 ();
 b15zdnd00an1n02x5 FILLER_162_2273 ();
 b15zdnd00an1n01x5 FILLER_162_2275 ();
 b15zdnd11an1n08x5 FILLER_163_0 ();
 b15zdnd11an1n04x5 FILLER_163_8 ();
 b15zdnd00an1n02x5 FILLER_163_12 ();
 b15zdnd11an1n64x5 FILLER_163_25 ();
 b15zdnd11an1n64x5 FILLER_163_89 ();
 b15zdnd11an1n64x5 FILLER_163_153 ();
 b15zdnd11an1n64x5 FILLER_163_217 ();
 b15zdnd11an1n64x5 FILLER_163_281 ();
 b15zdnd11an1n64x5 FILLER_163_345 ();
 b15zdnd11an1n64x5 FILLER_163_409 ();
 b15zdnd11an1n64x5 FILLER_163_473 ();
 b15zdnd11an1n64x5 FILLER_163_537 ();
 b15zdnd11an1n64x5 FILLER_163_601 ();
 b15zdnd11an1n64x5 FILLER_163_665 ();
 b15zdnd11an1n64x5 FILLER_163_729 ();
 b15zdnd11an1n64x5 FILLER_163_793 ();
 b15zdnd11an1n64x5 FILLER_163_857 ();
 b15zdnd11an1n64x5 FILLER_163_921 ();
 b15zdnd11an1n64x5 FILLER_163_985 ();
 b15zdnd11an1n64x5 FILLER_163_1049 ();
 b15zdnd11an1n64x5 FILLER_163_1113 ();
 b15zdnd11an1n64x5 FILLER_163_1177 ();
 b15zdnd11an1n64x5 FILLER_163_1241 ();
 b15zdnd11an1n64x5 FILLER_163_1305 ();
 b15zdnd11an1n64x5 FILLER_163_1369 ();
 b15zdnd11an1n32x5 FILLER_163_1433 ();
 b15zdnd11an1n16x5 FILLER_163_1465 ();
 b15zdnd11an1n04x5 FILLER_163_1481 ();
 b15zdnd00an1n01x5 FILLER_163_1485 ();
 b15zdnd00an1n02x5 FILLER_163_2257 ();
 b15zdnd11an1n16x5 FILLER_163_2265 ();
 b15zdnd00an1n02x5 FILLER_163_2281 ();
 b15zdnd00an1n01x5 FILLER_163_2283 ();
 b15zdnd11an1n64x5 FILLER_164_8 ();
 b15zdnd11an1n64x5 FILLER_164_72 ();
 b15zdnd11an1n64x5 FILLER_164_136 ();
 b15zdnd11an1n64x5 FILLER_164_200 ();
 b15zdnd11an1n64x5 FILLER_164_264 ();
 b15zdnd11an1n64x5 FILLER_164_328 ();
 b15zdnd11an1n32x5 FILLER_164_392 ();
 b15zdnd11an1n16x5 FILLER_164_424 ();
 b15zdnd00an1n02x5 FILLER_164_440 ();
 b15zdnd11an1n64x5 FILLER_164_484 ();
 b15zdnd11an1n64x5 FILLER_164_548 ();
 b15zdnd11an1n64x5 FILLER_164_612 ();
 b15zdnd11an1n32x5 FILLER_164_676 ();
 b15zdnd11an1n08x5 FILLER_164_708 ();
 b15zdnd00an1n02x5 FILLER_164_716 ();
 b15zdnd11an1n64x5 FILLER_164_726 ();
 b15zdnd11an1n64x5 FILLER_164_790 ();
 b15zdnd11an1n64x5 FILLER_164_854 ();
 b15zdnd11an1n64x5 FILLER_164_918 ();
 b15zdnd11an1n64x5 FILLER_164_982 ();
 b15zdnd11an1n64x5 FILLER_164_1046 ();
 b15zdnd11an1n64x5 FILLER_164_1110 ();
 b15zdnd11an1n64x5 FILLER_164_1174 ();
 b15zdnd11an1n64x5 FILLER_164_1238 ();
 b15zdnd11an1n64x5 FILLER_164_1302 ();
 b15zdnd11an1n64x5 FILLER_164_1366 ();
 b15zdnd11an1n32x5 FILLER_164_1430 ();
 b15zdnd11an1n16x5 FILLER_164_1462 ();
 b15zdnd00an1n02x5 FILLER_164_2265 ();
 b15zdnd00an1n01x5 FILLER_164_2267 ();
 b15zdnd00an1n02x5 FILLER_164_2274 ();
 b15zdnd11an1n64x5 FILLER_165_0 ();
 b15zdnd11an1n64x5 FILLER_165_64 ();
 b15zdnd11an1n64x5 FILLER_165_128 ();
 b15zdnd11an1n64x5 FILLER_165_192 ();
 b15zdnd11an1n64x5 FILLER_165_256 ();
 b15zdnd11an1n64x5 FILLER_165_320 ();
 b15zdnd11an1n64x5 FILLER_165_384 ();
 b15zdnd11an1n64x5 FILLER_165_448 ();
 b15zdnd11an1n64x5 FILLER_165_512 ();
 b15zdnd11an1n64x5 FILLER_165_576 ();
 b15zdnd11an1n64x5 FILLER_165_640 ();
 b15zdnd11an1n64x5 FILLER_165_704 ();
 b15zdnd11an1n64x5 FILLER_165_768 ();
 b15zdnd11an1n64x5 FILLER_165_832 ();
 b15zdnd11an1n64x5 FILLER_165_896 ();
 b15zdnd11an1n64x5 FILLER_165_960 ();
 b15zdnd11an1n64x5 FILLER_165_1024 ();
 b15zdnd11an1n32x5 FILLER_165_1088 ();
 b15zdnd11an1n08x5 FILLER_165_1120 ();
 b15zdnd11an1n04x5 FILLER_165_1128 ();
 b15zdnd00an1n01x5 FILLER_165_1132 ();
 b15zdnd11an1n64x5 FILLER_165_1175 ();
 b15zdnd11an1n64x5 FILLER_165_1239 ();
 b15zdnd11an1n64x5 FILLER_165_1303 ();
 b15zdnd11an1n64x5 FILLER_165_1367 ();
 b15zdnd11an1n32x5 FILLER_165_1431 ();
 b15zdnd11an1n16x5 FILLER_165_1463 ();
 b15zdnd11an1n04x5 FILLER_165_1479 ();
 b15zdnd00an1n02x5 FILLER_165_1483 ();
 b15zdnd00an1n01x5 FILLER_165_1485 ();
 b15zdnd11an1n16x5 FILLER_165_2257 ();
 b15zdnd11an1n08x5 FILLER_165_2273 ();
 b15zdnd00an1n02x5 FILLER_165_2281 ();
 b15zdnd00an1n01x5 FILLER_165_2283 ();
 b15zdnd11an1n64x5 FILLER_166_8 ();
 b15zdnd11an1n64x5 FILLER_166_72 ();
 b15zdnd11an1n64x5 FILLER_166_136 ();
 b15zdnd11an1n64x5 FILLER_166_200 ();
 b15zdnd11an1n64x5 FILLER_166_264 ();
 b15zdnd11an1n64x5 FILLER_166_328 ();
 b15zdnd11an1n32x5 FILLER_166_392 ();
 b15zdnd11an1n08x5 FILLER_166_424 ();
 b15zdnd11an1n04x5 FILLER_166_432 ();
 b15zdnd00an1n02x5 FILLER_166_436 ();
 b15zdnd00an1n01x5 FILLER_166_438 ();
 b15zdnd11an1n64x5 FILLER_166_451 ();
 b15zdnd11an1n64x5 FILLER_166_515 ();
 b15zdnd11an1n64x5 FILLER_166_579 ();
 b15zdnd11an1n64x5 FILLER_166_643 ();
 b15zdnd11an1n08x5 FILLER_166_707 ();
 b15zdnd00an1n02x5 FILLER_166_715 ();
 b15zdnd00an1n01x5 FILLER_166_717 ();
 b15zdnd11an1n64x5 FILLER_166_726 ();
 b15zdnd11an1n64x5 FILLER_166_790 ();
 b15zdnd11an1n64x5 FILLER_166_854 ();
 b15zdnd11an1n64x5 FILLER_166_918 ();
 b15zdnd11an1n64x5 FILLER_166_982 ();
 b15zdnd11an1n64x5 FILLER_166_1046 ();
 b15zdnd11an1n64x5 FILLER_166_1110 ();
 b15zdnd00an1n02x5 FILLER_166_1174 ();
 b15zdnd00an1n01x5 FILLER_166_1176 ();
 b15zdnd11an1n64x5 FILLER_166_1219 ();
 b15zdnd11an1n64x5 FILLER_166_1283 ();
 b15zdnd11an1n64x5 FILLER_166_1347 ();
 b15zdnd11an1n64x5 FILLER_166_1411 ();
 b15zdnd00an1n02x5 FILLER_166_1475 ();
 b15zdnd00an1n01x5 FILLER_166_1477 ();
 b15zdnd11an1n08x5 FILLER_166_2265 ();
 b15zdnd00an1n02x5 FILLER_166_2273 ();
 b15zdnd00an1n01x5 FILLER_166_2275 ();
 b15zdnd11an1n64x5 FILLER_167_0 ();
 b15zdnd11an1n64x5 FILLER_167_64 ();
 b15zdnd11an1n64x5 FILLER_167_128 ();
 b15zdnd11an1n64x5 FILLER_167_192 ();
 b15zdnd11an1n64x5 FILLER_167_256 ();
 b15zdnd11an1n64x5 FILLER_167_320 ();
 b15zdnd11an1n64x5 FILLER_167_384 ();
 b15zdnd11an1n64x5 FILLER_167_448 ();
 b15zdnd11an1n64x5 FILLER_167_512 ();
 b15zdnd11an1n64x5 FILLER_167_576 ();
 b15zdnd11an1n64x5 FILLER_167_640 ();
 b15zdnd11an1n64x5 FILLER_167_704 ();
 b15zdnd11an1n64x5 FILLER_167_768 ();
 b15zdnd11an1n64x5 FILLER_167_832 ();
 b15zdnd11an1n64x5 FILLER_167_896 ();
 b15zdnd11an1n64x5 FILLER_167_960 ();
 b15zdnd11an1n64x5 FILLER_167_1024 ();
 b15zdnd11an1n64x5 FILLER_167_1088 ();
 b15zdnd11an1n64x5 FILLER_167_1152 ();
 b15zdnd11an1n64x5 FILLER_167_1216 ();
 b15zdnd11an1n64x5 FILLER_167_1280 ();
 b15zdnd11an1n64x5 FILLER_167_1344 ();
 b15zdnd11an1n64x5 FILLER_167_1408 ();
 b15zdnd11an1n08x5 FILLER_167_1472 ();
 b15zdnd11an1n04x5 FILLER_167_1480 ();
 b15zdnd00an1n02x5 FILLER_167_1484 ();
 b15zdnd11an1n16x5 FILLER_167_2257 ();
 b15zdnd11an1n08x5 FILLER_167_2273 ();
 b15zdnd00an1n02x5 FILLER_167_2281 ();
 b15zdnd00an1n01x5 FILLER_167_2283 ();
 b15zdnd11an1n64x5 FILLER_168_8 ();
 b15zdnd11an1n64x5 FILLER_168_72 ();
 b15zdnd11an1n64x5 FILLER_168_136 ();
 b15zdnd11an1n32x5 FILLER_168_200 ();
 b15zdnd11an1n04x5 FILLER_168_232 ();
 b15zdnd11an1n64x5 FILLER_168_278 ();
 b15zdnd11an1n64x5 FILLER_168_342 ();
 b15zdnd11an1n32x5 FILLER_168_406 ();
 b15zdnd11an1n08x5 FILLER_168_438 ();
 b15zdnd11an1n04x5 FILLER_168_446 ();
 b15zdnd00an1n02x5 FILLER_168_450 ();
 b15zdnd11an1n64x5 FILLER_168_464 ();
 b15zdnd11an1n64x5 FILLER_168_528 ();
 b15zdnd11an1n64x5 FILLER_168_592 ();
 b15zdnd11an1n32x5 FILLER_168_656 ();
 b15zdnd11an1n16x5 FILLER_168_688 ();
 b15zdnd11an1n08x5 FILLER_168_704 ();
 b15zdnd11an1n04x5 FILLER_168_712 ();
 b15zdnd00an1n02x5 FILLER_168_716 ();
 b15zdnd11an1n64x5 FILLER_168_726 ();
 b15zdnd11an1n64x5 FILLER_168_790 ();
 b15zdnd11an1n64x5 FILLER_168_854 ();
 b15zdnd11an1n64x5 FILLER_168_918 ();
 b15zdnd11an1n32x5 FILLER_168_982 ();
 b15zdnd11an1n16x5 FILLER_168_1014 ();
 b15zdnd11an1n08x5 FILLER_168_1030 ();
 b15zdnd00an1n02x5 FILLER_168_1038 ();
 b15zdnd11an1n64x5 FILLER_168_1050 ();
 b15zdnd11an1n64x5 FILLER_168_1114 ();
 b15zdnd11an1n64x5 FILLER_168_1178 ();
 b15zdnd11an1n64x5 FILLER_168_1242 ();
 b15zdnd11an1n64x5 FILLER_168_1306 ();
 b15zdnd11an1n64x5 FILLER_168_1370 ();
 b15zdnd11an1n16x5 FILLER_168_1434 ();
 b15zdnd11an1n08x5 FILLER_168_1450 ();
 b15zdnd00an1n02x5 FILLER_168_1458 ();
 b15zdnd11an1n08x5 FILLER_168_1469 ();
 b15zdnd00an1n01x5 FILLER_168_1477 ();
 b15zdnd11an1n08x5 FILLER_168_2265 ();
 b15zdnd00an1n02x5 FILLER_168_2273 ();
 b15zdnd00an1n01x5 FILLER_168_2275 ();
 b15zdnd11an1n64x5 FILLER_169_0 ();
 b15zdnd11an1n64x5 FILLER_169_64 ();
 b15zdnd11an1n64x5 FILLER_169_128 ();
 b15zdnd11an1n64x5 FILLER_169_192 ();
 b15zdnd11an1n64x5 FILLER_169_256 ();
 b15zdnd11an1n64x5 FILLER_169_320 ();
 b15zdnd11an1n32x5 FILLER_169_384 ();
 b15zdnd11an1n16x5 FILLER_169_416 ();
 b15zdnd11an1n08x5 FILLER_169_432 ();
 b15zdnd11an1n64x5 FILLER_169_482 ();
 b15zdnd11an1n64x5 FILLER_169_546 ();
 b15zdnd11an1n64x5 FILLER_169_610 ();
 b15zdnd11an1n64x5 FILLER_169_674 ();
 b15zdnd11an1n64x5 FILLER_169_738 ();
 b15zdnd11an1n64x5 FILLER_169_802 ();
 b15zdnd11an1n64x5 FILLER_169_866 ();
 b15zdnd11an1n64x5 FILLER_169_930 ();
 b15zdnd11an1n64x5 FILLER_169_994 ();
 b15zdnd11an1n64x5 FILLER_169_1058 ();
 b15zdnd11an1n64x5 FILLER_169_1122 ();
 b15zdnd11an1n64x5 FILLER_169_1186 ();
 b15zdnd11an1n64x5 FILLER_169_1250 ();
 b15zdnd11an1n64x5 FILLER_169_1314 ();
 b15zdnd11an1n64x5 FILLER_169_1378 ();
 b15zdnd11an1n32x5 FILLER_169_1442 ();
 b15zdnd11an1n08x5 FILLER_169_1474 ();
 b15zdnd11an1n04x5 FILLER_169_1482 ();
 b15zdnd11an1n16x5 FILLER_169_2257 ();
 b15zdnd11an1n08x5 FILLER_169_2273 ();
 b15zdnd00an1n02x5 FILLER_169_2281 ();
 b15zdnd00an1n01x5 FILLER_169_2283 ();
 b15zdnd11an1n16x5 FILLER_170_8 ();
 b15zdnd11an1n64x5 FILLER_170_28 ();
 b15zdnd11an1n64x5 FILLER_170_92 ();
 b15zdnd11an1n64x5 FILLER_170_156 ();
 b15zdnd11an1n64x5 FILLER_170_220 ();
 b15zdnd11an1n64x5 FILLER_170_284 ();
 b15zdnd11an1n64x5 FILLER_170_348 ();
 b15zdnd11an1n32x5 FILLER_170_412 ();
 b15zdnd11an1n16x5 FILLER_170_444 ();
 b15zdnd11an1n04x5 FILLER_170_460 ();
 b15zdnd00an1n02x5 FILLER_170_464 ();
 b15zdnd00an1n01x5 FILLER_170_466 ();
 b15zdnd11an1n64x5 FILLER_170_483 ();
 b15zdnd11an1n64x5 FILLER_170_547 ();
 b15zdnd11an1n64x5 FILLER_170_611 ();
 b15zdnd11an1n32x5 FILLER_170_675 ();
 b15zdnd11an1n08x5 FILLER_170_707 ();
 b15zdnd00an1n02x5 FILLER_170_715 ();
 b15zdnd00an1n01x5 FILLER_170_717 ();
 b15zdnd11an1n64x5 FILLER_170_726 ();
 b15zdnd11an1n64x5 FILLER_170_790 ();
 b15zdnd11an1n64x5 FILLER_170_854 ();
 b15zdnd11an1n64x5 FILLER_170_918 ();
 b15zdnd11an1n64x5 FILLER_170_982 ();
 b15zdnd11an1n64x5 FILLER_170_1046 ();
 b15zdnd11an1n64x5 FILLER_170_1110 ();
 b15zdnd11an1n64x5 FILLER_170_1174 ();
 b15zdnd11an1n64x5 FILLER_170_1238 ();
 b15zdnd11an1n64x5 FILLER_170_1302 ();
 b15zdnd11an1n64x5 FILLER_170_1366 ();
 b15zdnd11an1n32x5 FILLER_170_1430 ();
 b15zdnd11an1n16x5 FILLER_170_1462 ();
 b15zdnd11an1n08x5 FILLER_170_2265 ();
 b15zdnd00an1n02x5 FILLER_170_2273 ();
 b15zdnd00an1n01x5 FILLER_170_2275 ();
 b15zdnd11an1n08x5 FILLER_171_0 ();
 b15zdnd11an1n64x5 FILLER_171_50 ();
 b15zdnd11an1n64x5 FILLER_171_114 ();
 b15zdnd11an1n64x5 FILLER_171_178 ();
 b15zdnd11an1n64x5 FILLER_171_242 ();
 b15zdnd11an1n64x5 FILLER_171_306 ();
 b15zdnd11an1n64x5 FILLER_171_370 ();
 b15zdnd11an1n08x5 FILLER_171_434 ();
 b15zdnd11an1n04x5 FILLER_171_442 ();
 b15zdnd00an1n02x5 FILLER_171_446 ();
 b15zdnd00an1n01x5 FILLER_171_448 ();
 b15zdnd11an1n64x5 FILLER_171_491 ();
 b15zdnd11an1n64x5 FILLER_171_555 ();
 b15zdnd11an1n64x5 FILLER_171_619 ();
 b15zdnd11an1n64x5 FILLER_171_683 ();
 b15zdnd11an1n64x5 FILLER_171_747 ();
 b15zdnd11an1n64x5 FILLER_171_811 ();
 b15zdnd11an1n64x5 FILLER_171_875 ();
 b15zdnd11an1n64x5 FILLER_171_939 ();
 b15zdnd11an1n64x5 FILLER_171_1003 ();
 b15zdnd11an1n64x5 FILLER_171_1067 ();
 b15zdnd11an1n64x5 FILLER_171_1131 ();
 b15zdnd11an1n64x5 FILLER_171_1195 ();
 b15zdnd11an1n64x5 FILLER_171_1259 ();
 b15zdnd11an1n64x5 FILLER_171_1323 ();
 b15zdnd11an1n64x5 FILLER_171_1387 ();
 b15zdnd11an1n32x5 FILLER_171_1451 ();
 b15zdnd00an1n02x5 FILLER_171_1483 ();
 b15zdnd00an1n01x5 FILLER_171_1485 ();
 b15zdnd11an1n16x5 FILLER_171_2257 ();
 b15zdnd11an1n08x5 FILLER_171_2273 ();
 b15zdnd00an1n02x5 FILLER_171_2281 ();
 b15zdnd00an1n01x5 FILLER_171_2283 ();
 b15zdnd11an1n64x5 FILLER_172_8 ();
 b15zdnd11an1n64x5 FILLER_172_72 ();
 b15zdnd11an1n64x5 FILLER_172_136 ();
 b15zdnd11an1n64x5 FILLER_172_200 ();
 b15zdnd11an1n64x5 FILLER_172_264 ();
 b15zdnd11an1n64x5 FILLER_172_328 ();
 b15zdnd11an1n64x5 FILLER_172_392 ();
 b15zdnd11an1n64x5 FILLER_172_456 ();
 b15zdnd11an1n64x5 FILLER_172_520 ();
 b15zdnd11an1n64x5 FILLER_172_584 ();
 b15zdnd11an1n64x5 FILLER_172_648 ();
 b15zdnd11an1n04x5 FILLER_172_712 ();
 b15zdnd00an1n02x5 FILLER_172_716 ();
 b15zdnd11an1n64x5 FILLER_172_726 ();
 b15zdnd11an1n64x5 FILLER_172_790 ();
 b15zdnd11an1n64x5 FILLER_172_854 ();
 b15zdnd11an1n64x5 FILLER_172_918 ();
 b15zdnd11an1n04x5 FILLER_172_982 ();
 b15zdnd00an1n02x5 FILLER_172_986 ();
 b15zdnd11an1n16x5 FILLER_172_997 ();
 b15zdnd00an1n02x5 FILLER_172_1013 ();
 b15zdnd00an1n01x5 FILLER_172_1015 ();
 b15zdnd11an1n04x5 FILLER_172_1025 ();
 b15zdnd11an1n32x5 FILLER_172_1032 ();
 b15zdnd11an1n16x5 FILLER_172_1064 ();
 b15zdnd11an1n04x5 FILLER_172_1080 ();
 b15zdnd00an1n02x5 FILLER_172_1084 ();
 b15zdnd00an1n01x5 FILLER_172_1086 ();
 b15zdnd11an1n64x5 FILLER_172_1095 ();
 b15zdnd11an1n64x5 FILLER_172_1159 ();
 b15zdnd11an1n64x5 FILLER_172_1223 ();
 b15zdnd11an1n64x5 FILLER_172_1287 ();
 b15zdnd11an1n64x5 FILLER_172_1351 ();
 b15zdnd11an1n32x5 FILLER_172_1415 ();
 b15zdnd11an1n16x5 FILLER_172_1447 ();
 b15zdnd11an1n08x5 FILLER_172_1463 ();
 b15zdnd11an1n04x5 FILLER_172_1471 ();
 b15zdnd00an1n02x5 FILLER_172_1475 ();
 b15zdnd00an1n01x5 FILLER_172_1477 ();
 b15zdnd11an1n08x5 FILLER_172_2265 ();
 b15zdnd00an1n02x5 FILLER_172_2273 ();
 b15zdnd00an1n01x5 FILLER_172_2275 ();
 b15zdnd11an1n64x5 FILLER_173_0 ();
 b15zdnd11an1n64x5 FILLER_173_64 ();
 b15zdnd11an1n64x5 FILLER_173_128 ();
 b15zdnd11an1n64x5 FILLER_173_192 ();
 b15zdnd11an1n64x5 FILLER_173_256 ();
 b15zdnd11an1n64x5 FILLER_173_320 ();
 b15zdnd11an1n04x5 FILLER_173_384 ();
 b15zdnd00an1n02x5 FILLER_173_388 ();
 b15zdnd00an1n01x5 FILLER_173_390 ();
 b15zdnd11an1n32x5 FILLER_173_403 ();
 b15zdnd11an1n16x5 FILLER_173_435 ();
 b15zdnd11an1n04x5 FILLER_173_451 ();
 b15zdnd00an1n02x5 FILLER_173_455 ();
 b15zdnd00an1n01x5 FILLER_173_457 ();
 b15zdnd11an1n64x5 FILLER_173_476 ();
 b15zdnd11an1n64x5 FILLER_173_540 ();
 b15zdnd11an1n64x5 FILLER_173_604 ();
 b15zdnd11an1n64x5 FILLER_173_668 ();
 b15zdnd11an1n64x5 FILLER_173_732 ();
 b15zdnd11an1n64x5 FILLER_173_796 ();
 b15zdnd11an1n64x5 FILLER_173_860 ();
 b15zdnd11an1n64x5 FILLER_173_924 ();
 b15zdnd11an1n64x5 FILLER_173_1032 ();
 b15zdnd11an1n64x5 FILLER_173_1096 ();
 b15zdnd11an1n64x5 FILLER_173_1160 ();
 b15zdnd11an1n64x5 FILLER_173_1224 ();
 b15zdnd11an1n64x5 FILLER_173_1288 ();
 b15zdnd11an1n64x5 FILLER_173_1352 ();
 b15zdnd11an1n64x5 FILLER_173_1416 ();
 b15zdnd11an1n04x5 FILLER_173_1480 ();
 b15zdnd00an1n02x5 FILLER_173_1484 ();
 b15zdnd11an1n16x5 FILLER_173_2257 ();
 b15zdnd11an1n08x5 FILLER_173_2273 ();
 b15zdnd00an1n02x5 FILLER_173_2281 ();
 b15zdnd00an1n01x5 FILLER_173_2283 ();
 b15zdnd11an1n64x5 FILLER_174_8 ();
 b15zdnd11an1n64x5 FILLER_174_72 ();
 b15zdnd11an1n64x5 FILLER_174_136 ();
 b15zdnd11an1n64x5 FILLER_174_200 ();
 b15zdnd11an1n64x5 FILLER_174_264 ();
 b15zdnd11an1n64x5 FILLER_174_328 ();
 b15zdnd11an1n64x5 FILLER_174_392 ();
 b15zdnd11an1n08x5 FILLER_174_456 ();
 b15zdnd11an1n04x5 FILLER_174_464 ();
 b15zdnd00an1n02x5 FILLER_174_468 ();
 b15zdnd11an1n64x5 FILLER_174_482 ();
 b15zdnd11an1n64x5 FILLER_174_546 ();
 b15zdnd11an1n64x5 FILLER_174_610 ();
 b15zdnd11an1n32x5 FILLER_174_674 ();
 b15zdnd11an1n08x5 FILLER_174_706 ();
 b15zdnd11an1n04x5 FILLER_174_714 ();
 b15zdnd11an1n64x5 FILLER_174_726 ();
 b15zdnd11an1n64x5 FILLER_174_790 ();
 b15zdnd11an1n64x5 FILLER_174_854 ();
 b15zdnd11an1n64x5 FILLER_174_918 ();
 b15zdnd11an1n16x5 FILLER_174_982 ();
 b15zdnd11an1n08x5 FILLER_174_998 ();
 b15zdnd00an1n02x5 FILLER_174_1006 ();
 b15zdnd11an1n04x5 FILLER_174_1017 ();
 b15zdnd11an1n08x5 FILLER_174_1024 ();
 b15zdnd11an1n04x5 FILLER_174_1032 ();
 b15zdnd00an1n02x5 FILLER_174_1036 ();
 b15zdnd00an1n01x5 FILLER_174_1038 ();
 b15zdnd11an1n64x5 FILLER_174_1042 ();
 b15zdnd11an1n64x5 FILLER_174_1106 ();
 b15zdnd11an1n64x5 FILLER_174_1170 ();
 b15zdnd11an1n64x5 FILLER_174_1234 ();
 b15zdnd11an1n64x5 FILLER_174_1298 ();
 b15zdnd11an1n64x5 FILLER_174_1362 ();
 b15zdnd11an1n32x5 FILLER_174_1426 ();
 b15zdnd11an1n16x5 FILLER_174_1458 ();
 b15zdnd11an1n04x5 FILLER_174_1474 ();
 b15zdnd11an1n08x5 FILLER_174_2265 ();
 b15zdnd00an1n02x5 FILLER_174_2273 ();
 b15zdnd00an1n01x5 FILLER_174_2275 ();
 b15zdnd11an1n64x5 FILLER_175_0 ();
 b15zdnd11an1n64x5 FILLER_175_64 ();
 b15zdnd11an1n64x5 FILLER_175_128 ();
 b15zdnd11an1n64x5 FILLER_175_192 ();
 b15zdnd11an1n64x5 FILLER_175_256 ();
 b15zdnd11an1n64x5 FILLER_175_320 ();
 b15zdnd11an1n32x5 FILLER_175_384 ();
 b15zdnd11an1n16x5 FILLER_175_416 ();
 b15zdnd11an1n04x5 FILLER_175_432 ();
 b15zdnd00an1n02x5 FILLER_175_436 ();
 b15zdnd11an1n64x5 FILLER_175_442 ();
 b15zdnd11an1n64x5 FILLER_175_506 ();
 b15zdnd11an1n64x5 FILLER_175_570 ();
 b15zdnd11an1n64x5 FILLER_175_634 ();
 b15zdnd11an1n64x5 FILLER_175_698 ();
 b15zdnd11an1n64x5 FILLER_175_762 ();
 b15zdnd11an1n64x5 FILLER_175_826 ();
 b15zdnd11an1n64x5 FILLER_175_890 ();
 b15zdnd11an1n32x5 FILLER_175_954 ();
 b15zdnd11an1n08x5 FILLER_175_986 ();
 b15zdnd11an1n04x5 FILLER_175_1038 ();
 b15zdnd11an1n08x5 FILLER_175_1045 ();
 b15zdnd11an1n64x5 FILLER_175_1056 ();
 b15zdnd11an1n64x5 FILLER_175_1120 ();
 b15zdnd11an1n64x5 FILLER_175_1184 ();
 b15zdnd11an1n64x5 FILLER_175_1248 ();
 b15zdnd11an1n64x5 FILLER_175_1312 ();
 b15zdnd11an1n64x5 FILLER_175_1376 ();
 b15zdnd11an1n32x5 FILLER_175_1440 ();
 b15zdnd11an1n08x5 FILLER_175_1472 ();
 b15zdnd11an1n04x5 FILLER_175_1480 ();
 b15zdnd00an1n02x5 FILLER_175_1484 ();
 b15zdnd11an1n16x5 FILLER_175_2257 ();
 b15zdnd11an1n08x5 FILLER_175_2273 ();
 b15zdnd00an1n02x5 FILLER_175_2281 ();
 b15zdnd00an1n01x5 FILLER_175_2283 ();
 b15zdnd11an1n64x5 FILLER_176_8 ();
 b15zdnd11an1n64x5 FILLER_176_72 ();
 b15zdnd11an1n64x5 FILLER_176_136 ();
 b15zdnd11an1n64x5 FILLER_176_200 ();
 b15zdnd11an1n64x5 FILLER_176_264 ();
 b15zdnd11an1n64x5 FILLER_176_328 ();
 b15zdnd11an1n64x5 FILLER_176_392 ();
 b15zdnd11an1n64x5 FILLER_176_456 ();
 b15zdnd11an1n64x5 FILLER_176_520 ();
 b15zdnd11an1n64x5 FILLER_176_584 ();
 b15zdnd11an1n64x5 FILLER_176_648 ();
 b15zdnd11an1n04x5 FILLER_176_712 ();
 b15zdnd00an1n02x5 FILLER_176_716 ();
 b15zdnd11an1n64x5 FILLER_176_726 ();
 b15zdnd11an1n64x5 FILLER_176_790 ();
 b15zdnd11an1n64x5 FILLER_176_854 ();
 b15zdnd11an1n64x5 FILLER_176_918 ();
 b15zdnd11an1n16x5 FILLER_176_982 ();
 b15zdnd11an1n08x5 FILLER_176_998 ();
 b15zdnd00an1n02x5 FILLER_176_1006 ();
 b15zdnd11an1n04x5 FILLER_176_1011 ();
 b15zdnd11an1n04x5 FILLER_176_1059 ();
 b15zdnd11an1n64x5 FILLER_176_1066 ();
 b15zdnd11an1n64x5 FILLER_176_1130 ();
 b15zdnd11an1n64x5 FILLER_176_1194 ();
 b15zdnd11an1n64x5 FILLER_176_1258 ();
 b15zdnd11an1n64x5 FILLER_176_1322 ();
 b15zdnd11an1n64x5 FILLER_176_1386 ();
 b15zdnd11an1n16x5 FILLER_176_1450 ();
 b15zdnd11an1n08x5 FILLER_176_1466 ();
 b15zdnd11an1n04x5 FILLER_176_1474 ();
 b15zdnd11an1n04x5 FILLER_176_2265 ();
 b15zdnd00an1n02x5 FILLER_176_2273 ();
 b15zdnd00an1n01x5 FILLER_176_2275 ();
 b15zdnd11an1n64x5 FILLER_177_0 ();
 b15zdnd11an1n64x5 FILLER_177_64 ();
 b15zdnd11an1n64x5 FILLER_177_128 ();
 b15zdnd11an1n64x5 FILLER_177_192 ();
 b15zdnd11an1n64x5 FILLER_177_256 ();
 b15zdnd11an1n64x5 FILLER_177_320 ();
 b15zdnd11an1n32x5 FILLER_177_384 ();
 b15zdnd11an1n16x5 FILLER_177_416 ();
 b15zdnd11an1n64x5 FILLER_177_440 ();
 b15zdnd11an1n64x5 FILLER_177_504 ();
 b15zdnd11an1n64x5 FILLER_177_568 ();
 b15zdnd11an1n64x5 FILLER_177_632 ();
 b15zdnd11an1n64x5 FILLER_177_696 ();
 b15zdnd11an1n64x5 FILLER_177_760 ();
 b15zdnd11an1n64x5 FILLER_177_824 ();
 b15zdnd11an1n64x5 FILLER_177_888 ();
 b15zdnd11an1n16x5 FILLER_177_952 ();
 b15zdnd00an1n01x5 FILLER_177_968 ();
 b15zdnd11an1n04x5 FILLER_177_996 ();
 b15zdnd11an1n08x5 FILLER_177_1003 ();
 b15zdnd00an1n02x5 FILLER_177_1011 ();
 b15zdnd00an1n01x5 FILLER_177_1013 ();
 b15zdnd11an1n64x5 FILLER_177_1058 ();
 b15zdnd11an1n64x5 FILLER_177_1122 ();
 b15zdnd11an1n64x5 FILLER_177_1186 ();
 b15zdnd11an1n64x5 FILLER_177_1250 ();
 b15zdnd11an1n64x5 FILLER_177_1314 ();
 b15zdnd11an1n64x5 FILLER_177_1378 ();
 b15zdnd11an1n32x5 FILLER_177_1442 ();
 b15zdnd11an1n08x5 FILLER_177_1474 ();
 b15zdnd11an1n04x5 FILLER_177_1482 ();
 b15zdnd11an1n16x5 FILLER_177_2257 ();
 b15zdnd11an1n08x5 FILLER_177_2273 ();
 b15zdnd00an1n02x5 FILLER_177_2281 ();
 b15zdnd00an1n01x5 FILLER_177_2283 ();
 b15zdnd11an1n64x5 FILLER_178_8 ();
 b15zdnd11an1n64x5 FILLER_178_72 ();
 b15zdnd11an1n64x5 FILLER_178_136 ();
 b15zdnd11an1n64x5 FILLER_178_200 ();
 b15zdnd11an1n64x5 FILLER_178_264 ();
 b15zdnd11an1n64x5 FILLER_178_328 ();
 b15zdnd11an1n64x5 FILLER_178_392 ();
 b15zdnd11an1n64x5 FILLER_178_456 ();
 b15zdnd11an1n64x5 FILLER_178_520 ();
 b15zdnd11an1n64x5 FILLER_178_584 ();
 b15zdnd11an1n64x5 FILLER_178_648 ();
 b15zdnd11an1n04x5 FILLER_178_712 ();
 b15zdnd00an1n02x5 FILLER_178_716 ();
 b15zdnd11an1n64x5 FILLER_178_726 ();
 b15zdnd11an1n64x5 FILLER_178_790 ();
 b15zdnd11an1n64x5 FILLER_178_854 ();
 b15zdnd11an1n64x5 FILLER_178_918 ();
 b15zdnd11an1n32x5 FILLER_178_982 ();
 b15zdnd00an1n01x5 FILLER_178_1014 ();
 b15zdnd11an1n08x5 FILLER_178_1018 ();
 b15zdnd00an1n02x5 FILLER_178_1026 ();
 b15zdnd00an1n01x5 FILLER_178_1028 ();
 b15zdnd11an1n04x5 FILLER_178_1032 ();
 b15zdnd11an1n04x5 FILLER_178_1039 ();
 b15zdnd11an1n08x5 FILLER_178_1046 ();
 b15zdnd00an1n02x5 FILLER_178_1054 ();
 b15zdnd11an1n64x5 FILLER_178_1059 ();
 b15zdnd11an1n64x5 FILLER_178_1123 ();
 b15zdnd11an1n64x5 FILLER_178_1187 ();
 b15zdnd11an1n64x5 FILLER_178_1251 ();
 b15zdnd11an1n64x5 FILLER_178_1315 ();
 b15zdnd11an1n64x5 FILLER_178_1379 ();
 b15zdnd11an1n32x5 FILLER_178_1443 ();
 b15zdnd00an1n02x5 FILLER_178_1475 ();
 b15zdnd00an1n01x5 FILLER_178_1477 ();
 b15zdnd11an1n08x5 FILLER_178_2265 ();
 b15zdnd00an1n02x5 FILLER_178_2273 ();
 b15zdnd00an1n01x5 FILLER_178_2275 ();
 b15zdnd11an1n64x5 FILLER_179_0 ();
 b15zdnd11an1n64x5 FILLER_179_64 ();
 b15zdnd11an1n64x5 FILLER_179_128 ();
 b15zdnd11an1n64x5 FILLER_179_192 ();
 b15zdnd11an1n32x5 FILLER_179_256 ();
 b15zdnd11an1n16x5 FILLER_179_288 ();
 b15zdnd11an1n08x5 FILLER_179_304 ();
 b15zdnd11an1n64x5 FILLER_179_328 ();
 b15zdnd11an1n64x5 FILLER_179_392 ();
 b15zdnd11an1n64x5 FILLER_179_456 ();
 b15zdnd11an1n64x5 FILLER_179_520 ();
 b15zdnd11an1n64x5 FILLER_179_584 ();
 b15zdnd11an1n64x5 FILLER_179_648 ();
 b15zdnd11an1n64x5 FILLER_179_712 ();
 b15zdnd11an1n64x5 FILLER_179_776 ();
 b15zdnd11an1n64x5 FILLER_179_840 ();
 b15zdnd11an1n64x5 FILLER_179_904 ();
 b15zdnd11an1n64x5 FILLER_179_968 ();
 b15zdnd11an1n04x5 FILLER_179_1032 ();
 b15zdnd00an1n01x5 FILLER_179_1036 ();
 b15zdnd11an1n64x5 FILLER_179_1040 ();
 b15zdnd11an1n64x5 FILLER_179_1104 ();
 b15zdnd11an1n32x5 FILLER_179_1168 ();
 b15zdnd11an1n16x5 FILLER_179_1200 ();
 b15zdnd11an1n04x5 FILLER_179_1216 ();
 b15zdnd11an1n64x5 FILLER_179_1262 ();
 b15zdnd11an1n64x5 FILLER_179_1326 ();
 b15zdnd11an1n64x5 FILLER_179_1390 ();
 b15zdnd11an1n32x5 FILLER_179_1454 ();
 b15zdnd11an1n04x5 FILLER_179_2257 ();
 b15zdnd00an1n01x5 FILLER_179_2261 ();
 b15zdnd11an1n16x5 FILLER_179_2266 ();
 b15zdnd00an1n02x5 FILLER_179_2282 ();
 b15zdnd11an1n64x5 FILLER_180_8 ();
 b15zdnd11an1n64x5 FILLER_180_72 ();
 b15zdnd11an1n64x5 FILLER_180_136 ();
 b15zdnd11an1n64x5 FILLER_180_200 ();
 b15zdnd11an1n64x5 FILLER_180_264 ();
 b15zdnd11an1n64x5 FILLER_180_328 ();
 b15zdnd11an1n64x5 FILLER_180_392 ();
 b15zdnd11an1n64x5 FILLER_180_456 ();
 b15zdnd11an1n64x5 FILLER_180_520 ();
 b15zdnd11an1n64x5 FILLER_180_584 ();
 b15zdnd11an1n64x5 FILLER_180_648 ();
 b15zdnd11an1n04x5 FILLER_180_712 ();
 b15zdnd00an1n02x5 FILLER_180_716 ();
 b15zdnd11an1n64x5 FILLER_180_726 ();
 b15zdnd11an1n64x5 FILLER_180_790 ();
 b15zdnd11an1n64x5 FILLER_180_854 ();
 b15zdnd11an1n64x5 FILLER_180_918 ();
 b15zdnd11an1n64x5 FILLER_180_982 ();
 b15zdnd11an1n64x5 FILLER_180_1046 ();
 b15zdnd11an1n64x5 FILLER_180_1110 ();
 b15zdnd11an1n16x5 FILLER_180_1174 ();
 b15zdnd11an1n04x5 FILLER_180_1190 ();
 b15zdnd00an1n01x5 FILLER_180_1194 ();
 b15zdnd11an1n64x5 FILLER_180_1237 ();
 b15zdnd11an1n64x5 FILLER_180_1301 ();
 b15zdnd11an1n64x5 FILLER_180_1365 ();
 b15zdnd11an1n32x5 FILLER_180_1429 ();
 b15zdnd11an1n16x5 FILLER_180_1461 ();
 b15zdnd00an1n01x5 FILLER_180_1477 ();
 b15zdnd11an1n04x5 FILLER_180_2265 ();
 b15zdnd00an1n01x5 FILLER_180_2269 ();
 b15zdnd00an1n02x5 FILLER_180_2274 ();
 b15zdnd11an1n64x5 FILLER_181_0 ();
 b15zdnd11an1n64x5 FILLER_181_64 ();
 b15zdnd11an1n64x5 FILLER_181_128 ();
 b15zdnd11an1n64x5 FILLER_181_192 ();
 b15zdnd11an1n64x5 FILLER_181_256 ();
 b15zdnd11an1n64x5 FILLER_181_320 ();
 b15zdnd11an1n64x5 FILLER_181_384 ();
 b15zdnd11an1n64x5 FILLER_181_448 ();
 b15zdnd11an1n64x5 FILLER_181_512 ();
 b15zdnd11an1n64x5 FILLER_181_576 ();
 b15zdnd11an1n64x5 FILLER_181_640 ();
 b15zdnd11an1n64x5 FILLER_181_704 ();
 b15zdnd11an1n64x5 FILLER_181_768 ();
 b15zdnd11an1n64x5 FILLER_181_832 ();
 b15zdnd11an1n64x5 FILLER_181_896 ();
 b15zdnd11an1n64x5 FILLER_181_960 ();
 b15zdnd11an1n64x5 FILLER_181_1024 ();
 b15zdnd11an1n64x5 FILLER_181_1088 ();
 b15zdnd11an1n64x5 FILLER_181_1152 ();
 b15zdnd11an1n64x5 FILLER_181_1216 ();
 b15zdnd11an1n64x5 FILLER_181_1280 ();
 b15zdnd11an1n64x5 FILLER_181_1344 ();
 b15zdnd11an1n64x5 FILLER_181_1408 ();
 b15zdnd11an1n08x5 FILLER_181_1472 ();
 b15zdnd11an1n04x5 FILLER_181_1480 ();
 b15zdnd00an1n02x5 FILLER_181_1484 ();
 b15zdnd11an1n16x5 FILLER_181_2257 ();
 b15zdnd11an1n08x5 FILLER_181_2273 ();
 b15zdnd00an1n02x5 FILLER_181_2281 ();
 b15zdnd00an1n01x5 FILLER_181_2283 ();
 b15zdnd11an1n64x5 FILLER_182_8 ();
 b15zdnd11an1n64x5 FILLER_182_72 ();
 b15zdnd11an1n64x5 FILLER_182_136 ();
 b15zdnd11an1n64x5 FILLER_182_200 ();
 b15zdnd11an1n64x5 FILLER_182_264 ();
 b15zdnd11an1n64x5 FILLER_182_328 ();
 b15zdnd11an1n32x5 FILLER_182_392 ();
 b15zdnd11an1n08x5 FILLER_182_424 ();
 b15zdnd00an1n02x5 FILLER_182_432 ();
 b15zdnd00an1n01x5 FILLER_182_434 ();
 b15zdnd11an1n64x5 FILLER_182_455 ();
 b15zdnd11an1n64x5 FILLER_182_519 ();
 b15zdnd11an1n64x5 FILLER_182_583 ();
 b15zdnd11an1n64x5 FILLER_182_647 ();
 b15zdnd11an1n04x5 FILLER_182_711 ();
 b15zdnd00an1n02x5 FILLER_182_715 ();
 b15zdnd00an1n01x5 FILLER_182_717 ();
 b15zdnd11an1n64x5 FILLER_182_726 ();
 b15zdnd11an1n64x5 FILLER_182_790 ();
 b15zdnd11an1n64x5 FILLER_182_854 ();
 b15zdnd11an1n64x5 FILLER_182_918 ();
 b15zdnd11an1n64x5 FILLER_182_982 ();
 b15zdnd11an1n64x5 FILLER_182_1046 ();
 b15zdnd11an1n64x5 FILLER_182_1110 ();
 b15zdnd11an1n64x5 FILLER_182_1174 ();
 b15zdnd11an1n64x5 FILLER_182_1238 ();
 b15zdnd11an1n32x5 FILLER_182_1302 ();
 b15zdnd11an1n16x5 FILLER_182_1334 ();
 b15zdnd00an1n02x5 FILLER_182_1350 ();
 b15zdnd11an1n64x5 FILLER_182_1355 ();
 b15zdnd11an1n32x5 FILLER_182_1419 ();
 b15zdnd11an1n16x5 FILLER_182_1451 ();
 b15zdnd11an1n08x5 FILLER_182_1467 ();
 b15zdnd00an1n02x5 FILLER_182_1475 ();
 b15zdnd00an1n01x5 FILLER_182_1477 ();
 b15zdnd11an1n08x5 FILLER_182_2265 ();
 b15zdnd00an1n02x5 FILLER_182_2273 ();
 b15zdnd00an1n01x5 FILLER_182_2275 ();
 b15zdnd11an1n64x5 FILLER_183_0 ();
 b15zdnd11an1n64x5 FILLER_183_64 ();
 b15zdnd11an1n64x5 FILLER_183_128 ();
 b15zdnd11an1n64x5 FILLER_183_192 ();
 b15zdnd11an1n64x5 FILLER_183_256 ();
 b15zdnd11an1n64x5 FILLER_183_320 ();
 b15zdnd11an1n32x5 FILLER_183_384 ();
 b15zdnd11an1n16x5 FILLER_183_416 ();
 b15zdnd11an1n08x5 FILLER_183_432 ();
 b15zdnd11an1n04x5 FILLER_183_440 ();
 b15zdnd00an1n02x5 FILLER_183_444 ();
 b15zdnd11an1n08x5 FILLER_183_449 ();
 b15zdnd11an1n04x5 FILLER_183_457 ();
 b15zdnd00an1n02x5 FILLER_183_461 ();
 b15zdnd11an1n64x5 FILLER_183_470 ();
 b15zdnd11an1n64x5 FILLER_183_534 ();
 b15zdnd11an1n32x5 FILLER_183_598 ();
 b15zdnd11an1n08x5 FILLER_183_630 ();
 b15zdnd11an1n04x5 FILLER_183_638 ();
 b15zdnd00an1n02x5 FILLER_183_642 ();
 b15zdnd00an1n01x5 FILLER_183_644 ();
 b15zdnd11an1n64x5 FILLER_183_648 ();
 b15zdnd11an1n64x5 FILLER_183_712 ();
 b15zdnd11an1n64x5 FILLER_183_776 ();
 b15zdnd11an1n64x5 FILLER_183_840 ();
 b15zdnd11an1n64x5 FILLER_183_904 ();
 b15zdnd11an1n64x5 FILLER_183_968 ();
 b15zdnd11an1n64x5 FILLER_183_1032 ();
 b15zdnd11an1n64x5 FILLER_183_1096 ();
 b15zdnd11an1n64x5 FILLER_183_1160 ();
 b15zdnd11an1n64x5 FILLER_183_1224 ();
 b15zdnd11an1n64x5 FILLER_183_1288 ();
 b15zdnd11an1n08x5 FILLER_183_1355 ();
 b15zdnd11an1n64x5 FILLER_183_1366 ();
 b15zdnd11an1n32x5 FILLER_183_1430 ();
 b15zdnd11an1n16x5 FILLER_183_1462 ();
 b15zdnd11an1n08x5 FILLER_183_1478 ();
 b15zdnd11an1n16x5 FILLER_183_2257 ();
 b15zdnd11an1n08x5 FILLER_183_2273 ();
 b15zdnd00an1n02x5 FILLER_183_2281 ();
 b15zdnd00an1n01x5 FILLER_183_2283 ();
 b15zdnd11an1n64x5 FILLER_184_8 ();
 b15zdnd11an1n64x5 FILLER_184_72 ();
 b15zdnd11an1n64x5 FILLER_184_136 ();
 b15zdnd11an1n64x5 FILLER_184_200 ();
 b15zdnd11an1n64x5 FILLER_184_264 ();
 b15zdnd11an1n64x5 FILLER_184_328 ();
 b15zdnd11an1n64x5 FILLER_184_392 ();
 b15zdnd11an1n64x5 FILLER_184_456 ();
 b15zdnd11an1n64x5 FILLER_184_520 ();
 b15zdnd11an1n16x5 FILLER_184_584 ();
 b15zdnd11an1n08x5 FILLER_184_600 ();
 b15zdnd00an1n02x5 FILLER_184_608 ();
 b15zdnd00an1n01x5 FILLER_184_610 ();
 b15zdnd11an1n04x5 FILLER_184_651 ();
 b15zdnd11an1n32x5 FILLER_184_658 ();
 b15zdnd11an1n16x5 FILLER_184_690 ();
 b15zdnd11an1n08x5 FILLER_184_706 ();
 b15zdnd11an1n04x5 FILLER_184_714 ();
 b15zdnd11an1n64x5 FILLER_184_726 ();
 b15zdnd11an1n64x5 FILLER_184_790 ();
 b15zdnd11an1n64x5 FILLER_184_854 ();
 b15zdnd11an1n64x5 FILLER_184_918 ();
 b15zdnd00an1n02x5 FILLER_184_982 ();
 b15zdnd00an1n01x5 FILLER_184_984 ();
 b15zdnd11an1n64x5 FILLER_184_996 ();
 b15zdnd11an1n64x5 FILLER_184_1060 ();
 b15zdnd11an1n64x5 FILLER_184_1124 ();
 b15zdnd11an1n64x5 FILLER_184_1188 ();
 b15zdnd11an1n64x5 FILLER_184_1252 ();
 b15zdnd11an1n08x5 FILLER_184_1316 ();
 b15zdnd11an1n04x5 FILLER_184_1324 ();
 b15zdnd00an1n01x5 FILLER_184_1328 ();
 b15zdnd11an1n64x5 FILLER_184_1381 ();
 b15zdnd11an1n32x5 FILLER_184_1445 ();
 b15zdnd00an1n01x5 FILLER_184_1477 ();
 b15zdnd11an1n08x5 FILLER_184_2265 ();
 b15zdnd00an1n02x5 FILLER_184_2273 ();
 b15zdnd00an1n01x5 FILLER_184_2275 ();
 b15zdnd11an1n64x5 FILLER_185_0 ();
 b15zdnd11an1n64x5 FILLER_185_64 ();
 b15zdnd11an1n64x5 FILLER_185_128 ();
 b15zdnd11an1n64x5 FILLER_185_192 ();
 b15zdnd11an1n64x5 FILLER_185_256 ();
 b15zdnd11an1n64x5 FILLER_185_320 ();
 b15zdnd11an1n32x5 FILLER_185_384 ();
 b15zdnd11an1n16x5 FILLER_185_416 ();
 b15zdnd11an1n08x5 FILLER_185_432 ();
 b15zdnd11an1n04x5 FILLER_185_440 ();
 b15zdnd00an1n01x5 FILLER_185_444 ();
 b15zdnd11an1n64x5 FILLER_185_487 ();
 b15zdnd11an1n64x5 FILLER_185_551 ();
 b15zdnd11an1n64x5 FILLER_185_615 ();
 b15zdnd11an1n64x5 FILLER_185_679 ();
 b15zdnd11an1n64x5 FILLER_185_743 ();
 b15zdnd11an1n64x5 FILLER_185_807 ();
 b15zdnd11an1n64x5 FILLER_185_871 ();
 b15zdnd11an1n64x5 FILLER_185_935 ();
 b15zdnd11an1n64x5 FILLER_185_999 ();
 b15zdnd11an1n64x5 FILLER_185_1063 ();
 b15zdnd11an1n64x5 FILLER_185_1127 ();
 b15zdnd11an1n64x5 FILLER_185_1191 ();
 b15zdnd11an1n64x5 FILLER_185_1255 ();
 b15zdnd11an1n64x5 FILLER_185_1319 ();
 b15zdnd11an1n64x5 FILLER_185_1383 ();
 b15zdnd11an1n32x5 FILLER_185_1447 ();
 b15zdnd11an1n04x5 FILLER_185_1479 ();
 b15zdnd00an1n02x5 FILLER_185_1483 ();
 b15zdnd00an1n01x5 FILLER_185_1485 ();
 b15zdnd11an1n16x5 FILLER_185_2257 ();
 b15zdnd11an1n08x5 FILLER_185_2273 ();
 b15zdnd00an1n02x5 FILLER_185_2281 ();
 b15zdnd00an1n01x5 FILLER_185_2283 ();
 b15zdnd11an1n64x5 FILLER_186_8 ();
 b15zdnd11an1n64x5 FILLER_186_72 ();
 b15zdnd11an1n64x5 FILLER_186_136 ();
 b15zdnd11an1n64x5 FILLER_186_200 ();
 b15zdnd11an1n64x5 FILLER_186_264 ();
 b15zdnd11an1n64x5 FILLER_186_328 ();
 b15zdnd11an1n64x5 FILLER_186_392 ();
 b15zdnd11an1n64x5 FILLER_186_456 ();
 b15zdnd11an1n64x5 FILLER_186_520 ();
 b15zdnd11an1n64x5 FILLER_186_584 ();
 b15zdnd11an1n64x5 FILLER_186_648 ();
 b15zdnd11an1n04x5 FILLER_186_712 ();
 b15zdnd00an1n02x5 FILLER_186_716 ();
 b15zdnd11an1n64x5 FILLER_186_726 ();
 b15zdnd11an1n64x5 FILLER_186_790 ();
 b15zdnd11an1n64x5 FILLER_186_854 ();
 b15zdnd11an1n64x5 FILLER_186_918 ();
 b15zdnd11an1n64x5 FILLER_186_982 ();
 b15zdnd11an1n64x5 FILLER_186_1046 ();
 b15zdnd11an1n64x5 FILLER_186_1110 ();
 b15zdnd11an1n64x5 FILLER_186_1174 ();
 b15zdnd11an1n64x5 FILLER_186_1238 ();
 b15zdnd11an1n08x5 FILLER_186_1302 ();
 b15zdnd11an1n04x5 FILLER_186_1310 ();
 b15zdnd00an1n01x5 FILLER_186_1314 ();
 b15zdnd11an1n32x5 FILLER_186_1318 ();
 b15zdnd11an1n16x5 FILLER_186_1350 ();
 b15zdnd11an1n04x5 FILLER_186_1366 ();
 b15zdnd00an1n02x5 FILLER_186_1370 ();
 b15zdnd11an1n64x5 FILLER_186_1414 ();
 b15zdnd11an1n08x5 FILLER_186_2265 ();
 b15zdnd00an1n02x5 FILLER_186_2273 ();
 b15zdnd00an1n01x5 FILLER_186_2275 ();
 b15zdnd11an1n64x5 FILLER_187_0 ();
 b15zdnd11an1n64x5 FILLER_187_64 ();
 b15zdnd11an1n64x5 FILLER_187_128 ();
 b15zdnd11an1n64x5 FILLER_187_192 ();
 b15zdnd11an1n64x5 FILLER_187_256 ();
 b15zdnd11an1n64x5 FILLER_187_320 ();
 b15zdnd11an1n64x5 FILLER_187_384 ();
 b15zdnd11an1n64x5 FILLER_187_448 ();
 b15zdnd11an1n64x5 FILLER_187_512 ();
 b15zdnd11an1n32x5 FILLER_187_576 ();
 b15zdnd00an1n02x5 FILLER_187_608 ();
 b15zdnd00an1n01x5 FILLER_187_610 ();
 b15zdnd11an1n04x5 FILLER_187_651 ();
 b15zdnd11an1n64x5 FILLER_187_658 ();
 b15zdnd11an1n64x5 FILLER_187_722 ();
 b15zdnd11an1n08x5 FILLER_187_786 ();
 b15zdnd11an1n04x5 FILLER_187_794 ();
 b15zdnd11an1n64x5 FILLER_187_801 ();
 b15zdnd11an1n64x5 FILLER_187_865 ();
 b15zdnd11an1n64x5 FILLER_187_929 ();
 b15zdnd11an1n64x5 FILLER_187_993 ();
 b15zdnd11an1n32x5 FILLER_187_1057 ();
 b15zdnd11an1n16x5 FILLER_187_1089 ();
 b15zdnd11an1n08x5 FILLER_187_1105 ();
 b15zdnd00an1n02x5 FILLER_187_1113 ();
 b15zdnd11an1n64x5 FILLER_187_1125 ();
 b15zdnd11an1n64x5 FILLER_187_1189 ();
 b15zdnd11an1n32x5 FILLER_187_1253 ();
 b15zdnd11an1n16x5 FILLER_187_1285 ();
 b15zdnd11an1n08x5 FILLER_187_1301 ();
 b15zdnd11an1n04x5 FILLER_187_1309 ();
 b15zdnd00an1n02x5 FILLER_187_1313 ();
 b15zdnd11an1n08x5 FILLER_187_1350 ();
 b15zdnd11an1n04x5 FILLER_187_1358 ();
 b15zdnd00an1n01x5 FILLER_187_1362 ();
 b15zdnd11an1n64x5 FILLER_187_1371 ();
 b15zdnd11an1n32x5 FILLER_187_1435 ();
 b15zdnd11an1n16x5 FILLER_187_1467 ();
 b15zdnd00an1n02x5 FILLER_187_1483 ();
 b15zdnd00an1n01x5 FILLER_187_1485 ();
 b15zdnd11an1n16x5 FILLER_187_2257 ();
 b15zdnd11an1n08x5 FILLER_187_2273 ();
 b15zdnd00an1n02x5 FILLER_187_2281 ();
 b15zdnd00an1n01x5 FILLER_187_2283 ();
 b15zdnd11an1n64x5 FILLER_188_8 ();
 b15zdnd11an1n64x5 FILLER_188_72 ();
 b15zdnd11an1n64x5 FILLER_188_136 ();
 b15zdnd11an1n64x5 FILLER_188_200 ();
 b15zdnd11an1n64x5 FILLER_188_264 ();
 b15zdnd11an1n64x5 FILLER_188_328 ();
 b15zdnd11an1n64x5 FILLER_188_392 ();
 b15zdnd11an1n64x5 FILLER_188_456 ();
 b15zdnd11an1n64x5 FILLER_188_520 ();
 b15zdnd11an1n64x5 FILLER_188_584 ();
 b15zdnd11an1n64x5 FILLER_188_651 ();
 b15zdnd00an1n02x5 FILLER_188_715 ();
 b15zdnd00an1n01x5 FILLER_188_717 ();
 b15zdnd11an1n32x5 FILLER_188_726 ();
 b15zdnd11an1n04x5 FILLER_188_758 ();
 b15zdnd00an1n01x5 FILLER_188_762 ();
 b15zdnd11an1n04x5 FILLER_188_803 ();
 b15zdnd11an1n16x5 FILLER_188_810 ();
 b15zdnd11an1n04x5 FILLER_188_826 ();
 b15zdnd11an1n64x5 FILLER_188_838 ();
 b15zdnd11an1n64x5 FILLER_188_902 ();
 b15zdnd11an1n64x5 FILLER_188_966 ();
 b15zdnd11an1n64x5 FILLER_188_1030 ();
 b15zdnd11an1n64x5 FILLER_188_1094 ();
 b15zdnd11an1n64x5 FILLER_188_1158 ();
 b15zdnd11an1n32x5 FILLER_188_1222 ();
 b15zdnd11an1n16x5 FILLER_188_1254 ();
 b15zdnd11an1n08x5 FILLER_188_1270 ();
 b15zdnd11an1n04x5 FILLER_188_1278 ();
 b15zdnd00an1n01x5 FILLER_188_1282 ();
 b15zdnd11an1n32x5 FILLER_188_1286 ();
 b15zdnd11an1n64x5 FILLER_188_1321 ();
 b15zdnd11an1n64x5 FILLER_188_1385 ();
 b15zdnd11an1n16x5 FILLER_188_1449 ();
 b15zdnd11an1n08x5 FILLER_188_1465 ();
 b15zdnd11an1n04x5 FILLER_188_1473 ();
 b15zdnd00an1n01x5 FILLER_188_1477 ();
 b15zdnd11an1n08x5 FILLER_188_2265 ();
 b15zdnd00an1n02x5 FILLER_188_2273 ();
 b15zdnd00an1n01x5 FILLER_188_2275 ();
 b15zdnd11an1n64x5 FILLER_189_0 ();
 b15zdnd11an1n64x5 FILLER_189_64 ();
 b15zdnd11an1n64x5 FILLER_189_128 ();
 b15zdnd11an1n64x5 FILLER_189_192 ();
 b15zdnd11an1n64x5 FILLER_189_256 ();
 b15zdnd11an1n64x5 FILLER_189_320 ();
 b15zdnd11an1n64x5 FILLER_189_384 ();
 b15zdnd11an1n64x5 FILLER_189_448 ();
 b15zdnd11an1n16x5 FILLER_189_512 ();
 b15zdnd11an1n08x5 FILLER_189_528 ();
 b15zdnd11an1n64x5 FILLER_189_578 ();
 b15zdnd11an1n64x5 FILLER_189_642 ();
 b15zdnd11an1n32x5 FILLER_189_706 ();
 b15zdnd11an1n16x5 FILLER_189_738 ();
 b15zdnd11an1n04x5 FILLER_189_754 ();
 b15zdnd11an1n04x5 FILLER_189_798 ();
 b15zdnd11an1n64x5 FILLER_189_805 ();
 b15zdnd11an1n64x5 FILLER_189_869 ();
 b15zdnd11an1n64x5 FILLER_189_933 ();
 b15zdnd11an1n64x5 FILLER_189_997 ();
 b15zdnd11an1n64x5 FILLER_189_1061 ();
 b15zdnd11an1n64x5 FILLER_189_1125 ();
 b15zdnd11an1n64x5 FILLER_189_1189 ();
 b15zdnd11an1n16x5 FILLER_189_1253 ();
 b15zdnd11an1n08x5 FILLER_189_1269 ();
 b15zdnd11an1n04x5 FILLER_189_1277 ();
 b15zdnd00an1n02x5 FILLER_189_1281 ();
 b15zdnd11an1n64x5 FILLER_189_1318 ();
 b15zdnd11an1n64x5 FILLER_189_1382 ();
 b15zdnd11an1n32x5 FILLER_189_1446 ();
 b15zdnd11an1n08x5 FILLER_189_1478 ();
 b15zdnd11an1n16x5 FILLER_189_2257 ();
 b15zdnd11an1n08x5 FILLER_189_2273 ();
 b15zdnd00an1n02x5 FILLER_189_2281 ();
 b15zdnd00an1n01x5 FILLER_189_2283 ();
 b15zdnd11an1n64x5 FILLER_190_8 ();
 b15zdnd11an1n64x5 FILLER_190_72 ();
 b15zdnd11an1n64x5 FILLER_190_136 ();
 b15zdnd11an1n64x5 FILLER_190_200 ();
 b15zdnd11an1n64x5 FILLER_190_264 ();
 b15zdnd11an1n64x5 FILLER_190_328 ();
 b15zdnd11an1n64x5 FILLER_190_392 ();
 b15zdnd11an1n64x5 FILLER_190_456 ();
 b15zdnd11an1n64x5 FILLER_190_520 ();
 b15zdnd11an1n64x5 FILLER_190_584 ();
 b15zdnd11an1n64x5 FILLER_190_648 ();
 b15zdnd11an1n04x5 FILLER_190_712 ();
 b15zdnd00an1n02x5 FILLER_190_716 ();
 b15zdnd11an1n04x5 FILLER_190_726 ();
 b15zdnd11an1n32x5 FILLER_190_737 ();
 b15zdnd00an1n01x5 FILLER_190_769 ();
 b15zdnd11an1n16x5 FILLER_190_773 ();
 b15zdnd11an1n08x5 FILLER_190_792 ();
 b15zdnd11an1n04x5 FILLER_190_800 ();
 b15zdnd00an1n02x5 FILLER_190_804 ();
 b15zdnd11an1n64x5 FILLER_190_820 ();
 b15zdnd11an1n64x5 FILLER_190_884 ();
 b15zdnd11an1n64x5 FILLER_190_948 ();
 b15zdnd11an1n64x5 FILLER_190_1012 ();
 b15zdnd11an1n64x5 FILLER_190_1076 ();
 b15zdnd11an1n64x5 FILLER_190_1140 ();
 b15zdnd11an1n32x5 FILLER_190_1204 ();
 b15zdnd00an1n02x5 FILLER_190_1236 ();
 b15zdnd00an1n01x5 FILLER_190_1238 ();
 b15zdnd11an1n04x5 FILLER_190_1242 ();
 b15zdnd11an1n04x5 FILLER_190_1281 ();
 b15zdnd11an1n64x5 FILLER_190_1288 ();
 b15zdnd11an1n64x5 FILLER_190_1352 ();
 b15zdnd11an1n32x5 FILLER_190_1416 ();
 b15zdnd11an1n16x5 FILLER_190_1448 ();
 b15zdnd11an1n08x5 FILLER_190_1464 ();
 b15zdnd11an1n04x5 FILLER_190_1472 ();
 b15zdnd00an1n02x5 FILLER_190_1476 ();
 b15zdnd11an1n08x5 FILLER_190_2265 ();
 b15zdnd00an1n02x5 FILLER_190_2273 ();
 b15zdnd00an1n01x5 FILLER_190_2275 ();
 b15zdnd11an1n64x5 FILLER_191_0 ();
 b15zdnd11an1n64x5 FILLER_191_64 ();
 b15zdnd11an1n64x5 FILLER_191_128 ();
 b15zdnd11an1n64x5 FILLER_191_192 ();
 b15zdnd11an1n64x5 FILLER_191_256 ();
 b15zdnd11an1n64x5 FILLER_191_320 ();
 b15zdnd11an1n64x5 FILLER_191_384 ();
 b15zdnd11an1n64x5 FILLER_191_448 ();
 b15zdnd11an1n64x5 FILLER_191_512 ();
 b15zdnd11an1n64x5 FILLER_191_576 ();
 b15zdnd11an1n64x5 FILLER_191_640 ();
 b15zdnd11an1n16x5 FILLER_191_704 ();
 b15zdnd11an1n08x5 FILLER_191_720 ();
 b15zdnd11an1n04x5 FILLER_191_728 ();
 b15zdnd00an1n02x5 FILLER_191_732 ();
 b15zdnd00an1n01x5 FILLER_191_734 ();
 b15zdnd11an1n04x5 FILLER_191_775 ();
 b15zdnd00an1n02x5 FILLER_191_779 ();
 b15zdnd11an1n64x5 FILLER_191_784 ();
 b15zdnd11an1n64x5 FILLER_191_848 ();
 b15zdnd11an1n64x5 FILLER_191_912 ();
 b15zdnd11an1n64x5 FILLER_191_976 ();
 b15zdnd11an1n64x5 FILLER_191_1040 ();
 b15zdnd11an1n64x5 FILLER_191_1104 ();
 b15zdnd11an1n64x5 FILLER_191_1168 ();
 b15zdnd11an1n08x5 FILLER_191_1232 ();
 b15zdnd11an1n04x5 FILLER_191_1240 ();
 b15zdnd00an1n02x5 FILLER_191_1244 ();
 b15zdnd00an1n01x5 FILLER_191_1246 ();
 b15zdnd11an1n64x5 FILLER_191_1250 ();
 b15zdnd11an1n64x5 FILLER_191_1314 ();
 b15zdnd11an1n64x5 FILLER_191_1378 ();
 b15zdnd11an1n32x5 FILLER_191_1442 ();
 b15zdnd11an1n08x5 FILLER_191_1474 ();
 b15zdnd11an1n04x5 FILLER_191_1482 ();
 b15zdnd11an1n16x5 FILLER_191_2257 ();
 b15zdnd11an1n08x5 FILLER_191_2273 ();
 b15zdnd00an1n02x5 FILLER_191_2281 ();
 b15zdnd00an1n01x5 FILLER_191_2283 ();
 b15zdnd11an1n64x5 FILLER_192_8 ();
 b15zdnd11an1n64x5 FILLER_192_72 ();
 b15zdnd11an1n64x5 FILLER_192_136 ();
 b15zdnd11an1n64x5 FILLER_192_200 ();
 b15zdnd11an1n64x5 FILLER_192_264 ();
 b15zdnd11an1n64x5 FILLER_192_328 ();
 b15zdnd11an1n64x5 FILLER_192_392 ();
 b15zdnd11an1n64x5 FILLER_192_456 ();
 b15zdnd11an1n64x5 FILLER_192_520 ();
 b15zdnd11an1n64x5 FILLER_192_584 ();
 b15zdnd11an1n64x5 FILLER_192_648 ();
 b15zdnd11an1n04x5 FILLER_192_712 ();
 b15zdnd00an1n02x5 FILLER_192_716 ();
 b15zdnd11an1n32x5 FILLER_192_726 ();
 b15zdnd00an1n02x5 FILLER_192_758 ();
 b15zdnd11an1n64x5 FILLER_192_802 ();
 b15zdnd11an1n64x5 FILLER_192_866 ();
 b15zdnd11an1n64x5 FILLER_192_930 ();
 b15zdnd11an1n64x5 FILLER_192_994 ();
 b15zdnd11an1n64x5 FILLER_192_1058 ();
 b15zdnd11an1n64x5 FILLER_192_1122 ();
 b15zdnd11an1n32x5 FILLER_192_1186 ();
 b15zdnd11an1n04x5 FILLER_192_1218 ();
 b15zdnd00an1n02x5 FILLER_192_1222 ();
 b15zdnd11an1n64x5 FILLER_192_1244 ();
 b15zdnd11an1n64x5 FILLER_192_1308 ();
 b15zdnd11an1n64x5 FILLER_192_1372 ();
 b15zdnd11an1n32x5 FILLER_192_1436 ();
 b15zdnd11an1n08x5 FILLER_192_1468 ();
 b15zdnd00an1n02x5 FILLER_192_1476 ();
 b15zdnd11an1n08x5 FILLER_192_2265 ();
 b15zdnd00an1n02x5 FILLER_192_2273 ();
 b15zdnd00an1n01x5 FILLER_192_2275 ();
 b15zdnd11an1n64x5 FILLER_193_0 ();
 b15zdnd11an1n64x5 FILLER_193_64 ();
 b15zdnd11an1n64x5 FILLER_193_128 ();
 b15zdnd11an1n64x5 FILLER_193_192 ();
 b15zdnd11an1n64x5 FILLER_193_256 ();
 b15zdnd11an1n64x5 FILLER_193_320 ();
 b15zdnd11an1n64x5 FILLER_193_384 ();
 b15zdnd11an1n64x5 FILLER_193_448 ();
 b15zdnd11an1n64x5 FILLER_193_512 ();
 b15zdnd11an1n64x5 FILLER_193_576 ();
 b15zdnd11an1n08x5 FILLER_193_640 ();
 b15zdnd00an1n01x5 FILLER_193_648 ();
 b15zdnd11an1n64x5 FILLER_193_652 ();
 b15zdnd11an1n64x5 FILLER_193_716 ();
 b15zdnd11an1n64x5 FILLER_193_780 ();
 b15zdnd11an1n64x5 FILLER_193_844 ();
 b15zdnd11an1n64x5 FILLER_193_908 ();
 b15zdnd11an1n64x5 FILLER_193_972 ();
 b15zdnd11an1n64x5 FILLER_193_1036 ();
 b15zdnd11an1n64x5 FILLER_193_1100 ();
 b15zdnd11an1n64x5 FILLER_193_1164 ();
 b15zdnd11an1n64x5 FILLER_193_1228 ();
 b15zdnd11an1n64x5 FILLER_193_1292 ();
 b15zdnd11an1n64x5 FILLER_193_1356 ();
 b15zdnd11an1n64x5 FILLER_193_1420 ();
 b15zdnd00an1n02x5 FILLER_193_1484 ();
 b15zdnd11an1n16x5 FILLER_193_2257 ();
 b15zdnd11an1n08x5 FILLER_193_2273 ();
 b15zdnd00an1n02x5 FILLER_193_2281 ();
 b15zdnd00an1n01x5 FILLER_193_2283 ();
 b15zdnd11an1n64x5 FILLER_194_8 ();
 b15zdnd11an1n64x5 FILLER_194_72 ();
 b15zdnd11an1n64x5 FILLER_194_136 ();
 b15zdnd11an1n64x5 FILLER_194_200 ();
 b15zdnd11an1n64x5 FILLER_194_264 ();
 b15zdnd11an1n64x5 FILLER_194_328 ();
 b15zdnd11an1n64x5 FILLER_194_392 ();
 b15zdnd11an1n64x5 FILLER_194_456 ();
 b15zdnd11an1n64x5 FILLER_194_520 ();
 b15zdnd11an1n32x5 FILLER_194_584 ();
 b15zdnd00an1n01x5 FILLER_194_616 ();
 b15zdnd11an1n04x5 FILLER_194_657 ();
 b15zdnd11an1n32x5 FILLER_194_664 ();
 b15zdnd11an1n16x5 FILLER_194_696 ();
 b15zdnd11an1n04x5 FILLER_194_712 ();
 b15zdnd00an1n02x5 FILLER_194_716 ();
 b15zdnd11an1n32x5 FILLER_194_726 ();
 b15zdnd11an1n64x5 FILLER_194_766 ();
 b15zdnd11an1n64x5 FILLER_194_830 ();
 b15zdnd11an1n64x5 FILLER_194_894 ();
 b15zdnd11an1n64x5 FILLER_194_958 ();
 b15zdnd11an1n64x5 FILLER_194_1022 ();
 b15zdnd11an1n64x5 FILLER_194_1086 ();
 b15zdnd11an1n64x5 FILLER_194_1150 ();
 b15zdnd11an1n64x5 FILLER_194_1214 ();
 b15zdnd11an1n64x5 FILLER_194_1278 ();
 b15zdnd11an1n64x5 FILLER_194_1342 ();
 b15zdnd11an1n64x5 FILLER_194_1406 ();
 b15zdnd11an1n08x5 FILLER_194_1470 ();
 b15zdnd11an1n08x5 FILLER_194_2265 ();
 b15zdnd00an1n02x5 FILLER_194_2273 ();
 b15zdnd00an1n01x5 FILLER_194_2275 ();
 b15zdnd11an1n64x5 FILLER_195_0 ();
 b15zdnd11an1n64x5 FILLER_195_64 ();
 b15zdnd11an1n64x5 FILLER_195_128 ();
 b15zdnd11an1n64x5 FILLER_195_192 ();
 b15zdnd11an1n64x5 FILLER_195_256 ();
 b15zdnd11an1n64x5 FILLER_195_320 ();
 b15zdnd11an1n64x5 FILLER_195_384 ();
 b15zdnd11an1n08x5 FILLER_195_448 ();
 b15zdnd11an1n64x5 FILLER_195_466 ();
 b15zdnd11an1n64x5 FILLER_195_530 ();
 b15zdnd11an1n64x5 FILLER_195_594 ();
 b15zdnd11an1n64x5 FILLER_195_658 ();
 b15zdnd11an1n64x5 FILLER_195_722 ();
 b15zdnd11an1n64x5 FILLER_195_786 ();
 b15zdnd11an1n64x5 FILLER_195_850 ();
 b15zdnd11an1n64x5 FILLER_195_914 ();
 b15zdnd11an1n64x5 FILLER_195_978 ();
 b15zdnd11an1n64x5 FILLER_195_1042 ();
 b15zdnd11an1n64x5 FILLER_195_1106 ();
 b15zdnd11an1n64x5 FILLER_195_1170 ();
 b15zdnd11an1n64x5 FILLER_195_1234 ();
 b15zdnd11an1n64x5 FILLER_195_1298 ();
 b15zdnd11an1n64x5 FILLER_195_1362 ();
 b15zdnd11an1n32x5 FILLER_195_1426 ();
 b15zdnd11an1n16x5 FILLER_195_1458 ();
 b15zdnd11an1n08x5 FILLER_195_1474 ();
 b15zdnd11an1n04x5 FILLER_195_1482 ();
 b15zdnd11an1n16x5 FILLER_195_2257 ();
 b15zdnd11an1n08x5 FILLER_195_2273 ();
 b15zdnd00an1n02x5 FILLER_195_2281 ();
 b15zdnd00an1n01x5 FILLER_195_2283 ();
 b15zdnd11an1n16x5 FILLER_196_8 ();
 b15zdnd00an1n01x5 FILLER_196_24 ();
 b15zdnd11an1n64x5 FILLER_196_29 ();
 b15zdnd11an1n64x5 FILLER_196_93 ();
 b15zdnd11an1n64x5 FILLER_196_157 ();
 b15zdnd11an1n64x5 FILLER_196_221 ();
 b15zdnd11an1n64x5 FILLER_196_285 ();
 b15zdnd11an1n64x5 FILLER_196_349 ();
 b15zdnd11an1n16x5 FILLER_196_413 ();
 b15zdnd11an1n04x5 FILLER_196_432 ();
 b15zdnd00an1n02x5 FILLER_196_436 ();
 b15zdnd11an1n64x5 FILLER_196_480 ();
 b15zdnd11an1n64x5 FILLER_196_544 ();
 b15zdnd11an1n64x5 FILLER_196_608 ();
 b15zdnd11an1n32x5 FILLER_196_672 ();
 b15zdnd11an1n08x5 FILLER_196_704 ();
 b15zdnd11an1n04x5 FILLER_196_712 ();
 b15zdnd00an1n02x5 FILLER_196_716 ();
 b15zdnd11an1n64x5 FILLER_196_726 ();
 b15zdnd11an1n64x5 FILLER_196_790 ();
 b15zdnd11an1n64x5 FILLER_196_854 ();
 b15zdnd11an1n64x5 FILLER_196_918 ();
 b15zdnd11an1n64x5 FILLER_196_982 ();
 b15zdnd11an1n64x5 FILLER_196_1046 ();
 b15zdnd11an1n64x5 FILLER_196_1110 ();
 b15zdnd11an1n64x5 FILLER_196_1174 ();
 b15zdnd11an1n64x5 FILLER_196_1238 ();
 b15zdnd11an1n64x5 FILLER_196_1302 ();
 b15zdnd11an1n64x5 FILLER_196_1366 ();
 b15zdnd11an1n32x5 FILLER_196_1430 ();
 b15zdnd11an1n16x5 FILLER_196_1462 ();
 b15zdnd11an1n08x5 FILLER_196_2265 ();
 b15zdnd00an1n02x5 FILLER_196_2273 ();
 b15zdnd00an1n01x5 FILLER_196_2275 ();
 b15zdnd11an1n08x5 FILLER_197_0 ();
 b15zdnd11an1n64x5 FILLER_197_50 ();
 b15zdnd11an1n64x5 FILLER_197_114 ();
 b15zdnd11an1n64x5 FILLER_197_178 ();
 b15zdnd11an1n64x5 FILLER_197_242 ();
 b15zdnd11an1n64x5 FILLER_197_306 ();
 b15zdnd11an1n64x5 FILLER_197_370 ();
 b15zdnd11an1n64x5 FILLER_197_434 ();
 b15zdnd11an1n64x5 FILLER_197_498 ();
 b15zdnd11an1n64x5 FILLER_197_562 ();
 b15zdnd11an1n64x5 FILLER_197_626 ();
 b15zdnd11an1n64x5 FILLER_197_690 ();
 b15zdnd11an1n64x5 FILLER_197_754 ();
 b15zdnd11an1n64x5 FILLER_197_818 ();
 b15zdnd11an1n64x5 FILLER_197_882 ();
 b15zdnd11an1n64x5 FILLER_197_946 ();
 b15zdnd11an1n64x5 FILLER_197_1010 ();
 b15zdnd11an1n64x5 FILLER_197_1074 ();
 b15zdnd11an1n64x5 FILLER_197_1138 ();
 b15zdnd00an1n02x5 FILLER_197_1202 ();
 b15zdnd00an1n01x5 FILLER_197_1204 ();
 b15zdnd11an1n64x5 FILLER_197_1247 ();
 b15zdnd11an1n64x5 FILLER_197_1311 ();
 b15zdnd11an1n64x5 FILLER_197_1375 ();
 b15zdnd11an1n32x5 FILLER_197_1439 ();
 b15zdnd11an1n08x5 FILLER_197_1471 ();
 b15zdnd11an1n04x5 FILLER_197_1479 ();
 b15zdnd00an1n02x5 FILLER_197_1483 ();
 b15zdnd00an1n01x5 FILLER_197_1485 ();
 b15zdnd11an1n16x5 FILLER_197_2257 ();
 b15zdnd11an1n08x5 FILLER_197_2273 ();
 b15zdnd00an1n02x5 FILLER_197_2281 ();
 b15zdnd00an1n01x5 FILLER_197_2283 ();
 b15zdnd00an1n02x5 FILLER_198_8 ();
 b15zdnd11an1n64x5 FILLER_198_52 ();
 b15zdnd11an1n64x5 FILLER_198_116 ();
 b15zdnd11an1n64x5 FILLER_198_180 ();
 b15zdnd11an1n64x5 FILLER_198_244 ();
 b15zdnd11an1n64x5 FILLER_198_308 ();
 b15zdnd11an1n64x5 FILLER_198_372 ();
 b15zdnd11an1n64x5 FILLER_198_436 ();
 b15zdnd11an1n64x5 FILLER_198_500 ();
 b15zdnd11an1n64x5 FILLER_198_564 ();
 b15zdnd11an1n64x5 FILLER_198_628 ();
 b15zdnd11an1n16x5 FILLER_198_692 ();
 b15zdnd11an1n08x5 FILLER_198_708 ();
 b15zdnd00an1n02x5 FILLER_198_716 ();
 b15zdnd11an1n64x5 FILLER_198_726 ();
 b15zdnd11an1n64x5 FILLER_198_790 ();
 b15zdnd11an1n64x5 FILLER_198_854 ();
 b15zdnd11an1n64x5 FILLER_198_918 ();
 b15zdnd11an1n64x5 FILLER_198_982 ();
 b15zdnd11an1n64x5 FILLER_198_1046 ();
 b15zdnd11an1n32x5 FILLER_198_1110 ();
 b15zdnd11an1n16x5 FILLER_198_1142 ();
 b15zdnd11an1n08x5 FILLER_198_1158 ();
 b15zdnd11an1n04x5 FILLER_198_1166 ();
 b15zdnd11an1n64x5 FILLER_198_1212 ();
 b15zdnd11an1n64x5 FILLER_198_1276 ();
 b15zdnd11an1n64x5 FILLER_198_1340 ();
 b15zdnd11an1n32x5 FILLER_198_1404 ();
 b15zdnd11an1n64x5 FILLER_198_1444 ();
 b15zdnd11an1n32x5 FILLER_198_1508 ();
 b15zdnd00an1n01x5 FILLER_198_1540 ();
 b15zdnd11an1n04x5 FILLER_198_1573 ();
 b15zdnd11an1n64x5 FILLER_198_1580 ();
 b15zdnd11an1n64x5 FILLER_198_1644 ();
 b15zdnd11an1n64x5 FILLER_198_1708 ();
 b15zdnd11an1n08x5 FILLER_198_1772 ();
 b15zdnd11an1n04x5 FILLER_198_1780 ();
 b15zdnd11an1n04x5 FILLER_198_1826 ();
 b15zdnd11an1n04x5 FILLER_198_1833 ();
 b15zdnd11an1n64x5 FILLER_198_1840 ();
 b15zdnd11an1n64x5 FILLER_198_1904 ();
 b15zdnd11an1n64x5 FILLER_198_1968 ();
 b15zdnd11an1n64x5 FILLER_198_2032 ();
 b15zdnd11an1n32x5 FILLER_198_2096 ();
 b15zdnd11an1n16x5 FILLER_198_2128 ();
 b15zdnd11an1n08x5 FILLER_198_2144 ();
 b15zdnd00an1n02x5 FILLER_198_2152 ();
 b15zdnd11an1n64x5 FILLER_198_2162 ();
 b15zdnd11an1n32x5 FILLER_198_2226 ();
 b15zdnd11an1n16x5 FILLER_198_2258 ();
 b15zdnd00an1n02x5 FILLER_198_2274 ();
 b15zdnd11an1n04x5 FILLER_199_0 ();
 b15zdnd00an1n02x5 FILLER_199_4 ();
 b15zdnd00an1n01x5 FILLER_199_6 ();
 b15zdnd11an1n08x5 FILLER_199_11 ();
 b15zdnd11an1n64x5 FILLER_199_23 ();
 b15zdnd11an1n64x5 FILLER_199_87 ();
 b15zdnd11an1n64x5 FILLER_199_151 ();
 b15zdnd11an1n16x5 FILLER_199_215 ();
 b15zdnd11an1n64x5 FILLER_199_273 ();
 b15zdnd11an1n64x5 FILLER_199_337 ();
 b15zdnd11an1n16x5 FILLER_199_401 ();
 b15zdnd00an1n02x5 FILLER_199_417 ();
 b15zdnd00an1n01x5 FILLER_199_419 ();
 b15zdnd11an1n64x5 FILLER_199_436 ();
 b15zdnd11an1n64x5 FILLER_199_500 ();
 b15zdnd11an1n64x5 FILLER_199_564 ();
 b15zdnd11an1n64x5 FILLER_199_628 ();
 b15zdnd11an1n64x5 FILLER_199_692 ();
 b15zdnd11an1n32x5 FILLER_199_756 ();
 b15zdnd11an1n64x5 FILLER_199_830 ();
 b15zdnd11an1n64x5 FILLER_199_894 ();
 b15zdnd11an1n32x5 FILLER_199_958 ();
 b15zdnd11an1n08x5 FILLER_199_990 ();
 b15zdnd00an1n02x5 FILLER_199_998 ();
 b15zdnd11an1n64x5 FILLER_199_1042 ();
 b15zdnd11an1n64x5 FILLER_199_1106 ();
 b15zdnd11an1n64x5 FILLER_199_1170 ();
 b15zdnd11an1n64x5 FILLER_199_1234 ();
 b15zdnd11an1n64x5 FILLER_199_1298 ();
 b15zdnd11an1n64x5 FILLER_199_1362 ();
 b15zdnd11an1n64x5 FILLER_199_1426 ();
 b15zdnd11an1n64x5 FILLER_199_1490 ();
 b15zdnd11an1n08x5 FILLER_199_1554 ();
 b15zdnd11an1n04x5 FILLER_199_1562 ();
 b15zdnd00an1n01x5 FILLER_199_1566 ();
 b15zdnd11an1n04x5 FILLER_199_1570 ();
 b15zdnd11an1n64x5 FILLER_199_1577 ();
 b15zdnd11an1n64x5 FILLER_199_1641 ();
 b15zdnd11an1n32x5 FILLER_199_1705 ();
 b15zdnd11an1n16x5 FILLER_199_1737 ();
 b15zdnd11an1n08x5 FILLER_199_1753 ();
 b15zdnd11an1n04x5 FILLER_199_1761 ();
 b15zdnd11an1n04x5 FILLER_199_1773 ();
 b15zdnd11an1n04x5 FILLER_199_1819 ();
 b15zdnd00an1n01x5 FILLER_199_1823 ();
 b15zdnd11an1n04x5 FILLER_199_1827 ();
 b15zdnd11an1n64x5 FILLER_199_1834 ();
 b15zdnd11an1n64x5 FILLER_199_1898 ();
 b15zdnd11an1n64x5 FILLER_199_1962 ();
 b15zdnd11an1n64x5 FILLER_199_2026 ();
 b15zdnd11an1n64x5 FILLER_199_2090 ();
 b15zdnd11an1n32x5 FILLER_199_2154 ();
 b15zdnd11an1n16x5 FILLER_199_2186 ();
 b15zdnd11an1n04x5 FILLER_199_2202 ();
 b15zdnd00an1n02x5 FILLER_199_2206 ();
 b15zdnd00an1n01x5 FILLER_199_2208 ();
 b15zdnd11an1n32x5 FILLER_199_2251 ();
 b15zdnd00an1n01x5 FILLER_199_2283 ();
 b15zdnd00an1n02x5 FILLER_200_8 ();
 b15zdnd11an1n64x5 FILLER_200_52 ();
 b15zdnd11an1n64x5 FILLER_200_116 ();
 b15zdnd11an1n32x5 FILLER_200_180 ();
 b15zdnd11an1n04x5 FILLER_200_212 ();
 b15zdnd11an1n64x5 FILLER_200_258 ();
 b15zdnd11an1n64x5 FILLER_200_322 ();
 b15zdnd11an1n64x5 FILLER_200_386 ();
 b15zdnd11an1n64x5 FILLER_200_450 ();
 b15zdnd11an1n64x5 FILLER_200_514 ();
 b15zdnd11an1n64x5 FILLER_200_578 ();
 b15zdnd11an1n64x5 FILLER_200_642 ();
 b15zdnd11an1n08x5 FILLER_200_706 ();
 b15zdnd11an1n04x5 FILLER_200_714 ();
 b15zdnd11an1n64x5 FILLER_200_726 ();
 b15zdnd11an1n64x5 FILLER_200_790 ();
 b15zdnd11an1n16x5 FILLER_200_854 ();
 b15zdnd11an1n08x5 FILLER_200_870 ();
 b15zdnd11an1n04x5 FILLER_200_878 ();
 b15zdnd00an1n02x5 FILLER_200_882 ();
 b15zdnd11an1n64x5 FILLER_200_895 ();
 b15zdnd11an1n64x5 FILLER_200_959 ();
 b15zdnd11an1n64x5 FILLER_200_1023 ();
 b15zdnd11an1n64x5 FILLER_200_1087 ();
 b15zdnd11an1n64x5 FILLER_200_1151 ();
 b15zdnd11an1n32x5 FILLER_200_1215 ();
 b15zdnd11an1n08x5 FILLER_200_1247 ();
 b15zdnd11an1n04x5 FILLER_200_1255 ();
 b15zdnd11an1n08x5 FILLER_200_1279 ();
 b15zdnd11an1n04x5 FILLER_200_1287 ();
 b15zdnd00an1n02x5 FILLER_200_1291 ();
 b15zdnd11an1n32x5 FILLER_200_1299 ();
 b15zdnd00an1n01x5 FILLER_200_1331 ();
 b15zdnd11an1n64x5 FILLER_200_1374 ();
 b15zdnd11an1n64x5 FILLER_200_1438 ();
 b15zdnd11an1n64x5 FILLER_200_1502 ();
 b15zdnd11an1n64x5 FILLER_200_1566 ();
 b15zdnd11an1n64x5 FILLER_200_1630 ();
 b15zdnd11an1n64x5 FILLER_200_1694 ();
 b15zdnd11an1n16x5 FILLER_200_1758 ();
 b15zdnd00an1n02x5 FILLER_200_1774 ();
 b15zdnd00an1n01x5 FILLER_200_1776 ();
 b15zdnd11an1n04x5 FILLER_200_1783 ();
 b15zdnd11an1n04x5 FILLER_200_1819 ();
 b15zdnd11an1n04x5 FILLER_200_1826 ();
 b15zdnd11an1n64x5 FILLER_200_1833 ();
 b15zdnd11an1n64x5 FILLER_200_1897 ();
 b15zdnd11an1n64x5 FILLER_200_1961 ();
 b15zdnd11an1n64x5 FILLER_200_2025 ();
 b15zdnd11an1n64x5 FILLER_200_2089 ();
 b15zdnd00an1n01x5 FILLER_200_2153 ();
 b15zdnd11an1n64x5 FILLER_200_2162 ();
 b15zdnd11an1n32x5 FILLER_200_2226 ();
 b15zdnd11an1n16x5 FILLER_200_2258 ();
 b15zdnd00an1n02x5 FILLER_200_2274 ();
 b15zdnd11an1n64x5 FILLER_201_0 ();
 b15zdnd11an1n64x5 FILLER_201_64 ();
 b15zdnd11an1n64x5 FILLER_201_128 ();
 b15zdnd11an1n64x5 FILLER_201_192 ();
 b15zdnd11an1n64x5 FILLER_201_256 ();
 b15zdnd11an1n64x5 FILLER_201_320 ();
 b15zdnd11an1n32x5 FILLER_201_384 ();
 b15zdnd11an1n04x5 FILLER_201_416 ();
 b15zdnd00an1n02x5 FILLER_201_420 ();
 b15zdnd00an1n01x5 FILLER_201_422 ();
 b15zdnd11an1n64x5 FILLER_201_437 ();
 b15zdnd11an1n64x5 FILLER_201_501 ();
 b15zdnd11an1n64x5 FILLER_201_565 ();
 b15zdnd11an1n64x5 FILLER_201_629 ();
 b15zdnd11an1n64x5 FILLER_201_693 ();
 b15zdnd11an1n64x5 FILLER_201_757 ();
 b15zdnd11an1n64x5 FILLER_201_821 ();
 b15zdnd11an1n64x5 FILLER_201_885 ();
 b15zdnd11an1n64x5 FILLER_201_949 ();
 b15zdnd11an1n64x5 FILLER_201_1013 ();
 b15zdnd11an1n16x5 FILLER_201_1077 ();
 b15zdnd11an1n04x5 FILLER_201_1093 ();
 b15zdnd00an1n02x5 FILLER_201_1097 ();
 b15zdnd00an1n01x5 FILLER_201_1099 ();
 b15zdnd11an1n64x5 FILLER_201_1142 ();
 b15zdnd11an1n64x5 FILLER_201_1206 ();
 b15zdnd11an1n64x5 FILLER_201_1270 ();
 b15zdnd11an1n08x5 FILLER_201_1334 ();
 b15zdnd11an1n64x5 FILLER_201_1384 ();
 b15zdnd11an1n64x5 FILLER_201_1448 ();
 b15zdnd11an1n64x5 FILLER_201_1512 ();
 b15zdnd11an1n64x5 FILLER_201_1576 ();
 b15zdnd11an1n64x5 FILLER_201_1640 ();
 b15zdnd11an1n64x5 FILLER_201_1704 ();
 b15zdnd11an1n16x5 FILLER_201_1768 ();
 b15zdnd11an1n04x5 FILLER_201_1784 ();
 b15zdnd11an1n64x5 FILLER_201_1820 ();
 b15zdnd11an1n64x5 FILLER_201_1884 ();
 b15zdnd11an1n64x5 FILLER_201_1948 ();
 b15zdnd11an1n64x5 FILLER_201_2012 ();
 b15zdnd11an1n64x5 FILLER_201_2076 ();
 b15zdnd11an1n64x5 FILLER_201_2140 ();
 b15zdnd11an1n64x5 FILLER_201_2204 ();
 b15zdnd11an1n16x5 FILLER_201_2268 ();
 b15zdnd11an1n64x5 FILLER_202_8 ();
 b15zdnd11an1n64x5 FILLER_202_72 ();
 b15zdnd11an1n64x5 FILLER_202_136 ();
 b15zdnd11an1n64x5 FILLER_202_200 ();
 b15zdnd11an1n64x5 FILLER_202_264 ();
 b15zdnd11an1n64x5 FILLER_202_328 ();
 b15zdnd11an1n32x5 FILLER_202_392 ();
 b15zdnd00an1n02x5 FILLER_202_424 ();
 b15zdnd11an1n64x5 FILLER_202_457 ();
 b15zdnd11an1n64x5 FILLER_202_521 ();
 b15zdnd11an1n64x5 FILLER_202_585 ();
 b15zdnd11an1n64x5 FILLER_202_649 ();
 b15zdnd11an1n04x5 FILLER_202_713 ();
 b15zdnd00an1n01x5 FILLER_202_717 ();
 b15zdnd11an1n64x5 FILLER_202_726 ();
 b15zdnd11an1n64x5 FILLER_202_790 ();
 b15zdnd11an1n64x5 FILLER_202_854 ();
 b15zdnd11an1n64x5 FILLER_202_918 ();
 b15zdnd11an1n64x5 FILLER_202_982 ();
 b15zdnd11an1n64x5 FILLER_202_1046 ();
 b15zdnd11an1n32x5 FILLER_202_1110 ();
 b15zdnd11an1n16x5 FILLER_202_1142 ();
 b15zdnd11an1n08x5 FILLER_202_1158 ();
 b15zdnd11an1n04x5 FILLER_202_1166 ();
 b15zdnd11an1n32x5 FILLER_202_1212 ();
 b15zdnd11an1n08x5 FILLER_202_1244 ();
 b15zdnd00an1n01x5 FILLER_202_1252 ();
 b15zdnd11an1n64x5 FILLER_202_1295 ();
 b15zdnd11an1n64x5 FILLER_202_1359 ();
 b15zdnd11an1n64x5 FILLER_202_1423 ();
 b15zdnd11an1n64x5 FILLER_202_1487 ();
 b15zdnd11an1n64x5 FILLER_202_1551 ();
 b15zdnd11an1n64x5 FILLER_202_1615 ();
 b15zdnd11an1n64x5 FILLER_202_1679 ();
 b15zdnd11an1n64x5 FILLER_202_1743 ();
 b15zdnd11an1n64x5 FILLER_202_1807 ();
 b15zdnd11an1n64x5 FILLER_202_1871 ();
 b15zdnd11an1n64x5 FILLER_202_1935 ();
 b15zdnd11an1n64x5 FILLER_202_1999 ();
 b15zdnd11an1n64x5 FILLER_202_2063 ();
 b15zdnd11an1n16x5 FILLER_202_2127 ();
 b15zdnd11an1n08x5 FILLER_202_2143 ();
 b15zdnd00an1n02x5 FILLER_202_2151 ();
 b15zdnd00an1n01x5 FILLER_202_2153 ();
 b15zdnd11an1n32x5 FILLER_202_2162 ();
 b15zdnd11an1n16x5 FILLER_202_2194 ();
 b15zdnd11an1n08x5 FILLER_202_2210 ();
 b15zdnd00an1n01x5 FILLER_202_2218 ();
 b15zdnd11an1n08x5 FILLER_202_2261 ();
 b15zdnd11an1n04x5 FILLER_202_2269 ();
 b15zdnd00an1n02x5 FILLER_202_2273 ();
 b15zdnd00an1n01x5 FILLER_202_2275 ();
 b15zdnd11an1n64x5 FILLER_203_0 ();
 b15zdnd11an1n64x5 FILLER_203_64 ();
 b15zdnd11an1n64x5 FILLER_203_128 ();
 b15zdnd11an1n64x5 FILLER_203_192 ();
 b15zdnd11an1n64x5 FILLER_203_256 ();
 b15zdnd11an1n64x5 FILLER_203_320 ();
 b15zdnd11an1n64x5 FILLER_203_384 ();
 b15zdnd11an1n64x5 FILLER_203_448 ();
 b15zdnd11an1n64x5 FILLER_203_512 ();
 b15zdnd11an1n64x5 FILLER_203_576 ();
 b15zdnd11an1n64x5 FILLER_203_640 ();
 b15zdnd11an1n64x5 FILLER_203_704 ();
 b15zdnd11an1n64x5 FILLER_203_768 ();
 b15zdnd11an1n64x5 FILLER_203_832 ();
 b15zdnd11an1n64x5 FILLER_203_896 ();
 b15zdnd11an1n64x5 FILLER_203_960 ();
 b15zdnd11an1n64x5 FILLER_203_1024 ();
 b15zdnd11an1n64x5 FILLER_203_1088 ();
 b15zdnd11an1n64x5 FILLER_203_1152 ();
 b15zdnd11an1n64x5 FILLER_203_1216 ();
 b15zdnd11an1n64x5 FILLER_203_1280 ();
 b15zdnd11an1n64x5 FILLER_203_1344 ();
 b15zdnd11an1n64x5 FILLER_203_1408 ();
 b15zdnd11an1n64x5 FILLER_203_1472 ();
 b15zdnd11an1n64x5 FILLER_203_1536 ();
 b15zdnd11an1n64x5 FILLER_203_1600 ();
 b15zdnd11an1n64x5 FILLER_203_1664 ();
 b15zdnd11an1n64x5 FILLER_203_1728 ();
 b15zdnd11an1n64x5 FILLER_203_1792 ();
 b15zdnd11an1n64x5 FILLER_203_1856 ();
 b15zdnd11an1n64x5 FILLER_203_1920 ();
 b15zdnd11an1n64x5 FILLER_203_1984 ();
 b15zdnd11an1n64x5 FILLER_203_2048 ();
 b15zdnd11an1n64x5 FILLER_203_2112 ();
 b15zdnd11an1n64x5 FILLER_203_2176 ();
 b15zdnd11an1n32x5 FILLER_203_2240 ();
 b15zdnd11an1n08x5 FILLER_203_2272 ();
 b15zdnd11an1n04x5 FILLER_203_2280 ();
 b15zdnd11an1n64x5 FILLER_204_8 ();
 b15zdnd11an1n64x5 FILLER_204_72 ();
 b15zdnd11an1n64x5 FILLER_204_136 ();
 b15zdnd11an1n64x5 FILLER_204_200 ();
 b15zdnd11an1n64x5 FILLER_204_264 ();
 b15zdnd11an1n64x5 FILLER_204_328 ();
 b15zdnd11an1n32x5 FILLER_204_392 ();
 b15zdnd11an1n08x5 FILLER_204_424 ();
 b15zdnd11an1n04x5 FILLER_204_432 ();
 b15zdnd00an1n02x5 FILLER_204_436 ();
 b15zdnd11an1n64x5 FILLER_204_456 ();
 b15zdnd11an1n64x5 FILLER_204_520 ();
 b15zdnd11an1n64x5 FILLER_204_584 ();
 b15zdnd11an1n64x5 FILLER_204_648 ();
 b15zdnd11an1n04x5 FILLER_204_712 ();
 b15zdnd00an1n02x5 FILLER_204_716 ();
 b15zdnd11an1n64x5 FILLER_204_726 ();
 b15zdnd11an1n64x5 FILLER_204_790 ();
 b15zdnd11an1n64x5 FILLER_204_854 ();
 b15zdnd11an1n64x5 FILLER_204_918 ();
 b15zdnd11an1n64x5 FILLER_204_982 ();
 b15zdnd11an1n64x5 FILLER_204_1046 ();
 b15zdnd11an1n64x5 FILLER_204_1110 ();
 b15zdnd11an1n32x5 FILLER_204_1174 ();
 b15zdnd11an1n16x5 FILLER_204_1206 ();
 b15zdnd11an1n04x5 FILLER_204_1222 ();
 b15zdnd00an1n01x5 FILLER_204_1226 ();
 b15zdnd11an1n64x5 FILLER_204_1269 ();
 b15zdnd11an1n64x5 FILLER_204_1333 ();
 b15zdnd11an1n64x5 FILLER_204_1397 ();
 b15zdnd11an1n64x5 FILLER_204_1461 ();
 b15zdnd11an1n64x5 FILLER_204_1525 ();
 b15zdnd11an1n64x5 FILLER_204_1589 ();
 b15zdnd11an1n64x5 FILLER_204_1653 ();
 b15zdnd11an1n64x5 FILLER_204_1717 ();
 b15zdnd11an1n64x5 FILLER_204_1781 ();
 b15zdnd11an1n64x5 FILLER_204_1845 ();
 b15zdnd11an1n64x5 FILLER_204_1909 ();
 b15zdnd11an1n64x5 FILLER_204_1973 ();
 b15zdnd11an1n64x5 FILLER_204_2037 ();
 b15zdnd11an1n32x5 FILLER_204_2101 ();
 b15zdnd11an1n16x5 FILLER_204_2133 ();
 b15zdnd11an1n04x5 FILLER_204_2149 ();
 b15zdnd00an1n01x5 FILLER_204_2153 ();
 b15zdnd11an1n32x5 FILLER_204_2162 ();
 b15zdnd11an1n04x5 FILLER_204_2194 ();
 b15zdnd00an1n01x5 FILLER_204_2198 ();
 b15zdnd11an1n32x5 FILLER_204_2241 ();
 b15zdnd00an1n02x5 FILLER_204_2273 ();
 b15zdnd00an1n01x5 FILLER_204_2275 ();
 b15zdnd11an1n64x5 FILLER_205_0 ();
 b15zdnd11an1n64x5 FILLER_205_64 ();
 b15zdnd11an1n64x5 FILLER_205_128 ();
 b15zdnd11an1n32x5 FILLER_205_192 ();
 b15zdnd11an1n16x5 FILLER_205_224 ();
 b15zdnd11an1n08x5 FILLER_205_240 ();
 b15zdnd00an1n01x5 FILLER_205_248 ();
 b15zdnd11an1n64x5 FILLER_205_257 ();
 b15zdnd11an1n64x5 FILLER_205_321 ();
 b15zdnd11an1n64x5 FILLER_205_385 ();
 b15zdnd11an1n64x5 FILLER_205_449 ();
 b15zdnd11an1n64x5 FILLER_205_513 ();
 b15zdnd11an1n64x5 FILLER_205_577 ();
 b15zdnd11an1n64x5 FILLER_205_641 ();
 b15zdnd11an1n64x5 FILLER_205_705 ();
 b15zdnd11an1n64x5 FILLER_205_769 ();
 b15zdnd11an1n64x5 FILLER_205_833 ();
 b15zdnd11an1n16x5 FILLER_205_897 ();
 b15zdnd11an1n04x5 FILLER_205_913 ();
 b15zdnd00an1n01x5 FILLER_205_917 ();
 b15zdnd11an1n64x5 FILLER_205_960 ();
 b15zdnd11an1n64x5 FILLER_205_1024 ();
 b15zdnd11an1n64x5 FILLER_205_1088 ();
 b15zdnd11an1n64x5 FILLER_205_1152 ();
 b15zdnd11an1n64x5 FILLER_205_1216 ();
 b15zdnd11an1n64x5 FILLER_205_1280 ();
 b15zdnd11an1n64x5 FILLER_205_1344 ();
 b15zdnd11an1n64x5 FILLER_205_1408 ();
 b15zdnd11an1n32x5 FILLER_205_1472 ();
 b15zdnd00an1n02x5 FILLER_205_1504 ();
 b15zdnd11an1n64x5 FILLER_205_1548 ();
 b15zdnd11an1n64x5 FILLER_205_1612 ();
 b15zdnd11an1n64x5 FILLER_205_1676 ();
 b15zdnd11an1n64x5 FILLER_205_1740 ();
 b15zdnd11an1n64x5 FILLER_205_1804 ();
 b15zdnd11an1n64x5 FILLER_205_1868 ();
 b15zdnd11an1n64x5 FILLER_205_1932 ();
 b15zdnd11an1n64x5 FILLER_205_1996 ();
 b15zdnd11an1n64x5 FILLER_205_2060 ();
 b15zdnd11an1n64x5 FILLER_205_2124 ();
 b15zdnd11an1n64x5 FILLER_205_2188 ();
 b15zdnd11an1n32x5 FILLER_205_2252 ();
 b15zdnd11an1n64x5 FILLER_206_8 ();
 b15zdnd11an1n64x5 FILLER_206_72 ();
 b15zdnd11an1n64x5 FILLER_206_136 ();
 b15zdnd11an1n16x5 FILLER_206_200 ();
 b15zdnd11an1n04x5 FILLER_206_216 ();
 b15zdnd00an1n01x5 FILLER_206_220 ();
 b15zdnd11an1n64x5 FILLER_206_263 ();
 b15zdnd11an1n64x5 FILLER_206_327 ();
 b15zdnd11an1n64x5 FILLER_206_391 ();
 b15zdnd11an1n64x5 FILLER_206_455 ();
 b15zdnd11an1n32x5 FILLER_206_519 ();
 b15zdnd11an1n16x5 FILLER_206_551 ();
 b15zdnd11an1n08x5 FILLER_206_567 ();
 b15zdnd11an1n04x5 FILLER_206_575 ();
 b15zdnd11an1n64x5 FILLER_206_621 ();
 b15zdnd11an1n32x5 FILLER_206_685 ();
 b15zdnd00an1n01x5 FILLER_206_717 ();
 b15zdnd11an1n64x5 FILLER_206_726 ();
 b15zdnd11an1n64x5 FILLER_206_790 ();
 b15zdnd11an1n64x5 FILLER_206_854 ();
 b15zdnd11an1n64x5 FILLER_206_918 ();
 b15zdnd11an1n64x5 FILLER_206_982 ();
 b15zdnd11an1n64x5 FILLER_206_1046 ();
 b15zdnd11an1n64x5 FILLER_206_1110 ();
 b15zdnd11an1n16x5 FILLER_206_1174 ();
 b15zdnd11an1n08x5 FILLER_206_1190 ();
 b15zdnd11an1n04x5 FILLER_206_1198 ();
 b15zdnd11an1n64x5 FILLER_206_1244 ();
 b15zdnd11an1n64x5 FILLER_206_1308 ();
 b15zdnd11an1n64x5 FILLER_206_1372 ();
 b15zdnd11an1n64x5 FILLER_206_1436 ();
 b15zdnd11an1n64x5 FILLER_206_1500 ();
 b15zdnd11an1n64x5 FILLER_206_1564 ();
 b15zdnd11an1n64x5 FILLER_206_1628 ();
 b15zdnd11an1n64x5 FILLER_206_1692 ();
 b15zdnd11an1n64x5 FILLER_206_1756 ();
 b15zdnd11an1n64x5 FILLER_206_1820 ();
 b15zdnd11an1n64x5 FILLER_206_1884 ();
 b15zdnd11an1n64x5 FILLER_206_1948 ();
 b15zdnd11an1n64x5 FILLER_206_2012 ();
 b15zdnd11an1n64x5 FILLER_206_2076 ();
 b15zdnd11an1n08x5 FILLER_206_2140 ();
 b15zdnd11an1n04x5 FILLER_206_2148 ();
 b15zdnd00an1n02x5 FILLER_206_2152 ();
 b15zdnd11an1n64x5 FILLER_206_2162 ();
 b15zdnd11an1n16x5 FILLER_206_2226 ();
 b15zdnd11an1n08x5 FILLER_206_2242 ();
 b15zdnd11an1n04x5 FILLER_206_2250 ();
 b15zdnd00an1n02x5 FILLER_206_2254 ();
 b15zdnd11an1n08x5 FILLER_206_2261 ();
 b15zdnd11an1n04x5 FILLER_206_2269 ();
 b15zdnd00an1n02x5 FILLER_206_2273 ();
 b15zdnd00an1n01x5 FILLER_206_2275 ();
 b15zdnd11an1n64x5 FILLER_207_0 ();
 b15zdnd11an1n64x5 FILLER_207_64 ();
 b15zdnd11an1n64x5 FILLER_207_128 ();
 b15zdnd11an1n64x5 FILLER_207_192 ();
 b15zdnd11an1n64x5 FILLER_207_256 ();
 b15zdnd11an1n64x5 FILLER_207_320 ();
 b15zdnd11an1n64x5 FILLER_207_384 ();
 b15zdnd11an1n64x5 FILLER_207_448 ();
 b15zdnd11an1n64x5 FILLER_207_512 ();
 b15zdnd11an1n64x5 FILLER_207_576 ();
 b15zdnd11an1n64x5 FILLER_207_640 ();
 b15zdnd11an1n64x5 FILLER_207_704 ();
 b15zdnd11an1n64x5 FILLER_207_768 ();
 b15zdnd11an1n64x5 FILLER_207_832 ();
 b15zdnd11an1n64x5 FILLER_207_896 ();
 b15zdnd11an1n64x5 FILLER_207_960 ();
 b15zdnd11an1n64x5 FILLER_207_1024 ();
 b15zdnd11an1n64x5 FILLER_207_1088 ();
 b15zdnd11an1n64x5 FILLER_207_1152 ();
 b15zdnd11an1n16x5 FILLER_207_1216 ();
 b15zdnd11an1n08x5 FILLER_207_1232 ();
 b15zdnd11an1n04x5 FILLER_207_1240 ();
 b15zdnd00an1n02x5 FILLER_207_1244 ();
 b15zdnd11an1n64x5 FILLER_207_1291 ();
 b15zdnd11an1n64x5 FILLER_207_1355 ();
 b15zdnd11an1n64x5 FILLER_207_1419 ();
 b15zdnd11an1n64x5 FILLER_207_1483 ();
 b15zdnd11an1n64x5 FILLER_207_1547 ();
 b15zdnd11an1n64x5 FILLER_207_1611 ();
 b15zdnd11an1n64x5 FILLER_207_1675 ();
 b15zdnd11an1n64x5 FILLER_207_1739 ();
 b15zdnd11an1n64x5 FILLER_207_1803 ();
 b15zdnd11an1n64x5 FILLER_207_1867 ();
 b15zdnd11an1n64x5 FILLER_207_1931 ();
 b15zdnd11an1n64x5 FILLER_207_1995 ();
 b15zdnd11an1n64x5 FILLER_207_2059 ();
 b15zdnd11an1n64x5 FILLER_207_2123 ();
 b15zdnd11an1n32x5 FILLER_207_2187 ();
 b15zdnd11an1n08x5 FILLER_207_2219 ();
 b15zdnd11an1n04x5 FILLER_207_2227 ();
 b15zdnd11an1n16x5 FILLER_207_2236 ();
 b15zdnd11an1n04x5 FILLER_207_2252 ();
 b15zdnd00an1n02x5 FILLER_207_2256 ();
 b15zdnd00an1n01x5 FILLER_207_2258 ();
 b15zdnd11an1n16x5 FILLER_207_2264 ();
 b15zdnd11an1n04x5 FILLER_207_2280 ();
 b15zdnd11an1n64x5 FILLER_208_8 ();
 b15zdnd11an1n64x5 FILLER_208_72 ();
 b15zdnd11an1n64x5 FILLER_208_136 ();
 b15zdnd11an1n64x5 FILLER_208_200 ();
 b15zdnd11an1n64x5 FILLER_208_264 ();
 b15zdnd11an1n64x5 FILLER_208_328 ();
 b15zdnd11an1n64x5 FILLER_208_392 ();
 b15zdnd11an1n64x5 FILLER_208_456 ();
 b15zdnd11an1n64x5 FILLER_208_520 ();
 b15zdnd11an1n64x5 FILLER_208_584 ();
 b15zdnd11an1n64x5 FILLER_208_648 ();
 b15zdnd11an1n04x5 FILLER_208_712 ();
 b15zdnd00an1n02x5 FILLER_208_716 ();
 b15zdnd11an1n64x5 FILLER_208_726 ();
 b15zdnd11an1n64x5 FILLER_208_790 ();
 b15zdnd11an1n64x5 FILLER_208_854 ();
 b15zdnd11an1n64x5 FILLER_208_918 ();
 b15zdnd11an1n64x5 FILLER_208_982 ();
 b15zdnd11an1n64x5 FILLER_208_1046 ();
 b15zdnd11an1n64x5 FILLER_208_1110 ();
 b15zdnd11an1n64x5 FILLER_208_1174 ();
 b15zdnd11an1n64x5 FILLER_208_1238 ();
 b15zdnd11an1n64x5 FILLER_208_1302 ();
 b15zdnd11an1n64x5 FILLER_208_1366 ();
 b15zdnd11an1n64x5 FILLER_208_1430 ();
 b15zdnd11an1n64x5 FILLER_208_1494 ();
 b15zdnd11an1n64x5 FILLER_208_1558 ();
 b15zdnd11an1n64x5 FILLER_208_1622 ();
 b15zdnd11an1n64x5 FILLER_208_1686 ();
 b15zdnd11an1n64x5 FILLER_208_1750 ();
 b15zdnd11an1n64x5 FILLER_208_1814 ();
 b15zdnd11an1n64x5 FILLER_208_1878 ();
 b15zdnd11an1n64x5 FILLER_208_1942 ();
 b15zdnd11an1n64x5 FILLER_208_2006 ();
 b15zdnd11an1n64x5 FILLER_208_2070 ();
 b15zdnd11an1n16x5 FILLER_208_2134 ();
 b15zdnd11an1n04x5 FILLER_208_2150 ();
 b15zdnd11an1n64x5 FILLER_208_2162 ();
 b15zdnd11an1n16x5 FILLER_208_2226 ();
 b15zdnd00an1n02x5 FILLER_208_2242 ();
 b15zdnd11an1n08x5 FILLER_208_2249 ();
 b15zdnd00an1n02x5 FILLER_208_2257 ();
 b15zdnd00an1n01x5 FILLER_208_2259 ();
 b15zdnd11an1n04x5 FILLER_208_2265 ();
 b15zdnd00an1n02x5 FILLER_208_2274 ();
 b15zdnd11an1n64x5 FILLER_209_0 ();
 b15zdnd11an1n64x5 FILLER_209_64 ();
 b15zdnd11an1n64x5 FILLER_209_128 ();
 b15zdnd11an1n64x5 FILLER_209_192 ();
 b15zdnd11an1n64x5 FILLER_209_256 ();
 b15zdnd11an1n64x5 FILLER_209_320 ();
 b15zdnd11an1n64x5 FILLER_209_384 ();
 b15zdnd11an1n64x5 FILLER_209_448 ();
 b15zdnd11an1n64x5 FILLER_209_512 ();
 b15zdnd11an1n64x5 FILLER_209_576 ();
 b15zdnd11an1n64x5 FILLER_209_640 ();
 b15zdnd11an1n64x5 FILLER_209_704 ();
 b15zdnd11an1n64x5 FILLER_209_768 ();
 b15zdnd11an1n64x5 FILLER_209_832 ();
 b15zdnd11an1n64x5 FILLER_209_896 ();
 b15zdnd11an1n64x5 FILLER_209_960 ();
 b15zdnd11an1n64x5 FILLER_209_1024 ();
 b15zdnd11an1n64x5 FILLER_209_1088 ();
 b15zdnd11an1n64x5 FILLER_209_1152 ();
 b15zdnd11an1n16x5 FILLER_209_1216 ();
 b15zdnd11an1n04x5 FILLER_209_1232 ();
 b15zdnd11an1n64x5 FILLER_209_1281 ();
 b15zdnd11an1n64x5 FILLER_209_1345 ();
 b15zdnd11an1n64x5 FILLER_209_1409 ();
 b15zdnd11an1n64x5 FILLER_209_1473 ();
 b15zdnd11an1n64x5 FILLER_209_1537 ();
 b15zdnd11an1n64x5 FILLER_209_1601 ();
 b15zdnd11an1n64x5 FILLER_209_1665 ();
 b15zdnd11an1n64x5 FILLER_209_1729 ();
 b15zdnd11an1n64x5 FILLER_209_1793 ();
 b15zdnd11an1n64x5 FILLER_209_1857 ();
 b15zdnd11an1n64x5 FILLER_209_1921 ();
 b15zdnd11an1n64x5 FILLER_209_1985 ();
 b15zdnd11an1n64x5 FILLER_209_2049 ();
 b15zdnd11an1n64x5 FILLER_209_2113 ();
 b15zdnd11an1n64x5 FILLER_209_2177 ();
 b15zdnd11an1n16x5 FILLER_209_2241 ();
 b15zdnd00an1n02x5 FILLER_209_2257 ();
 b15zdnd11an1n16x5 FILLER_209_2264 ();
 b15zdnd11an1n04x5 FILLER_209_2280 ();
 b15zdnd11an1n64x5 FILLER_210_8 ();
 b15zdnd11an1n64x5 FILLER_210_72 ();
 b15zdnd11an1n64x5 FILLER_210_136 ();
 b15zdnd11an1n64x5 FILLER_210_200 ();
 b15zdnd11an1n64x5 FILLER_210_264 ();
 b15zdnd11an1n64x5 FILLER_210_328 ();
 b15zdnd11an1n64x5 FILLER_210_392 ();
 b15zdnd11an1n64x5 FILLER_210_456 ();
 b15zdnd11an1n64x5 FILLER_210_520 ();
 b15zdnd11an1n64x5 FILLER_210_584 ();
 b15zdnd11an1n64x5 FILLER_210_648 ();
 b15zdnd11an1n04x5 FILLER_210_712 ();
 b15zdnd00an1n02x5 FILLER_210_716 ();
 b15zdnd11an1n64x5 FILLER_210_726 ();
 b15zdnd11an1n64x5 FILLER_210_790 ();
 b15zdnd11an1n64x5 FILLER_210_854 ();
 b15zdnd11an1n64x5 FILLER_210_918 ();
 b15zdnd11an1n64x5 FILLER_210_982 ();
 b15zdnd11an1n64x5 FILLER_210_1046 ();
 b15zdnd11an1n32x5 FILLER_210_1110 ();
 b15zdnd11an1n08x5 FILLER_210_1142 ();
 b15zdnd00an1n02x5 FILLER_210_1150 ();
 b15zdnd00an1n01x5 FILLER_210_1152 ();
 b15zdnd11an1n32x5 FILLER_210_1169 ();
 b15zdnd11an1n16x5 FILLER_210_1201 ();
 b15zdnd11an1n08x5 FILLER_210_1217 ();
 b15zdnd11an1n04x5 FILLER_210_1225 ();
 b15zdnd00an1n01x5 FILLER_210_1229 ();
 b15zdnd11an1n16x5 FILLER_210_1240 ();
 b15zdnd11an1n04x5 FILLER_210_1256 ();
 b15zdnd00an1n02x5 FILLER_210_1260 ();
 b15zdnd00an1n01x5 FILLER_210_1262 ();
 b15zdnd11an1n64x5 FILLER_210_1283 ();
 b15zdnd11an1n64x5 FILLER_210_1347 ();
 b15zdnd11an1n64x5 FILLER_210_1411 ();
 b15zdnd11an1n64x5 FILLER_210_1475 ();
 b15zdnd11an1n64x5 FILLER_210_1539 ();
 b15zdnd11an1n64x5 FILLER_210_1603 ();
 b15zdnd11an1n64x5 FILLER_210_1667 ();
 b15zdnd11an1n64x5 FILLER_210_1731 ();
 b15zdnd11an1n64x5 FILLER_210_1795 ();
 b15zdnd11an1n64x5 FILLER_210_1859 ();
 b15zdnd11an1n64x5 FILLER_210_1923 ();
 b15zdnd11an1n64x5 FILLER_210_1987 ();
 b15zdnd11an1n64x5 FILLER_210_2051 ();
 b15zdnd11an1n32x5 FILLER_210_2115 ();
 b15zdnd11an1n04x5 FILLER_210_2147 ();
 b15zdnd00an1n02x5 FILLER_210_2151 ();
 b15zdnd00an1n01x5 FILLER_210_2153 ();
 b15zdnd11an1n64x5 FILLER_210_2162 ();
 b15zdnd11an1n16x5 FILLER_210_2226 ();
 b15zdnd11an1n08x5 FILLER_210_2242 ();
 b15zdnd00an1n01x5 FILLER_210_2250 ();
 b15zdnd11an1n16x5 FILLER_210_2256 ();
 b15zdnd11an1n04x5 FILLER_210_2272 ();
 b15zdnd11an1n64x5 FILLER_211_0 ();
 b15zdnd11an1n64x5 FILLER_211_64 ();
 b15zdnd11an1n64x5 FILLER_211_128 ();
 b15zdnd11an1n64x5 FILLER_211_192 ();
 b15zdnd11an1n64x5 FILLER_211_256 ();
 b15zdnd11an1n64x5 FILLER_211_320 ();
 b15zdnd11an1n64x5 FILLER_211_384 ();
 b15zdnd11an1n64x5 FILLER_211_448 ();
 b15zdnd11an1n64x5 FILLER_211_512 ();
 b15zdnd11an1n64x5 FILLER_211_576 ();
 b15zdnd11an1n64x5 FILLER_211_640 ();
 b15zdnd11an1n64x5 FILLER_211_704 ();
 b15zdnd11an1n64x5 FILLER_211_768 ();
 b15zdnd11an1n64x5 FILLER_211_832 ();
 b15zdnd11an1n64x5 FILLER_211_896 ();
 b15zdnd11an1n64x5 FILLER_211_960 ();
 b15zdnd11an1n64x5 FILLER_211_1024 ();
 b15zdnd11an1n32x5 FILLER_211_1088 ();
 b15zdnd11an1n16x5 FILLER_211_1120 ();
 b15zdnd11an1n08x5 FILLER_211_1136 ();
 b15zdnd11an1n04x5 FILLER_211_1144 ();
 b15zdnd11an1n64x5 FILLER_211_1193 ();
 b15zdnd11an1n64x5 FILLER_211_1257 ();
 b15zdnd11an1n64x5 FILLER_211_1321 ();
 b15zdnd11an1n64x5 FILLER_211_1385 ();
 b15zdnd11an1n64x5 FILLER_211_1449 ();
 b15zdnd11an1n64x5 FILLER_211_1513 ();
 b15zdnd11an1n64x5 FILLER_211_1577 ();
 b15zdnd11an1n64x5 FILLER_211_1641 ();
 b15zdnd11an1n64x5 FILLER_211_1705 ();
 b15zdnd11an1n64x5 FILLER_211_1769 ();
 b15zdnd11an1n64x5 FILLER_211_1833 ();
 b15zdnd11an1n64x5 FILLER_211_1897 ();
 b15zdnd11an1n64x5 FILLER_211_1961 ();
 b15zdnd11an1n64x5 FILLER_211_2025 ();
 b15zdnd11an1n64x5 FILLER_211_2089 ();
 b15zdnd11an1n64x5 FILLER_211_2153 ();
 b15zdnd11an1n64x5 FILLER_211_2217 ();
 b15zdnd00an1n02x5 FILLER_211_2281 ();
 b15zdnd00an1n01x5 FILLER_211_2283 ();
 b15zdnd11an1n64x5 FILLER_212_8 ();
 b15zdnd11an1n64x5 FILLER_212_72 ();
 b15zdnd11an1n64x5 FILLER_212_136 ();
 b15zdnd11an1n64x5 FILLER_212_200 ();
 b15zdnd11an1n64x5 FILLER_212_264 ();
 b15zdnd11an1n64x5 FILLER_212_328 ();
 b15zdnd11an1n16x5 FILLER_212_392 ();
 b15zdnd11an1n08x5 FILLER_212_408 ();
 b15zdnd00an1n01x5 FILLER_212_416 ();
 b15zdnd11an1n64x5 FILLER_212_428 ();
 b15zdnd11an1n64x5 FILLER_212_492 ();
 b15zdnd11an1n64x5 FILLER_212_556 ();
 b15zdnd11an1n64x5 FILLER_212_620 ();
 b15zdnd11an1n32x5 FILLER_212_684 ();
 b15zdnd00an1n02x5 FILLER_212_716 ();
 b15zdnd11an1n64x5 FILLER_212_726 ();
 b15zdnd11an1n64x5 FILLER_212_790 ();
 b15zdnd11an1n64x5 FILLER_212_854 ();
 b15zdnd11an1n64x5 FILLER_212_918 ();
 b15zdnd11an1n64x5 FILLER_212_982 ();
 b15zdnd11an1n64x5 FILLER_212_1046 ();
 b15zdnd11an1n16x5 FILLER_212_1110 ();
 b15zdnd11an1n04x5 FILLER_212_1126 ();
 b15zdnd00an1n02x5 FILLER_212_1130 ();
 b15zdnd11an1n64x5 FILLER_212_1177 ();
 b15zdnd11an1n64x5 FILLER_212_1241 ();
 b15zdnd11an1n64x5 FILLER_212_1305 ();
 b15zdnd11an1n64x5 FILLER_212_1369 ();
 b15zdnd11an1n64x5 FILLER_212_1433 ();
 b15zdnd11an1n64x5 FILLER_212_1497 ();
 b15zdnd11an1n64x5 FILLER_212_1561 ();
 b15zdnd11an1n64x5 FILLER_212_1625 ();
 b15zdnd11an1n64x5 FILLER_212_1689 ();
 b15zdnd11an1n64x5 FILLER_212_1753 ();
 b15zdnd11an1n64x5 FILLER_212_1817 ();
 b15zdnd11an1n64x5 FILLER_212_1881 ();
 b15zdnd11an1n64x5 FILLER_212_1945 ();
 b15zdnd11an1n64x5 FILLER_212_2009 ();
 b15zdnd11an1n64x5 FILLER_212_2073 ();
 b15zdnd11an1n16x5 FILLER_212_2137 ();
 b15zdnd00an1n01x5 FILLER_212_2153 ();
 b15zdnd11an1n64x5 FILLER_212_2162 ();
 b15zdnd11an1n32x5 FILLER_212_2226 ();
 b15zdnd11an1n16x5 FILLER_212_2258 ();
 b15zdnd00an1n02x5 FILLER_212_2274 ();
 b15zdnd11an1n64x5 FILLER_213_0 ();
 b15zdnd11an1n64x5 FILLER_213_64 ();
 b15zdnd11an1n64x5 FILLER_213_128 ();
 b15zdnd11an1n64x5 FILLER_213_192 ();
 b15zdnd11an1n64x5 FILLER_213_256 ();
 b15zdnd11an1n64x5 FILLER_213_320 ();
 b15zdnd11an1n32x5 FILLER_213_388 ();
 b15zdnd11an1n16x5 FILLER_213_420 ();
 b15zdnd00an1n01x5 FILLER_213_436 ();
 b15zdnd11an1n64x5 FILLER_213_441 ();
 b15zdnd11an1n64x5 FILLER_213_505 ();
 b15zdnd11an1n64x5 FILLER_213_569 ();
 b15zdnd11an1n64x5 FILLER_213_633 ();
 b15zdnd11an1n64x5 FILLER_213_697 ();
 b15zdnd11an1n64x5 FILLER_213_761 ();
 b15zdnd11an1n64x5 FILLER_213_825 ();
 b15zdnd11an1n64x5 FILLER_213_889 ();
 b15zdnd11an1n64x5 FILLER_213_953 ();
 b15zdnd11an1n64x5 FILLER_213_1017 ();
 b15zdnd11an1n32x5 FILLER_213_1081 ();
 b15zdnd11an1n16x5 FILLER_213_1113 ();
 b15zdnd11an1n08x5 FILLER_213_1129 ();
 b15zdnd11an1n04x5 FILLER_213_1137 ();
 b15zdnd00an1n02x5 FILLER_213_1141 ();
 b15zdnd11an1n64x5 FILLER_213_1155 ();
 b15zdnd11an1n64x5 FILLER_213_1219 ();
 b15zdnd11an1n16x5 FILLER_213_1283 ();
 b15zdnd11an1n08x5 FILLER_213_1299 ();
 b15zdnd11an1n04x5 FILLER_213_1307 ();
 b15zdnd00an1n01x5 FILLER_213_1311 ();
 b15zdnd11an1n64x5 FILLER_213_1335 ();
 b15zdnd11an1n04x5 FILLER_213_1399 ();
 b15zdnd11an1n64x5 FILLER_213_1414 ();
 b15zdnd11an1n64x5 FILLER_213_1478 ();
 b15zdnd11an1n64x5 FILLER_213_1542 ();
 b15zdnd11an1n64x5 FILLER_213_1606 ();
 b15zdnd11an1n64x5 FILLER_213_1670 ();
 b15zdnd11an1n64x5 FILLER_213_1734 ();
 b15zdnd11an1n64x5 FILLER_213_1798 ();
 b15zdnd11an1n64x5 FILLER_213_1862 ();
 b15zdnd11an1n64x5 FILLER_213_1926 ();
 b15zdnd11an1n64x5 FILLER_213_1990 ();
 b15zdnd11an1n64x5 FILLER_213_2054 ();
 b15zdnd11an1n64x5 FILLER_213_2118 ();
 b15zdnd11an1n64x5 FILLER_213_2182 ();
 b15zdnd11an1n32x5 FILLER_213_2246 ();
 b15zdnd11an1n04x5 FILLER_213_2278 ();
 b15zdnd00an1n02x5 FILLER_213_2282 ();
 b15zdnd11an1n64x5 FILLER_214_8 ();
 b15zdnd11an1n64x5 FILLER_214_72 ();
 b15zdnd11an1n64x5 FILLER_214_136 ();
 b15zdnd11an1n64x5 FILLER_214_200 ();
 b15zdnd11an1n64x5 FILLER_214_264 ();
 b15zdnd11an1n64x5 FILLER_214_328 ();
 b15zdnd11an1n32x5 FILLER_214_392 ();
 b15zdnd00an1n02x5 FILLER_214_424 ();
 b15zdnd00an1n01x5 FILLER_214_426 ();
 b15zdnd11an1n64x5 FILLER_214_448 ();
 b15zdnd11an1n64x5 FILLER_214_512 ();
 b15zdnd11an1n64x5 FILLER_214_576 ();
 b15zdnd11an1n64x5 FILLER_214_640 ();
 b15zdnd11an1n08x5 FILLER_214_704 ();
 b15zdnd11an1n04x5 FILLER_214_712 ();
 b15zdnd00an1n02x5 FILLER_214_716 ();
 b15zdnd11an1n64x5 FILLER_214_726 ();
 b15zdnd11an1n64x5 FILLER_214_790 ();
 b15zdnd11an1n64x5 FILLER_214_854 ();
 b15zdnd11an1n64x5 FILLER_214_918 ();
 b15zdnd11an1n64x5 FILLER_214_982 ();
 b15zdnd11an1n64x5 FILLER_214_1046 ();
 b15zdnd11an1n16x5 FILLER_214_1110 ();
 b15zdnd00an1n01x5 FILLER_214_1126 ();
 b15zdnd11an1n64x5 FILLER_214_1159 ();
 b15zdnd00an1n01x5 FILLER_214_1223 ();
 b15zdnd11an1n64x5 FILLER_214_1235 ();
 b15zdnd11an1n64x5 FILLER_214_1299 ();
 b15zdnd11an1n32x5 FILLER_214_1363 ();
 b15zdnd11an1n04x5 FILLER_214_1437 ();
 b15zdnd11an1n08x5 FILLER_214_1447 ();
 b15zdnd11an1n64x5 FILLER_214_1471 ();
 b15zdnd11an1n64x5 FILLER_214_1535 ();
 b15zdnd11an1n64x5 FILLER_214_1599 ();
 b15zdnd11an1n64x5 FILLER_214_1663 ();
 b15zdnd11an1n64x5 FILLER_214_1727 ();
 b15zdnd11an1n64x5 FILLER_214_1791 ();
 b15zdnd11an1n64x5 FILLER_214_1855 ();
 b15zdnd11an1n64x5 FILLER_214_1919 ();
 b15zdnd11an1n64x5 FILLER_214_1983 ();
 b15zdnd11an1n64x5 FILLER_214_2047 ();
 b15zdnd11an1n32x5 FILLER_214_2111 ();
 b15zdnd11an1n08x5 FILLER_214_2143 ();
 b15zdnd00an1n02x5 FILLER_214_2151 ();
 b15zdnd00an1n01x5 FILLER_214_2153 ();
 b15zdnd11an1n64x5 FILLER_214_2162 ();
 b15zdnd11an1n32x5 FILLER_214_2226 ();
 b15zdnd11an1n16x5 FILLER_214_2258 ();
 b15zdnd00an1n02x5 FILLER_214_2274 ();
 b15zdnd11an1n64x5 FILLER_215_0 ();
 b15zdnd11an1n64x5 FILLER_215_64 ();
 b15zdnd11an1n64x5 FILLER_215_128 ();
 b15zdnd11an1n64x5 FILLER_215_192 ();
 b15zdnd11an1n64x5 FILLER_215_256 ();
 b15zdnd11an1n64x5 FILLER_215_320 ();
 b15zdnd11an1n64x5 FILLER_215_384 ();
 b15zdnd11an1n64x5 FILLER_215_448 ();
 b15zdnd11an1n64x5 FILLER_215_512 ();
 b15zdnd11an1n64x5 FILLER_215_576 ();
 b15zdnd11an1n32x5 FILLER_215_640 ();
 b15zdnd11an1n16x5 FILLER_215_672 ();
 b15zdnd11an1n08x5 FILLER_215_688 ();
 b15zdnd11an1n04x5 FILLER_215_696 ();
 b15zdnd00an1n02x5 FILLER_215_700 ();
 b15zdnd11an1n64x5 FILLER_215_744 ();
 b15zdnd11an1n64x5 FILLER_215_808 ();
 b15zdnd11an1n64x5 FILLER_215_872 ();
 b15zdnd11an1n64x5 FILLER_215_936 ();
 b15zdnd11an1n64x5 FILLER_215_1000 ();
 b15zdnd11an1n64x5 FILLER_215_1064 ();
 b15zdnd11an1n64x5 FILLER_215_1128 ();
 b15zdnd11an1n64x5 FILLER_215_1192 ();
 b15zdnd11an1n64x5 FILLER_215_1256 ();
 b15zdnd11an1n32x5 FILLER_215_1320 ();
 b15zdnd11an1n04x5 FILLER_215_1352 ();
 b15zdnd00an1n01x5 FILLER_215_1356 ();
 b15zdnd11an1n64x5 FILLER_215_1373 ();
 b15zdnd11an1n64x5 FILLER_215_1437 ();
 b15zdnd11an1n64x5 FILLER_215_1501 ();
 b15zdnd11an1n64x5 FILLER_215_1565 ();
 b15zdnd11an1n64x5 FILLER_215_1629 ();
 b15zdnd11an1n16x5 FILLER_215_1693 ();
 b15zdnd11an1n08x5 FILLER_215_1709 ();
 b15zdnd00an1n02x5 FILLER_215_1717 ();
 b15zdnd11an1n64x5 FILLER_215_1761 ();
 b15zdnd11an1n64x5 FILLER_215_1825 ();
 b15zdnd11an1n64x5 FILLER_215_1889 ();
 b15zdnd11an1n64x5 FILLER_215_1953 ();
 b15zdnd11an1n64x5 FILLER_215_2017 ();
 b15zdnd11an1n64x5 FILLER_215_2081 ();
 b15zdnd11an1n64x5 FILLER_215_2145 ();
 b15zdnd11an1n64x5 FILLER_215_2209 ();
 b15zdnd11an1n08x5 FILLER_215_2273 ();
 b15zdnd00an1n02x5 FILLER_215_2281 ();
 b15zdnd00an1n01x5 FILLER_215_2283 ();
 b15zdnd11an1n64x5 FILLER_216_8 ();
 b15zdnd11an1n64x5 FILLER_216_72 ();
 b15zdnd11an1n64x5 FILLER_216_136 ();
 b15zdnd11an1n64x5 FILLER_216_200 ();
 b15zdnd11an1n64x5 FILLER_216_264 ();
 b15zdnd11an1n64x5 FILLER_216_328 ();
 b15zdnd11an1n64x5 FILLER_216_392 ();
 b15zdnd11an1n64x5 FILLER_216_456 ();
 b15zdnd11an1n64x5 FILLER_216_520 ();
 b15zdnd11an1n64x5 FILLER_216_584 ();
 b15zdnd11an1n64x5 FILLER_216_648 ();
 b15zdnd11an1n04x5 FILLER_216_712 ();
 b15zdnd00an1n02x5 FILLER_216_716 ();
 b15zdnd11an1n64x5 FILLER_216_726 ();
 b15zdnd11an1n64x5 FILLER_216_790 ();
 b15zdnd11an1n64x5 FILLER_216_854 ();
 b15zdnd11an1n32x5 FILLER_216_918 ();
 b15zdnd11an1n16x5 FILLER_216_950 ();
 b15zdnd00an1n02x5 FILLER_216_966 ();
 b15zdnd00an1n01x5 FILLER_216_968 ();
 b15zdnd11an1n04x5 FILLER_216_973 ();
 b15zdnd11an1n64x5 FILLER_216_988 ();
 b15zdnd11an1n64x5 FILLER_216_1052 ();
 b15zdnd11an1n64x5 FILLER_216_1116 ();
 b15zdnd11an1n64x5 FILLER_216_1180 ();
 b15zdnd11an1n64x5 FILLER_216_1244 ();
 b15zdnd11an1n64x5 FILLER_216_1308 ();
 b15zdnd11an1n32x5 FILLER_216_1372 ();
 b15zdnd11an1n08x5 FILLER_216_1404 ();
 b15zdnd00an1n02x5 FILLER_216_1412 ();
 b15zdnd00an1n01x5 FILLER_216_1414 ();
 b15zdnd11an1n64x5 FILLER_216_1431 ();
 b15zdnd11an1n64x5 FILLER_216_1495 ();
 b15zdnd11an1n64x5 FILLER_216_1559 ();
 b15zdnd11an1n32x5 FILLER_216_1623 ();
 b15zdnd11an1n08x5 FILLER_216_1655 ();
 b15zdnd11an1n08x5 FILLER_216_1705 ();
 b15zdnd00an1n02x5 FILLER_216_1713 ();
 b15zdnd00an1n01x5 FILLER_216_1715 ();
 b15zdnd11an1n64x5 FILLER_216_1758 ();
 b15zdnd11an1n64x5 FILLER_216_1822 ();
 b15zdnd11an1n64x5 FILLER_216_1886 ();
 b15zdnd11an1n64x5 FILLER_216_1950 ();
 b15zdnd11an1n64x5 FILLER_216_2014 ();
 b15zdnd11an1n64x5 FILLER_216_2078 ();
 b15zdnd11an1n08x5 FILLER_216_2142 ();
 b15zdnd11an1n04x5 FILLER_216_2150 ();
 b15zdnd11an1n64x5 FILLER_216_2162 ();
 b15zdnd11an1n32x5 FILLER_216_2226 ();
 b15zdnd11an1n16x5 FILLER_216_2258 ();
 b15zdnd00an1n02x5 FILLER_216_2274 ();
 b15zdnd11an1n64x5 FILLER_217_0 ();
 b15zdnd11an1n64x5 FILLER_217_64 ();
 b15zdnd11an1n64x5 FILLER_217_128 ();
 b15zdnd11an1n64x5 FILLER_217_192 ();
 b15zdnd11an1n64x5 FILLER_217_256 ();
 b15zdnd11an1n64x5 FILLER_217_320 ();
 b15zdnd11an1n08x5 FILLER_217_384 ();
 b15zdnd00an1n01x5 FILLER_217_392 ();
 b15zdnd11an1n64x5 FILLER_217_425 ();
 b15zdnd11an1n64x5 FILLER_217_489 ();
 b15zdnd11an1n64x5 FILLER_217_553 ();
 b15zdnd11an1n64x5 FILLER_217_617 ();
 b15zdnd11an1n64x5 FILLER_217_681 ();
 b15zdnd11an1n64x5 FILLER_217_745 ();
 b15zdnd11an1n64x5 FILLER_217_809 ();
 b15zdnd11an1n64x5 FILLER_217_873 ();
 b15zdnd11an1n16x5 FILLER_217_937 ();
 b15zdnd11an1n08x5 FILLER_217_953 ();
 b15zdnd11an1n64x5 FILLER_217_992 ();
 b15zdnd11an1n64x5 FILLER_217_1056 ();
 b15zdnd11an1n64x5 FILLER_217_1120 ();
 b15zdnd11an1n64x5 FILLER_217_1184 ();
 b15zdnd11an1n64x5 FILLER_217_1248 ();
 b15zdnd11an1n64x5 FILLER_217_1312 ();
 b15zdnd11an1n64x5 FILLER_217_1376 ();
 b15zdnd11an1n64x5 FILLER_217_1440 ();
 b15zdnd11an1n64x5 FILLER_217_1504 ();
 b15zdnd11an1n64x5 FILLER_217_1568 ();
 b15zdnd11an1n64x5 FILLER_217_1632 ();
 b15zdnd11an1n64x5 FILLER_217_1696 ();
 b15zdnd11an1n64x5 FILLER_217_1760 ();
 b15zdnd11an1n64x5 FILLER_217_1824 ();
 b15zdnd11an1n64x5 FILLER_217_1888 ();
 b15zdnd11an1n64x5 FILLER_217_1952 ();
 b15zdnd11an1n64x5 FILLER_217_2016 ();
 b15zdnd11an1n64x5 FILLER_217_2080 ();
 b15zdnd11an1n64x5 FILLER_217_2144 ();
 b15zdnd11an1n32x5 FILLER_217_2208 ();
 b15zdnd11an1n08x5 FILLER_217_2240 ();
 b15zdnd11an1n04x5 FILLER_217_2248 ();
 b15zdnd00an1n02x5 FILLER_217_2252 ();
 b15zdnd11an1n08x5 FILLER_217_2258 ();
 b15zdnd00an1n02x5 FILLER_217_2266 ();
 b15zdnd11an1n08x5 FILLER_217_2272 ();
 b15zdnd11an1n04x5 FILLER_217_2280 ();
 b15zdnd11an1n64x5 FILLER_218_8 ();
 b15zdnd11an1n64x5 FILLER_218_72 ();
 b15zdnd11an1n64x5 FILLER_218_136 ();
 b15zdnd11an1n64x5 FILLER_218_200 ();
 b15zdnd11an1n64x5 FILLER_218_264 ();
 b15zdnd11an1n64x5 FILLER_218_328 ();
 b15zdnd11an1n32x5 FILLER_218_392 ();
 b15zdnd11an1n16x5 FILLER_218_424 ();
 b15zdnd11an1n08x5 FILLER_218_440 ();
 b15zdnd11an1n04x5 FILLER_218_448 ();
 b15zdnd00an1n02x5 FILLER_218_452 ();
 b15zdnd11an1n32x5 FILLER_218_472 ();
 b15zdnd11an1n16x5 FILLER_218_504 ();
 b15zdnd11an1n08x5 FILLER_218_520 ();
 b15zdnd00an1n02x5 FILLER_218_528 ();
 b15zdnd00an1n01x5 FILLER_218_530 ();
 b15zdnd11an1n64x5 FILLER_218_573 ();
 b15zdnd11an1n64x5 FILLER_218_637 ();
 b15zdnd11an1n16x5 FILLER_218_701 ();
 b15zdnd00an1n01x5 FILLER_218_717 ();
 b15zdnd11an1n64x5 FILLER_218_726 ();
 b15zdnd11an1n64x5 FILLER_218_790 ();
 b15zdnd11an1n64x5 FILLER_218_854 ();
 b15zdnd11an1n64x5 FILLER_218_918 ();
 b15zdnd11an1n64x5 FILLER_218_982 ();
 b15zdnd11an1n64x5 FILLER_218_1046 ();
 b15zdnd11an1n64x5 FILLER_218_1110 ();
 b15zdnd11an1n64x5 FILLER_218_1174 ();
 b15zdnd11an1n64x5 FILLER_218_1238 ();
 b15zdnd11an1n64x5 FILLER_218_1302 ();
 b15zdnd11an1n64x5 FILLER_218_1366 ();
 b15zdnd11an1n64x5 FILLER_218_1430 ();
 b15zdnd11an1n64x5 FILLER_218_1494 ();
 b15zdnd11an1n64x5 FILLER_218_1558 ();
 b15zdnd11an1n32x5 FILLER_218_1622 ();
 b15zdnd11an1n64x5 FILLER_218_1696 ();
 b15zdnd11an1n64x5 FILLER_218_1760 ();
 b15zdnd11an1n64x5 FILLER_218_1824 ();
 b15zdnd11an1n64x5 FILLER_218_1888 ();
 b15zdnd11an1n64x5 FILLER_218_1952 ();
 b15zdnd11an1n64x5 FILLER_218_2016 ();
 b15zdnd11an1n32x5 FILLER_218_2080 ();
 b15zdnd00an1n02x5 FILLER_218_2112 ();
 b15zdnd11an1n16x5 FILLER_218_2126 ();
 b15zdnd11an1n08x5 FILLER_218_2142 ();
 b15zdnd11an1n04x5 FILLER_218_2150 ();
 b15zdnd11an1n64x5 FILLER_218_2162 ();
 b15zdnd11an1n04x5 FILLER_218_2226 ();
 b15zdnd00an1n02x5 FILLER_218_2230 ();
 b15zdnd00an1n02x5 FILLER_218_2274 ();
 b15zdnd11an1n16x5 FILLER_219_0 ();
 b15zdnd11an1n08x5 FILLER_219_16 ();
 b15zdnd11an1n04x5 FILLER_219_24 ();
 b15zdnd00an1n02x5 FILLER_219_28 ();
 b15zdnd11an1n64x5 FILLER_219_40 ();
 b15zdnd11an1n64x5 FILLER_219_104 ();
 b15zdnd11an1n64x5 FILLER_219_168 ();
 b15zdnd11an1n64x5 FILLER_219_232 ();
 b15zdnd11an1n64x5 FILLER_219_296 ();
 b15zdnd11an1n64x5 FILLER_219_360 ();
 b15zdnd11an1n16x5 FILLER_219_424 ();
 b15zdnd11an1n08x5 FILLER_219_440 ();
 b15zdnd11an1n04x5 FILLER_219_448 ();
 b15zdnd00an1n02x5 FILLER_219_452 ();
 b15zdnd11an1n64x5 FILLER_219_496 ();
 b15zdnd11an1n64x5 FILLER_219_560 ();
 b15zdnd11an1n64x5 FILLER_219_624 ();
 b15zdnd11an1n64x5 FILLER_219_688 ();
 b15zdnd11an1n64x5 FILLER_219_752 ();
 b15zdnd11an1n64x5 FILLER_219_816 ();
 b15zdnd11an1n64x5 FILLER_219_880 ();
 b15zdnd11an1n08x5 FILLER_219_944 ();
 b15zdnd11an1n04x5 FILLER_219_952 ();
 b15zdnd00an1n02x5 FILLER_219_956 ();
 b15zdnd00an1n01x5 FILLER_219_958 ();
 b15zdnd11an1n04x5 FILLER_219_965 ();
 b15zdnd11an1n08x5 FILLER_219_987 ();
 b15zdnd11an1n04x5 FILLER_219_995 ();
 b15zdnd00an1n01x5 FILLER_219_999 ();
 b15zdnd11an1n64x5 FILLER_219_1012 ();
 b15zdnd11an1n64x5 FILLER_219_1076 ();
 b15zdnd11an1n64x5 FILLER_219_1140 ();
 b15zdnd11an1n64x5 FILLER_219_1204 ();
 b15zdnd11an1n64x5 FILLER_219_1268 ();
 b15zdnd11an1n64x5 FILLER_219_1332 ();
 b15zdnd11an1n64x5 FILLER_219_1396 ();
 b15zdnd11an1n64x5 FILLER_219_1460 ();
 b15zdnd11an1n64x5 FILLER_219_1524 ();
 b15zdnd11an1n64x5 FILLER_219_1588 ();
 b15zdnd11an1n64x5 FILLER_219_1652 ();
 b15zdnd11an1n64x5 FILLER_219_1716 ();
 b15zdnd11an1n64x5 FILLER_219_1780 ();
 b15zdnd11an1n64x5 FILLER_219_1844 ();
 b15zdnd11an1n64x5 FILLER_219_1908 ();
 b15zdnd11an1n64x5 FILLER_219_1972 ();
 b15zdnd11an1n16x5 FILLER_219_2036 ();
 b15zdnd11an1n04x5 FILLER_219_2052 ();
 b15zdnd00an1n02x5 FILLER_219_2056 ();
 b15zdnd00an1n01x5 FILLER_219_2058 ();
 b15zdnd11an1n08x5 FILLER_219_2071 ();
 b15zdnd11an1n32x5 FILLER_219_2095 ();
 b15zdnd11an1n16x5 FILLER_219_2127 ();
 b15zdnd11an1n08x5 FILLER_219_2143 ();
 b15zdnd11an1n04x5 FILLER_219_2151 ();
 b15zdnd00an1n02x5 FILLER_219_2155 ();
 b15zdnd11an1n64x5 FILLER_219_2173 ();
 b15zdnd11an1n32x5 FILLER_219_2237 ();
 b15zdnd11an1n08x5 FILLER_219_2269 ();
 b15zdnd11an1n04x5 FILLER_219_2277 ();
 b15zdnd00an1n02x5 FILLER_219_2281 ();
 b15zdnd00an1n01x5 FILLER_219_2283 ();
 b15zdnd11an1n16x5 FILLER_220_8 ();
 b15zdnd11an1n04x5 FILLER_220_24 ();
 b15zdnd00an1n02x5 FILLER_220_28 ();
 b15zdnd00an1n01x5 FILLER_220_30 ();
 b15zdnd11an1n64x5 FILLER_220_51 ();
 b15zdnd11an1n64x5 FILLER_220_115 ();
 b15zdnd11an1n64x5 FILLER_220_179 ();
 b15zdnd11an1n64x5 FILLER_220_243 ();
 b15zdnd11an1n64x5 FILLER_220_307 ();
 b15zdnd11an1n64x5 FILLER_220_371 ();
 b15zdnd11an1n64x5 FILLER_220_435 ();
 b15zdnd11an1n32x5 FILLER_220_499 ();
 b15zdnd11an1n08x5 FILLER_220_531 ();
 b15zdnd00an1n01x5 FILLER_220_539 ();
 b15zdnd11an1n64x5 FILLER_220_582 ();
 b15zdnd11an1n64x5 FILLER_220_646 ();
 b15zdnd11an1n08x5 FILLER_220_710 ();
 b15zdnd11an1n64x5 FILLER_220_726 ();
 b15zdnd11an1n64x5 FILLER_220_790 ();
 b15zdnd11an1n64x5 FILLER_220_854 ();
 b15zdnd11an1n32x5 FILLER_220_918 ();
 b15zdnd11an1n04x5 FILLER_220_950 ();
 b15zdnd00an1n01x5 FILLER_220_954 ();
 b15zdnd11an1n64x5 FILLER_220_968 ();
 b15zdnd11an1n64x5 FILLER_220_1032 ();
 b15zdnd11an1n64x5 FILLER_220_1096 ();
 b15zdnd11an1n64x5 FILLER_220_1160 ();
 b15zdnd11an1n64x5 FILLER_220_1224 ();
 b15zdnd11an1n64x5 FILLER_220_1288 ();
 b15zdnd11an1n64x5 FILLER_220_1352 ();
 b15zdnd11an1n64x5 FILLER_220_1416 ();
 b15zdnd11an1n64x5 FILLER_220_1480 ();
 b15zdnd11an1n64x5 FILLER_220_1544 ();
 b15zdnd11an1n64x5 FILLER_220_1608 ();
 b15zdnd11an1n64x5 FILLER_220_1672 ();
 b15zdnd11an1n64x5 FILLER_220_1736 ();
 b15zdnd11an1n64x5 FILLER_220_1800 ();
 b15zdnd11an1n64x5 FILLER_220_1864 ();
 b15zdnd11an1n64x5 FILLER_220_1928 ();
 b15zdnd11an1n32x5 FILLER_220_1992 ();
 b15zdnd11an1n08x5 FILLER_220_2024 ();
 b15zdnd00an1n01x5 FILLER_220_2032 ();
 b15zdnd11an1n64x5 FILLER_220_2045 ();
 b15zdnd11an1n32x5 FILLER_220_2109 ();
 b15zdnd11an1n04x5 FILLER_220_2141 ();
 b15zdnd00an1n02x5 FILLER_220_2145 ();
 b15zdnd00an1n01x5 FILLER_220_2147 ();
 b15zdnd00an1n02x5 FILLER_220_2152 ();
 b15zdnd11an1n04x5 FILLER_220_2162 ();
 b15zdnd00an1n02x5 FILLER_220_2166 ();
 b15zdnd00an1n01x5 FILLER_220_2168 ();
 b15zdnd11an1n64x5 FILLER_220_2185 ();
 b15zdnd11an1n16x5 FILLER_220_2249 ();
 b15zdnd11an1n08x5 FILLER_220_2265 ();
 b15zdnd00an1n02x5 FILLER_220_2273 ();
 b15zdnd00an1n01x5 FILLER_220_2275 ();
 b15zdnd11an1n64x5 FILLER_221_0 ();
 b15zdnd11an1n64x5 FILLER_221_64 ();
 b15zdnd11an1n64x5 FILLER_221_128 ();
 b15zdnd11an1n64x5 FILLER_221_192 ();
 b15zdnd11an1n64x5 FILLER_221_256 ();
 b15zdnd11an1n64x5 FILLER_221_320 ();
 b15zdnd11an1n64x5 FILLER_221_384 ();
 b15zdnd11an1n16x5 FILLER_221_448 ();
 b15zdnd11an1n08x5 FILLER_221_464 ();
 b15zdnd11an1n04x5 FILLER_221_472 ();
 b15zdnd11an1n64x5 FILLER_221_484 ();
 b15zdnd11an1n64x5 FILLER_221_548 ();
 b15zdnd11an1n08x5 FILLER_221_612 ();
 b15zdnd11an1n04x5 FILLER_221_620 ();
 b15zdnd00an1n02x5 FILLER_221_624 ();
 b15zdnd11an1n64x5 FILLER_221_668 ();
 b15zdnd11an1n64x5 FILLER_221_732 ();
 b15zdnd11an1n64x5 FILLER_221_796 ();
 b15zdnd11an1n64x5 FILLER_221_860 ();
 b15zdnd11an1n32x5 FILLER_221_924 ();
 b15zdnd00an1n02x5 FILLER_221_956 ();
 b15zdnd00an1n01x5 FILLER_221_958 ();
 b15zdnd11an1n64x5 FILLER_221_972 ();
 b15zdnd11an1n16x5 FILLER_221_1036 ();
 b15zdnd11an1n08x5 FILLER_221_1052 ();
 b15zdnd11an1n04x5 FILLER_221_1060 ();
 b15zdnd11an1n64x5 FILLER_221_1087 ();
 b15zdnd11an1n64x5 FILLER_221_1151 ();
 b15zdnd11an1n32x5 FILLER_221_1215 ();
 b15zdnd11an1n08x5 FILLER_221_1247 ();
 b15zdnd00an1n02x5 FILLER_221_1255 ();
 b15zdnd11an1n64x5 FILLER_221_1299 ();
 b15zdnd11an1n64x5 FILLER_221_1363 ();
 b15zdnd11an1n64x5 FILLER_221_1443 ();
 b15zdnd11an1n64x5 FILLER_221_1507 ();
 b15zdnd11an1n64x5 FILLER_221_1571 ();
 b15zdnd11an1n64x5 FILLER_221_1635 ();
 b15zdnd11an1n64x5 FILLER_221_1699 ();
 b15zdnd11an1n64x5 FILLER_221_1763 ();
 b15zdnd11an1n64x5 FILLER_221_1827 ();
 b15zdnd11an1n64x5 FILLER_221_1891 ();
 b15zdnd11an1n64x5 FILLER_221_1955 ();
 b15zdnd11an1n64x5 FILLER_221_2019 ();
 b15zdnd11an1n32x5 FILLER_221_2083 ();
 b15zdnd11an1n16x5 FILLER_221_2115 ();
 b15zdnd11an1n08x5 FILLER_221_2131 ();
 b15zdnd11an1n04x5 FILLER_221_2139 ();
 b15zdnd11an1n08x5 FILLER_221_2154 ();
 b15zdnd00an1n01x5 FILLER_221_2162 ();
 b15zdnd11an1n04x5 FILLER_221_2167 ();
 b15zdnd11an1n08x5 FILLER_221_2187 ();
 b15zdnd11an1n32x5 FILLER_221_2237 ();
 b15zdnd11an1n08x5 FILLER_221_2269 ();
 b15zdnd11an1n04x5 FILLER_221_2277 ();
 b15zdnd00an1n02x5 FILLER_221_2281 ();
 b15zdnd00an1n01x5 FILLER_221_2283 ();
 b15zdnd11an1n64x5 FILLER_222_8 ();
 b15zdnd11an1n64x5 FILLER_222_72 ();
 b15zdnd11an1n64x5 FILLER_222_136 ();
 b15zdnd11an1n64x5 FILLER_222_200 ();
 b15zdnd11an1n64x5 FILLER_222_264 ();
 b15zdnd11an1n64x5 FILLER_222_328 ();
 b15zdnd11an1n64x5 FILLER_222_392 ();
 b15zdnd11an1n64x5 FILLER_222_456 ();
 b15zdnd11an1n64x5 FILLER_222_520 ();
 b15zdnd11an1n64x5 FILLER_222_584 ();
 b15zdnd11an1n64x5 FILLER_222_648 ();
 b15zdnd11an1n04x5 FILLER_222_712 ();
 b15zdnd00an1n02x5 FILLER_222_716 ();
 b15zdnd11an1n64x5 FILLER_222_726 ();
 b15zdnd11an1n64x5 FILLER_222_790 ();
 b15zdnd11an1n08x5 FILLER_222_854 ();
 b15zdnd11an1n64x5 FILLER_222_872 ();
 b15zdnd11an1n16x5 FILLER_222_936 ();
 b15zdnd11an1n08x5 FILLER_222_952 ();
 b15zdnd00an1n01x5 FILLER_222_960 ();
 b15zdnd11an1n64x5 FILLER_222_974 ();
 b15zdnd11an1n64x5 FILLER_222_1038 ();
 b15zdnd11an1n64x5 FILLER_222_1102 ();
 b15zdnd11an1n64x5 FILLER_222_1166 ();
 b15zdnd11an1n64x5 FILLER_222_1230 ();
 b15zdnd11an1n64x5 FILLER_222_1294 ();
 b15zdnd11an1n64x5 FILLER_222_1358 ();
 b15zdnd11an1n64x5 FILLER_222_1422 ();
 b15zdnd11an1n64x5 FILLER_222_1486 ();
 b15zdnd11an1n64x5 FILLER_222_1550 ();
 b15zdnd11an1n64x5 FILLER_222_1614 ();
 b15zdnd11an1n64x5 FILLER_222_1678 ();
 b15zdnd11an1n64x5 FILLER_222_1742 ();
 b15zdnd11an1n64x5 FILLER_222_1806 ();
 b15zdnd11an1n64x5 FILLER_222_1870 ();
 b15zdnd11an1n64x5 FILLER_222_1934 ();
 b15zdnd11an1n64x5 FILLER_222_1998 ();
 b15zdnd11an1n64x5 FILLER_222_2062 ();
 b15zdnd11an1n04x5 FILLER_222_2126 ();
 b15zdnd00an1n02x5 FILLER_222_2130 ();
 b15zdnd00an1n01x5 FILLER_222_2132 ();
 b15zdnd11an1n16x5 FILLER_222_2137 ();
 b15zdnd00an1n01x5 FILLER_222_2153 ();
 b15zdnd11an1n04x5 FILLER_222_2162 ();
 b15zdnd11an1n04x5 FILLER_222_2172 ();
 b15zdnd11an1n16x5 FILLER_222_2192 ();
 b15zdnd11an1n08x5 FILLER_222_2208 ();
 b15zdnd11an1n04x5 FILLER_222_2216 ();
 b15zdnd11an1n08x5 FILLER_222_2262 ();
 b15zdnd11an1n04x5 FILLER_222_2270 ();
 b15zdnd00an1n02x5 FILLER_222_2274 ();
 b15zdnd11an1n64x5 FILLER_223_0 ();
 b15zdnd11an1n64x5 FILLER_223_64 ();
 b15zdnd11an1n64x5 FILLER_223_128 ();
 b15zdnd11an1n64x5 FILLER_223_192 ();
 b15zdnd11an1n64x5 FILLER_223_256 ();
 b15zdnd11an1n64x5 FILLER_223_320 ();
 b15zdnd11an1n64x5 FILLER_223_384 ();
 b15zdnd11an1n16x5 FILLER_223_448 ();
 b15zdnd11an1n04x5 FILLER_223_464 ();
 b15zdnd00an1n01x5 FILLER_223_468 ();
 b15zdnd11an1n64x5 FILLER_223_481 ();
 b15zdnd11an1n64x5 FILLER_223_545 ();
 b15zdnd11an1n64x5 FILLER_223_609 ();
 b15zdnd11an1n64x5 FILLER_223_673 ();
 b15zdnd11an1n64x5 FILLER_223_737 ();
 b15zdnd11an1n64x5 FILLER_223_801 ();
 b15zdnd11an1n64x5 FILLER_223_865 ();
 b15zdnd11an1n64x5 FILLER_223_929 ();
 b15zdnd11an1n64x5 FILLER_223_993 ();
 b15zdnd11an1n64x5 FILLER_223_1057 ();
 b15zdnd11an1n64x5 FILLER_223_1121 ();
 b15zdnd11an1n64x5 FILLER_223_1185 ();
 b15zdnd11an1n64x5 FILLER_223_1249 ();
 b15zdnd11an1n16x5 FILLER_223_1313 ();
 b15zdnd11an1n08x5 FILLER_223_1329 ();
 b15zdnd11an1n04x5 FILLER_223_1337 ();
 b15zdnd11an1n64x5 FILLER_223_1383 ();
 b15zdnd11an1n64x5 FILLER_223_1447 ();
 b15zdnd11an1n64x5 FILLER_223_1511 ();
 b15zdnd11an1n64x5 FILLER_223_1575 ();
 b15zdnd11an1n64x5 FILLER_223_1639 ();
 b15zdnd11an1n64x5 FILLER_223_1703 ();
 b15zdnd11an1n64x5 FILLER_223_1767 ();
 b15zdnd11an1n64x5 FILLER_223_1831 ();
 b15zdnd11an1n64x5 FILLER_223_1895 ();
 b15zdnd11an1n08x5 FILLER_223_1959 ();
 b15zdnd00an1n02x5 FILLER_223_1967 ();
 b15zdnd00an1n01x5 FILLER_223_1969 ();
 b15zdnd11an1n64x5 FILLER_223_1979 ();
 b15zdnd11an1n64x5 FILLER_223_2043 ();
 b15zdnd11an1n32x5 FILLER_223_2107 ();
 b15zdnd11an1n04x5 FILLER_223_2139 ();
 b15zdnd00an1n02x5 FILLER_223_2143 ();
 b15zdnd00an1n01x5 FILLER_223_2145 ();
 b15zdnd11an1n32x5 FILLER_223_2152 ();
 b15zdnd11an1n16x5 FILLER_223_2184 ();
 b15zdnd11an1n32x5 FILLER_223_2242 ();
 b15zdnd11an1n08x5 FILLER_223_2274 ();
 b15zdnd00an1n02x5 FILLER_223_2282 ();
 b15zdnd11an1n64x5 FILLER_224_8 ();
 b15zdnd11an1n64x5 FILLER_224_72 ();
 b15zdnd11an1n64x5 FILLER_224_136 ();
 b15zdnd11an1n64x5 FILLER_224_200 ();
 b15zdnd11an1n64x5 FILLER_224_264 ();
 b15zdnd11an1n64x5 FILLER_224_328 ();
 b15zdnd11an1n64x5 FILLER_224_392 ();
 b15zdnd11an1n16x5 FILLER_224_456 ();
 b15zdnd11an1n04x5 FILLER_224_472 ();
 b15zdnd00an1n02x5 FILLER_224_476 ();
 b15zdnd11an1n64x5 FILLER_224_520 ();
 b15zdnd11an1n64x5 FILLER_224_584 ();
 b15zdnd11an1n64x5 FILLER_224_648 ();
 b15zdnd11an1n04x5 FILLER_224_712 ();
 b15zdnd00an1n02x5 FILLER_224_716 ();
 b15zdnd11an1n08x5 FILLER_224_726 ();
 b15zdnd11an1n04x5 FILLER_224_734 ();
 b15zdnd00an1n01x5 FILLER_224_738 ();
 b15zdnd11an1n16x5 FILLER_224_781 ();
 b15zdnd11an1n04x5 FILLER_224_797 ();
 b15zdnd00an1n02x5 FILLER_224_801 ();
 b15zdnd00an1n01x5 FILLER_224_803 ();
 b15zdnd11an1n64x5 FILLER_224_823 ();
 b15zdnd11an1n64x5 FILLER_224_887 ();
 b15zdnd11an1n64x5 FILLER_224_951 ();
 b15zdnd11an1n64x5 FILLER_224_1015 ();
 b15zdnd11an1n64x5 FILLER_224_1079 ();
 b15zdnd11an1n64x5 FILLER_224_1143 ();
 b15zdnd11an1n64x5 FILLER_224_1207 ();
 b15zdnd11an1n64x5 FILLER_224_1271 ();
 b15zdnd11an1n64x5 FILLER_224_1335 ();
 b15zdnd11an1n64x5 FILLER_224_1399 ();
 b15zdnd11an1n64x5 FILLER_224_1463 ();
 b15zdnd11an1n64x5 FILLER_224_1527 ();
 b15zdnd11an1n08x5 FILLER_224_1591 ();
 b15zdnd11an1n64x5 FILLER_224_1615 ();
 b15zdnd11an1n64x5 FILLER_224_1679 ();
 b15zdnd11an1n64x5 FILLER_224_1743 ();
 b15zdnd11an1n64x5 FILLER_224_1807 ();
 b15zdnd11an1n64x5 FILLER_224_1871 ();
 b15zdnd11an1n16x5 FILLER_224_1935 ();
 b15zdnd00an1n02x5 FILLER_224_1951 ();
 b15zdnd00an1n01x5 FILLER_224_1953 ();
 b15zdnd11an1n08x5 FILLER_224_1964 ();
 b15zdnd00an1n02x5 FILLER_224_1972 ();
 b15zdnd00an1n01x5 FILLER_224_1974 ();
 b15zdnd11an1n64x5 FILLER_224_1984 ();
 b15zdnd11an1n64x5 FILLER_224_2048 ();
 b15zdnd11an1n32x5 FILLER_224_2112 ();
 b15zdnd11an1n08x5 FILLER_224_2144 ();
 b15zdnd00an1n02x5 FILLER_224_2152 ();
 b15zdnd11an1n08x5 FILLER_224_2162 ();
 b15zdnd11an1n32x5 FILLER_224_2178 ();
 b15zdnd00an1n02x5 FILLER_224_2210 ();
 b15zdnd11an1n16x5 FILLER_224_2254 ();
 b15zdnd11an1n04x5 FILLER_224_2270 ();
 b15zdnd00an1n02x5 FILLER_224_2274 ();
 b15zdnd11an1n64x5 FILLER_225_0 ();
 b15zdnd11an1n64x5 FILLER_225_64 ();
 b15zdnd11an1n64x5 FILLER_225_128 ();
 b15zdnd11an1n64x5 FILLER_225_192 ();
 b15zdnd11an1n64x5 FILLER_225_256 ();
 b15zdnd11an1n64x5 FILLER_225_320 ();
 b15zdnd11an1n64x5 FILLER_225_384 ();
 b15zdnd11an1n16x5 FILLER_225_448 ();
 b15zdnd11an1n08x5 FILLER_225_464 ();
 b15zdnd11an1n04x5 FILLER_225_472 ();
 b15zdnd11an1n16x5 FILLER_225_484 ();
 b15zdnd00an1n02x5 FILLER_225_500 ();
 b15zdnd00an1n01x5 FILLER_225_502 ();
 b15zdnd11an1n64x5 FILLER_225_545 ();
 b15zdnd11an1n64x5 FILLER_225_609 ();
 b15zdnd11an1n64x5 FILLER_225_673 ();
 b15zdnd11an1n32x5 FILLER_225_737 ();
 b15zdnd11an1n08x5 FILLER_225_769 ();
 b15zdnd11an1n04x5 FILLER_225_777 ();
 b15zdnd00an1n02x5 FILLER_225_781 ();
 b15zdnd00an1n01x5 FILLER_225_783 ();
 b15zdnd11an1n64x5 FILLER_225_826 ();
 b15zdnd11an1n64x5 FILLER_225_890 ();
 b15zdnd11an1n64x5 FILLER_225_954 ();
 b15zdnd11an1n64x5 FILLER_225_1018 ();
 b15zdnd11an1n32x5 FILLER_225_1082 ();
 b15zdnd11an1n04x5 FILLER_225_1114 ();
 b15zdnd00an1n01x5 FILLER_225_1118 ();
 b15zdnd11an1n64x5 FILLER_225_1129 ();
 b15zdnd11an1n64x5 FILLER_225_1193 ();
 b15zdnd11an1n64x5 FILLER_225_1257 ();
 b15zdnd11an1n64x5 FILLER_225_1321 ();
 b15zdnd11an1n64x5 FILLER_225_1385 ();
 b15zdnd11an1n64x5 FILLER_225_1449 ();
 b15zdnd11an1n64x5 FILLER_225_1513 ();
 b15zdnd11an1n64x5 FILLER_225_1577 ();
 b15zdnd11an1n64x5 FILLER_225_1641 ();
 b15zdnd11an1n64x5 FILLER_225_1705 ();
 b15zdnd11an1n64x5 FILLER_225_1769 ();
 b15zdnd11an1n64x5 FILLER_225_1833 ();
 b15zdnd11an1n32x5 FILLER_225_1897 ();
 b15zdnd11an1n04x5 FILLER_225_1929 ();
 b15zdnd00an1n02x5 FILLER_225_1933 ();
 b15zdnd00an1n01x5 FILLER_225_1935 ();
 b15zdnd11an1n16x5 FILLER_225_1948 ();
 b15zdnd11an1n64x5 FILLER_225_1974 ();
 b15zdnd11an1n64x5 FILLER_225_2038 ();
 b15zdnd11an1n64x5 FILLER_225_2102 ();
 b15zdnd00an1n02x5 FILLER_225_2166 ();
 b15zdnd00an1n01x5 FILLER_225_2168 ();
 b15zdnd11an1n16x5 FILLER_225_2173 ();
 b15zdnd11an1n08x5 FILLER_225_2189 ();
 b15zdnd11an1n08x5 FILLER_225_2239 ();
 b15zdnd00an1n01x5 FILLER_225_2247 ();
 b15zdnd11an1n32x5 FILLER_225_2252 ();
 b15zdnd11an1n64x5 FILLER_226_8 ();
 b15zdnd11an1n64x5 FILLER_226_72 ();
 b15zdnd11an1n64x5 FILLER_226_136 ();
 b15zdnd11an1n64x5 FILLER_226_200 ();
 b15zdnd11an1n64x5 FILLER_226_264 ();
 b15zdnd11an1n64x5 FILLER_226_328 ();
 b15zdnd11an1n64x5 FILLER_226_392 ();
 b15zdnd11an1n64x5 FILLER_226_456 ();
 b15zdnd11an1n64x5 FILLER_226_520 ();
 b15zdnd11an1n32x5 FILLER_226_584 ();
 b15zdnd00an1n02x5 FILLER_226_616 ();
 b15zdnd00an1n01x5 FILLER_226_618 ();
 b15zdnd11an1n64x5 FILLER_226_629 ();
 b15zdnd11an1n16x5 FILLER_226_693 ();
 b15zdnd11an1n08x5 FILLER_226_709 ();
 b15zdnd00an1n01x5 FILLER_226_717 ();
 b15zdnd11an1n32x5 FILLER_226_726 ();
 b15zdnd11an1n16x5 FILLER_226_758 ();
 b15zdnd11an1n04x5 FILLER_226_774 ();
 b15zdnd00an1n02x5 FILLER_226_778 ();
 b15zdnd00an1n01x5 FILLER_226_780 ();
 b15zdnd11an1n64x5 FILLER_226_800 ();
 b15zdnd11an1n64x5 FILLER_226_864 ();
 b15zdnd11an1n64x5 FILLER_226_928 ();
 b15zdnd11an1n64x5 FILLER_226_992 ();
 b15zdnd11an1n64x5 FILLER_226_1056 ();
 b15zdnd11an1n64x5 FILLER_226_1120 ();
 b15zdnd11an1n64x5 FILLER_226_1184 ();
 b15zdnd11an1n64x5 FILLER_226_1248 ();
 b15zdnd11an1n64x5 FILLER_226_1312 ();
 b15zdnd11an1n64x5 FILLER_226_1376 ();
 b15zdnd11an1n64x5 FILLER_226_1440 ();
 b15zdnd11an1n64x5 FILLER_226_1504 ();
 b15zdnd11an1n64x5 FILLER_226_1568 ();
 b15zdnd11an1n64x5 FILLER_226_1632 ();
 b15zdnd11an1n16x5 FILLER_226_1696 ();
 b15zdnd11an1n08x5 FILLER_226_1712 ();
 b15zdnd11an1n04x5 FILLER_226_1720 ();
 b15zdnd00an1n02x5 FILLER_226_1724 ();
 b15zdnd00an1n01x5 FILLER_226_1726 ();
 b15zdnd11an1n64x5 FILLER_226_1736 ();
 b15zdnd11an1n64x5 FILLER_226_1800 ();
 b15zdnd11an1n64x5 FILLER_226_1864 ();
 b15zdnd11an1n16x5 FILLER_226_1928 ();
 b15zdnd00an1n01x5 FILLER_226_1944 ();
 b15zdnd11an1n04x5 FILLER_226_1957 ();
 b15zdnd00an1n02x5 FILLER_226_1961 ();
 b15zdnd11an1n32x5 FILLER_226_1973 ();
 b15zdnd00an1n02x5 FILLER_226_2005 ();
 b15zdnd00an1n01x5 FILLER_226_2007 ();
 b15zdnd11an1n64x5 FILLER_226_2028 ();
 b15zdnd11an1n16x5 FILLER_226_2092 ();
 b15zdnd11an1n08x5 FILLER_226_2108 ();
 b15zdnd11an1n04x5 FILLER_226_2116 ();
 b15zdnd00an1n02x5 FILLER_226_2120 ();
 b15zdnd11an1n16x5 FILLER_226_2130 ();
 b15zdnd11an1n08x5 FILLER_226_2146 ();
 b15zdnd11an1n32x5 FILLER_226_2162 ();
 b15zdnd11an1n16x5 FILLER_226_2194 ();
 b15zdnd11an1n04x5 FILLER_226_2252 ();
 b15zdnd11an1n16x5 FILLER_226_2260 ();
 b15zdnd11an1n64x5 FILLER_227_0 ();
 b15zdnd11an1n64x5 FILLER_227_64 ();
 b15zdnd11an1n64x5 FILLER_227_128 ();
 b15zdnd11an1n64x5 FILLER_227_192 ();
 b15zdnd11an1n64x5 FILLER_227_256 ();
 b15zdnd11an1n64x5 FILLER_227_320 ();
 b15zdnd11an1n64x5 FILLER_227_384 ();
 b15zdnd11an1n64x5 FILLER_227_448 ();
 b15zdnd11an1n64x5 FILLER_227_512 ();
 b15zdnd11an1n64x5 FILLER_227_576 ();
 b15zdnd11an1n16x5 FILLER_227_640 ();
 b15zdnd11an1n08x5 FILLER_227_656 ();
 b15zdnd00an1n01x5 FILLER_227_664 ();
 b15zdnd11an1n64x5 FILLER_227_674 ();
 b15zdnd11an1n64x5 FILLER_227_738 ();
 b15zdnd11an1n32x5 FILLER_227_821 ();
 b15zdnd11an1n04x5 FILLER_227_853 ();
 b15zdnd00an1n01x5 FILLER_227_857 ();
 b15zdnd11an1n64x5 FILLER_227_880 ();
 b15zdnd11an1n64x5 FILLER_227_944 ();
 b15zdnd11an1n64x5 FILLER_227_1008 ();
 b15zdnd11an1n64x5 FILLER_227_1072 ();
 b15zdnd11an1n64x5 FILLER_227_1136 ();
 b15zdnd11an1n32x5 FILLER_227_1200 ();
 b15zdnd11an1n16x5 FILLER_227_1232 ();
 b15zdnd11an1n08x5 FILLER_227_1248 ();
 b15zdnd00an1n01x5 FILLER_227_1256 ();
 b15zdnd11an1n16x5 FILLER_227_1268 ();
 b15zdnd11an1n04x5 FILLER_227_1284 ();
 b15zdnd00an1n01x5 FILLER_227_1288 ();
 b15zdnd11an1n64x5 FILLER_227_1295 ();
 b15zdnd11an1n64x5 FILLER_227_1359 ();
 b15zdnd11an1n64x5 FILLER_227_1423 ();
 b15zdnd11an1n64x5 FILLER_227_1487 ();
 b15zdnd11an1n64x5 FILLER_227_1551 ();
 b15zdnd11an1n64x5 FILLER_227_1615 ();
 b15zdnd11an1n08x5 FILLER_227_1679 ();
 b15zdnd00an1n01x5 FILLER_227_1687 ();
 b15zdnd11an1n04x5 FILLER_227_1730 ();
 b15zdnd11an1n04x5 FILLER_227_1748 ();
 b15zdnd11an1n64x5 FILLER_227_1761 ();
 b15zdnd11an1n64x5 FILLER_227_1825 ();
 b15zdnd11an1n32x5 FILLER_227_1889 ();
 b15zdnd11an1n04x5 FILLER_227_1921 ();
 b15zdnd00an1n02x5 FILLER_227_1925 ();
 b15zdnd11an1n04x5 FILLER_227_1939 ();
 b15zdnd11an1n64x5 FILLER_227_1955 ();
 b15zdnd11an1n64x5 FILLER_227_2019 ();
 b15zdnd11an1n64x5 FILLER_227_2083 ();
 b15zdnd11an1n64x5 FILLER_227_2147 ();
 b15zdnd11an1n32x5 FILLER_227_2211 ();
 b15zdnd00an1n01x5 FILLER_227_2243 ();
 b15zdnd11an1n32x5 FILLER_227_2248 ();
 b15zdnd11an1n04x5 FILLER_227_2280 ();
 b15zdnd11an1n64x5 FILLER_228_8 ();
 b15zdnd11an1n64x5 FILLER_228_72 ();
 b15zdnd11an1n64x5 FILLER_228_136 ();
 b15zdnd11an1n64x5 FILLER_228_200 ();
 b15zdnd11an1n64x5 FILLER_228_264 ();
 b15zdnd11an1n64x5 FILLER_228_328 ();
 b15zdnd11an1n64x5 FILLER_228_392 ();
 b15zdnd11an1n64x5 FILLER_228_456 ();
 b15zdnd11an1n32x5 FILLER_228_520 ();
 b15zdnd11an1n08x5 FILLER_228_552 ();
 b15zdnd11an1n04x5 FILLER_228_560 ();
 b15zdnd00an1n01x5 FILLER_228_564 ();
 b15zdnd11an1n32x5 FILLER_228_585 ();
 b15zdnd11an1n16x5 FILLER_228_617 ();
 b15zdnd11an1n08x5 FILLER_228_633 ();
 b15zdnd11an1n04x5 FILLER_228_641 ();
 b15zdnd11an1n64x5 FILLER_228_652 ();
 b15zdnd00an1n02x5 FILLER_228_716 ();
 b15zdnd11an1n64x5 FILLER_228_726 ();
 b15zdnd11an1n64x5 FILLER_228_790 ();
 b15zdnd11an1n64x5 FILLER_228_854 ();
 b15zdnd11an1n64x5 FILLER_228_918 ();
 b15zdnd11an1n16x5 FILLER_228_982 ();
 b15zdnd00an1n02x5 FILLER_228_998 ();
 b15zdnd00an1n01x5 FILLER_228_1000 ();
 b15zdnd11an1n64x5 FILLER_228_1046 ();
 b15zdnd11an1n64x5 FILLER_228_1110 ();
 b15zdnd11an1n64x5 FILLER_228_1174 ();
 b15zdnd11an1n64x5 FILLER_228_1238 ();
 b15zdnd11an1n32x5 FILLER_228_1302 ();
 b15zdnd11an1n08x5 FILLER_228_1334 ();
 b15zdnd11an1n04x5 FILLER_228_1342 ();
 b15zdnd11an1n64x5 FILLER_228_1388 ();
 b15zdnd11an1n64x5 FILLER_228_1452 ();
 b15zdnd11an1n64x5 FILLER_228_1516 ();
 b15zdnd11an1n64x5 FILLER_228_1580 ();
 b15zdnd11an1n32x5 FILLER_228_1644 ();
 b15zdnd11an1n04x5 FILLER_228_1676 ();
 b15zdnd00an1n02x5 FILLER_228_1680 ();
 b15zdnd00an1n01x5 FILLER_228_1682 ();
 b15zdnd11an1n08x5 FILLER_228_1699 ();
 b15zdnd11an1n04x5 FILLER_228_1707 ();
 b15zdnd00an1n01x5 FILLER_228_1711 ();
 b15zdnd11an1n64x5 FILLER_228_1754 ();
 b15zdnd11an1n64x5 FILLER_228_1818 ();
 b15zdnd11an1n64x5 FILLER_228_1882 ();
 b15zdnd11an1n64x5 FILLER_228_1946 ();
 b15zdnd11an1n64x5 FILLER_228_2010 ();
 b15zdnd11an1n64x5 FILLER_228_2074 ();
 b15zdnd11an1n16x5 FILLER_228_2138 ();
 b15zdnd11an1n64x5 FILLER_228_2162 ();
 b15zdnd11an1n16x5 FILLER_228_2226 ();
 b15zdnd11an1n08x5 FILLER_228_2242 ();
 b15zdnd11an1n04x5 FILLER_228_2250 ();
 b15zdnd11an1n16x5 FILLER_228_2258 ();
 b15zdnd00an1n02x5 FILLER_228_2274 ();
 b15zdnd11an1n64x5 FILLER_229_0 ();
 b15zdnd11an1n64x5 FILLER_229_64 ();
 b15zdnd11an1n64x5 FILLER_229_128 ();
 b15zdnd11an1n64x5 FILLER_229_192 ();
 b15zdnd11an1n64x5 FILLER_229_256 ();
 b15zdnd11an1n64x5 FILLER_229_320 ();
 b15zdnd11an1n64x5 FILLER_229_384 ();
 b15zdnd11an1n64x5 FILLER_229_448 ();
 b15zdnd11an1n16x5 FILLER_229_512 ();
 b15zdnd11an1n08x5 FILLER_229_528 ();
 b15zdnd11an1n04x5 FILLER_229_536 ();
 b15zdnd00an1n02x5 FILLER_229_540 ();
 b15zdnd00an1n01x5 FILLER_229_542 ();
 b15zdnd11an1n64x5 FILLER_229_564 ();
 b15zdnd11an1n64x5 FILLER_229_628 ();
 b15zdnd11an1n32x5 FILLER_229_692 ();
 b15zdnd11an1n16x5 FILLER_229_724 ();
 b15zdnd11an1n08x5 FILLER_229_740 ();
 b15zdnd11an1n04x5 FILLER_229_748 ();
 b15zdnd00an1n02x5 FILLER_229_752 ();
 b15zdnd11an1n32x5 FILLER_229_762 ();
 b15zdnd11an1n16x5 FILLER_229_794 ();
 b15zdnd00an1n02x5 FILLER_229_810 ();
 b15zdnd11an1n64x5 FILLER_229_836 ();
 b15zdnd11an1n64x5 FILLER_229_900 ();
 b15zdnd11an1n64x5 FILLER_229_964 ();
 b15zdnd11an1n64x5 FILLER_229_1028 ();
 b15zdnd11an1n32x5 FILLER_229_1092 ();
 b15zdnd11an1n16x5 FILLER_229_1124 ();
 b15zdnd00an1n01x5 FILLER_229_1140 ();
 b15zdnd11an1n64x5 FILLER_229_1157 ();
 b15zdnd11an1n64x5 FILLER_229_1221 ();
 b15zdnd11an1n64x5 FILLER_229_1285 ();
 b15zdnd11an1n64x5 FILLER_229_1349 ();
 b15zdnd11an1n64x5 FILLER_229_1413 ();
 b15zdnd11an1n64x5 FILLER_229_1477 ();
 b15zdnd11an1n64x5 FILLER_229_1541 ();
 b15zdnd11an1n32x5 FILLER_229_1605 ();
 b15zdnd11an1n16x5 FILLER_229_1637 ();
 b15zdnd00an1n02x5 FILLER_229_1653 ();
 b15zdnd00an1n01x5 FILLER_229_1655 ();
 b15zdnd11an1n16x5 FILLER_229_1698 ();
 b15zdnd11an1n04x5 FILLER_229_1756 ();
 b15zdnd11an1n64x5 FILLER_229_1766 ();
 b15zdnd11an1n64x5 FILLER_229_1830 ();
 b15zdnd11an1n64x5 FILLER_229_1894 ();
 b15zdnd11an1n64x5 FILLER_229_1958 ();
 b15zdnd11an1n64x5 FILLER_229_2022 ();
 b15zdnd11an1n64x5 FILLER_229_2086 ();
 b15zdnd11an1n64x5 FILLER_229_2150 ();
 b15zdnd11an1n64x5 FILLER_229_2214 ();
 b15zdnd11an1n04x5 FILLER_229_2278 ();
 b15zdnd00an1n02x5 FILLER_229_2282 ();
 b15zdnd11an1n64x5 FILLER_230_8 ();
 b15zdnd11an1n64x5 FILLER_230_72 ();
 b15zdnd11an1n64x5 FILLER_230_136 ();
 b15zdnd11an1n64x5 FILLER_230_200 ();
 b15zdnd11an1n64x5 FILLER_230_264 ();
 b15zdnd11an1n64x5 FILLER_230_328 ();
 b15zdnd11an1n64x5 FILLER_230_392 ();
 b15zdnd11an1n64x5 FILLER_230_456 ();
 b15zdnd11an1n64x5 FILLER_230_520 ();
 b15zdnd11an1n32x5 FILLER_230_584 ();
 b15zdnd11an1n04x5 FILLER_230_616 ();
 b15zdnd00an1n01x5 FILLER_230_620 ();
 b15zdnd11an1n32x5 FILLER_230_663 ();
 b15zdnd11an1n16x5 FILLER_230_695 ();
 b15zdnd11an1n04x5 FILLER_230_711 ();
 b15zdnd00an1n02x5 FILLER_230_715 ();
 b15zdnd00an1n01x5 FILLER_230_717 ();
 b15zdnd11an1n64x5 FILLER_230_726 ();
 b15zdnd11an1n64x5 FILLER_230_790 ();
 b15zdnd11an1n64x5 FILLER_230_854 ();
 b15zdnd11an1n32x5 FILLER_230_918 ();
 b15zdnd11an1n16x5 FILLER_230_950 ();
 b15zdnd11an1n08x5 FILLER_230_966 ();
 b15zdnd00an1n01x5 FILLER_230_974 ();
 b15zdnd11an1n64x5 FILLER_230_981 ();
 b15zdnd11an1n64x5 FILLER_230_1045 ();
 b15zdnd11an1n64x5 FILLER_230_1109 ();
 b15zdnd11an1n64x5 FILLER_230_1173 ();
 b15zdnd11an1n64x5 FILLER_230_1237 ();
 b15zdnd11an1n64x5 FILLER_230_1301 ();
 b15zdnd11an1n64x5 FILLER_230_1365 ();
 b15zdnd11an1n64x5 FILLER_230_1429 ();
 b15zdnd11an1n64x5 FILLER_230_1493 ();
 b15zdnd11an1n64x5 FILLER_230_1557 ();
 b15zdnd11an1n64x5 FILLER_230_1621 ();
 b15zdnd11an1n16x5 FILLER_230_1685 ();
 b15zdnd00an1n02x5 FILLER_230_1701 ();
 b15zdnd11an1n04x5 FILLER_230_1719 ();
 b15zdnd00an1n01x5 FILLER_230_1723 ();
 b15zdnd11an1n08x5 FILLER_230_1738 ();
 b15zdnd00an1n02x5 FILLER_230_1746 ();
 b15zdnd00an1n01x5 FILLER_230_1748 ();
 b15zdnd11an1n64x5 FILLER_230_1765 ();
 b15zdnd11an1n64x5 FILLER_230_1829 ();
 b15zdnd11an1n64x5 FILLER_230_1893 ();
 b15zdnd11an1n64x5 FILLER_230_1957 ();
 b15zdnd11an1n64x5 FILLER_230_2021 ();
 b15zdnd11an1n64x5 FILLER_230_2085 ();
 b15zdnd11an1n04x5 FILLER_230_2149 ();
 b15zdnd00an1n01x5 FILLER_230_2153 ();
 b15zdnd11an1n64x5 FILLER_230_2162 ();
 b15zdnd11an1n32x5 FILLER_230_2226 ();
 b15zdnd11an1n16x5 FILLER_230_2258 ();
 b15zdnd00an1n02x5 FILLER_230_2274 ();
 b15zdnd11an1n64x5 FILLER_231_0 ();
 b15zdnd11an1n64x5 FILLER_231_64 ();
 b15zdnd11an1n64x5 FILLER_231_128 ();
 b15zdnd11an1n64x5 FILLER_231_192 ();
 b15zdnd11an1n64x5 FILLER_231_256 ();
 b15zdnd11an1n64x5 FILLER_231_320 ();
 b15zdnd11an1n64x5 FILLER_231_384 ();
 b15zdnd11an1n64x5 FILLER_231_448 ();
 b15zdnd11an1n64x5 FILLER_231_512 ();
 b15zdnd11an1n64x5 FILLER_231_576 ();
 b15zdnd11an1n64x5 FILLER_231_640 ();
 b15zdnd11an1n04x5 FILLER_231_704 ();
 b15zdnd00an1n02x5 FILLER_231_708 ();
 b15zdnd00an1n01x5 FILLER_231_710 ();
 b15zdnd11an1n64x5 FILLER_231_727 ();
 b15zdnd11an1n64x5 FILLER_231_791 ();
 b15zdnd11an1n64x5 FILLER_231_855 ();
 b15zdnd11an1n64x5 FILLER_231_919 ();
 b15zdnd11an1n64x5 FILLER_231_983 ();
 b15zdnd11an1n16x5 FILLER_231_1047 ();
 b15zdnd11an1n04x5 FILLER_231_1063 ();
 b15zdnd00an1n02x5 FILLER_231_1067 ();
 b15zdnd11an1n64x5 FILLER_231_1076 ();
 b15zdnd11an1n64x5 FILLER_231_1140 ();
 b15zdnd11an1n08x5 FILLER_231_1204 ();
 b15zdnd00an1n01x5 FILLER_231_1212 ();
 b15zdnd11an1n64x5 FILLER_231_1258 ();
 b15zdnd11an1n64x5 FILLER_231_1322 ();
 b15zdnd11an1n64x5 FILLER_231_1386 ();
 b15zdnd11an1n64x5 FILLER_231_1450 ();
 b15zdnd11an1n64x5 FILLER_231_1514 ();
 b15zdnd11an1n64x5 FILLER_231_1578 ();
 b15zdnd11an1n32x5 FILLER_231_1642 ();
 b15zdnd11an1n16x5 FILLER_231_1674 ();
 b15zdnd00an1n02x5 FILLER_231_1690 ();
 b15zdnd11an1n16x5 FILLER_231_1734 ();
 b15zdnd00an1n02x5 FILLER_231_1750 ();
 b15zdnd00an1n01x5 FILLER_231_1752 ();
 b15zdnd11an1n64x5 FILLER_231_1764 ();
 b15zdnd11an1n64x5 FILLER_231_1828 ();
 b15zdnd11an1n64x5 FILLER_231_1892 ();
 b15zdnd11an1n64x5 FILLER_231_1956 ();
 b15zdnd11an1n64x5 FILLER_231_2020 ();
 b15zdnd11an1n64x5 FILLER_231_2084 ();
 b15zdnd11an1n64x5 FILLER_231_2148 ();
 b15zdnd11an1n64x5 FILLER_231_2212 ();
 b15zdnd11an1n08x5 FILLER_231_2276 ();
 b15zdnd11an1n64x5 FILLER_232_8 ();
 b15zdnd11an1n64x5 FILLER_232_72 ();
 b15zdnd11an1n64x5 FILLER_232_136 ();
 b15zdnd11an1n64x5 FILLER_232_200 ();
 b15zdnd11an1n64x5 FILLER_232_264 ();
 b15zdnd11an1n64x5 FILLER_232_328 ();
 b15zdnd11an1n64x5 FILLER_232_392 ();
 b15zdnd11an1n64x5 FILLER_232_456 ();
 b15zdnd11an1n64x5 FILLER_232_520 ();
 b15zdnd00an1n02x5 FILLER_232_584 ();
 b15zdnd11an1n04x5 FILLER_232_602 ();
 b15zdnd00an1n02x5 FILLER_232_606 ();
 b15zdnd00an1n01x5 FILLER_232_608 ();
 b15zdnd11an1n64x5 FILLER_232_651 ();
 b15zdnd00an1n02x5 FILLER_232_715 ();
 b15zdnd00an1n01x5 FILLER_232_717 ();
 b15zdnd11an1n64x5 FILLER_232_726 ();
 b15zdnd11an1n64x5 FILLER_232_790 ();
 b15zdnd11an1n64x5 FILLER_232_854 ();
 b15zdnd11an1n64x5 FILLER_232_918 ();
 b15zdnd11an1n64x5 FILLER_232_982 ();
 b15zdnd11an1n08x5 FILLER_232_1046 ();
 b15zdnd11an1n04x5 FILLER_232_1054 ();
 b15zdnd00an1n01x5 FILLER_232_1058 ();
 b15zdnd11an1n64x5 FILLER_232_1066 ();
 b15zdnd11an1n64x5 FILLER_232_1130 ();
 b15zdnd11an1n32x5 FILLER_232_1194 ();
 b15zdnd11an1n04x5 FILLER_232_1226 ();
 b15zdnd11an1n64x5 FILLER_232_1275 ();
 b15zdnd11an1n64x5 FILLER_232_1339 ();
 b15zdnd11an1n64x5 FILLER_232_1403 ();
 b15zdnd11an1n64x5 FILLER_232_1467 ();
 b15zdnd11an1n64x5 FILLER_232_1531 ();
 b15zdnd11an1n64x5 FILLER_232_1595 ();
 b15zdnd11an1n64x5 FILLER_232_1659 ();
 b15zdnd11an1n64x5 FILLER_232_1723 ();
 b15zdnd11an1n64x5 FILLER_232_1787 ();
 b15zdnd11an1n64x5 FILLER_232_1851 ();
 b15zdnd11an1n64x5 FILLER_232_1915 ();
 b15zdnd11an1n64x5 FILLER_232_1979 ();
 b15zdnd11an1n64x5 FILLER_232_2043 ();
 b15zdnd11an1n32x5 FILLER_232_2107 ();
 b15zdnd11an1n08x5 FILLER_232_2139 ();
 b15zdnd11an1n04x5 FILLER_232_2147 ();
 b15zdnd00an1n02x5 FILLER_232_2151 ();
 b15zdnd00an1n01x5 FILLER_232_2153 ();
 b15zdnd11an1n64x5 FILLER_232_2162 ();
 b15zdnd11an1n32x5 FILLER_232_2226 ();
 b15zdnd11an1n16x5 FILLER_232_2258 ();
 b15zdnd00an1n02x5 FILLER_232_2274 ();
 b15zdnd11an1n64x5 FILLER_233_0 ();
 b15zdnd11an1n64x5 FILLER_233_64 ();
 b15zdnd11an1n64x5 FILLER_233_128 ();
 b15zdnd11an1n64x5 FILLER_233_192 ();
 b15zdnd11an1n64x5 FILLER_233_256 ();
 b15zdnd11an1n64x5 FILLER_233_320 ();
 b15zdnd11an1n64x5 FILLER_233_384 ();
 b15zdnd11an1n64x5 FILLER_233_448 ();
 b15zdnd11an1n64x5 FILLER_233_512 ();
 b15zdnd11an1n64x5 FILLER_233_576 ();
 b15zdnd11an1n64x5 FILLER_233_640 ();
 b15zdnd11an1n64x5 FILLER_233_704 ();
 b15zdnd11an1n32x5 FILLER_233_768 ();
 b15zdnd11an1n16x5 FILLER_233_800 ();
 b15zdnd11an1n08x5 FILLER_233_816 ();
 b15zdnd11an1n04x5 FILLER_233_824 ();
 b15zdnd00an1n02x5 FILLER_233_828 ();
 b15zdnd00an1n01x5 FILLER_233_830 ();
 b15zdnd11an1n64x5 FILLER_233_850 ();
 b15zdnd11an1n64x5 FILLER_233_914 ();
 b15zdnd11an1n64x5 FILLER_233_978 ();
 b15zdnd11an1n64x5 FILLER_233_1042 ();
 b15zdnd11an1n04x5 FILLER_233_1106 ();
 b15zdnd00an1n02x5 FILLER_233_1110 ();
 b15zdnd11an1n64x5 FILLER_233_1157 ();
 b15zdnd11an1n16x5 FILLER_233_1221 ();
 b15zdnd11an1n08x5 FILLER_233_1237 ();
 b15zdnd11an1n04x5 FILLER_233_1245 ();
 b15zdnd00an1n02x5 FILLER_233_1249 ();
 b15zdnd11an1n64x5 FILLER_233_1296 ();
 b15zdnd11an1n64x5 FILLER_233_1360 ();
 b15zdnd11an1n64x5 FILLER_233_1424 ();
 b15zdnd11an1n64x5 FILLER_233_1488 ();
 b15zdnd11an1n64x5 FILLER_233_1552 ();
 b15zdnd11an1n64x5 FILLER_233_1616 ();
 b15zdnd11an1n64x5 FILLER_233_1680 ();
 b15zdnd11an1n64x5 FILLER_233_1744 ();
 b15zdnd11an1n64x5 FILLER_233_1808 ();
 b15zdnd11an1n64x5 FILLER_233_1872 ();
 b15zdnd11an1n64x5 FILLER_233_1936 ();
 b15zdnd11an1n64x5 FILLER_233_2000 ();
 b15zdnd11an1n64x5 FILLER_233_2064 ();
 b15zdnd11an1n64x5 FILLER_233_2128 ();
 b15zdnd11an1n64x5 FILLER_233_2192 ();
 b15zdnd11an1n16x5 FILLER_233_2256 ();
 b15zdnd11an1n08x5 FILLER_233_2272 ();
 b15zdnd11an1n04x5 FILLER_233_2280 ();
 b15zdnd11an1n64x5 FILLER_234_8 ();
 b15zdnd11an1n64x5 FILLER_234_72 ();
 b15zdnd11an1n64x5 FILLER_234_136 ();
 b15zdnd11an1n64x5 FILLER_234_200 ();
 b15zdnd11an1n64x5 FILLER_234_264 ();
 b15zdnd11an1n64x5 FILLER_234_328 ();
 b15zdnd11an1n64x5 FILLER_234_392 ();
 b15zdnd11an1n64x5 FILLER_234_456 ();
 b15zdnd11an1n64x5 FILLER_234_520 ();
 b15zdnd11an1n64x5 FILLER_234_584 ();
 b15zdnd11an1n64x5 FILLER_234_648 ();
 b15zdnd11an1n04x5 FILLER_234_712 ();
 b15zdnd00an1n02x5 FILLER_234_716 ();
 b15zdnd11an1n08x5 FILLER_234_726 ();
 b15zdnd00an1n01x5 FILLER_234_734 ();
 b15zdnd11an1n64x5 FILLER_234_743 ();
 b15zdnd11an1n64x5 FILLER_234_807 ();
 b15zdnd11an1n64x5 FILLER_234_871 ();
 b15zdnd11an1n64x5 FILLER_234_935 ();
 b15zdnd11an1n64x5 FILLER_234_999 ();
 b15zdnd11an1n64x5 FILLER_234_1063 ();
 b15zdnd11an1n64x5 FILLER_234_1159 ();
 b15zdnd11an1n32x5 FILLER_234_1223 ();
 b15zdnd11an1n08x5 FILLER_234_1255 ();
 b15zdnd11an1n04x5 FILLER_234_1263 ();
 b15zdnd00an1n02x5 FILLER_234_1267 ();
 b15zdnd00an1n01x5 FILLER_234_1269 ();
 b15zdnd11an1n64x5 FILLER_234_1312 ();
 b15zdnd11an1n64x5 FILLER_234_1376 ();
 b15zdnd11an1n64x5 FILLER_234_1440 ();
 b15zdnd11an1n64x5 FILLER_234_1504 ();
 b15zdnd11an1n64x5 FILLER_234_1568 ();
 b15zdnd11an1n64x5 FILLER_234_1632 ();
 b15zdnd11an1n64x5 FILLER_234_1696 ();
 b15zdnd11an1n64x5 FILLER_234_1760 ();
 b15zdnd11an1n64x5 FILLER_234_1824 ();
 b15zdnd11an1n64x5 FILLER_234_1888 ();
 b15zdnd11an1n64x5 FILLER_234_1952 ();
 b15zdnd11an1n64x5 FILLER_234_2016 ();
 b15zdnd11an1n64x5 FILLER_234_2080 ();
 b15zdnd11an1n08x5 FILLER_234_2144 ();
 b15zdnd00an1n02x5 FILLER_234_2152 ();
 b15zdnd11an1n64x5 FILLER_234_2162 ();
 b15zdnd11an1n32x5 FILLER_234_2226 ();
 b15zdnd11an1n16x5 FILLER_234_2258 ();
 b15zdnd00an1n02x5 FILLER_234_2274 ();
 b15zdnd11an1n64x5 FILLER_235_0 ();
 b15zdnd11an1n64x5 FILLER_235_64 ();
 b15zdnd11an1n64x5 FILLER_235_128 ();
 b15zdnd11an1n64x5 FILLER_235_192 ();
 b15zdnd11an1n64x5 FILLER_235_256 ();
 b15zdnd11an1n64x5 FILLER_235_320 ();
 b15zdnd11an1n64x5 FILLER_235_384 ();
 b15zdnd11an1n64x5 FILLER_235_448 ();
 b15zdnd11an1n64x5 FILLER_235_512 ();
 b15zdnd11an1n64x5 FILLER_235_576 ();
 b15zdnd11an1n08x5 FILLER_235_640 ();
 b15zdnd00an1n01x5 FILLER_235_648 ();
 b15zdnd11an1n64x5 FILLER_235_691 ();
 b15zdnd11an1n64x5 FILLER_235_755 ();
 b15zdnd11an1n64x5 FILLER_235_819 ();
 b15zdnd11an1n64x5 FILLER_235_883 ();
 b15zdnd11an1n64x5 FILLER_235_947 ();
 b15zdnd11an1n64x5 FILLER_235_1011 ();
 b15zdnd11an1n64x5 FILLER_235_1075 ();
 b15zdnd11an1n64x5 FILLER_235_1139 ();
 b15zdnd11an1n64x5 FILLER_235_1203 ();
 b15zdnd11an1n64x5 FILLER_235_1267 ();
 b15zdnd11an1n64x5 FILLER_235_1331 ();
 b15zdnd11an1n64x5 FILLER_235_1395 ();
 b15zdnd11an1n64x5 FILLER_235_1459 ();
 b15zdnd11an1n64x5 FILLER_235_1523 ();
 b15zdnd11an1n64x5 FILLER_235_1587 ();
 b15zdnd11an1n64x5 FILLER_235_1651 ();
 b15zdnd11an1n64x5 FILLER_235_1715 ();
 b15zdnd11an1n64x5 FILLER_235_1779 ();
 b15zdnd11an1n64x5 FILLER_235_1843 ();
 b15zdnd11an1n64x5 FILLER_235_1907 ();
 b15zdnd11an1n64x5 FILLER_235_1971 ();
 b15zdnd11an1n64x5 FILLER_235_2035 ();
 b15zdnd11an1n64x5 FILLER_235_2099 ();
 b15zdnd11an1n64x5 FILLER_235_2163 ();
 b15zdnd11an1n32x5 FILLER_235_2227 ();
 b15zdnd11an1n16x5 FILLER_235_2259 ();
 b15zdnd11an1n08x5 FILLER_235_2275 ();
 b15zdnd00an1n01x5 FILLER_235_2283 ();
 b15zdnd11an1n64x5 FILLER_236_8 ();
 b15zdnd11an1n64x5 FILLER_236_72 ();
 b15zdnd11an1n64x5 FILLER_236_136 ();
 b15zdnd11an1n64x5 FILLER_236_200 ();
 b15zdnd11an1n64x5 FILLER_236_264 ();
 b15zdnd11an1n64x5 FILLER_236_328 ();
 b15zdnd11an1n64x5 FILLER_236_392 ();
 b15zdnd11an1n64x5 FILLER_236_456 ();
 b15zdnd11an1n64x5 FILLER_236_520 ();
 b15zdnd11an1n64x5 FILLER_236_584 ();
 b15zdnd11an1n64x5 FILLER_236_648 ();
 b15zdnd11an1n04x5 FILLER_236_712 ();
 b15zdnd00an1n02x5 FILLER_236_716 ();
 b15zdnd11an1n64x5 FILLER_236_726 ();
 b15zdnd11an1n64x5 FILLER_236_790 ();
 b15zdnd11an1n64x5 FILLER_236_854 ();
 b15zdnd11an1n64x5 FILLER_236_918 ();
 b15zdnd11an1n64x5 FILLER_236_982 ();
 b15zdnd11an1n64x5 FILLER_236_1046 ();
 b15zdnd11an1n64x5 FILLER_236_1110 ();
 b15zdnd11an1n32x5 FILLER_236_1174 ();
 b15zdnd11an1n16x5 FILLER_236_1206 ();
 b15zdnd11an1n08x5 FILLER_236_1222 ();
 b15zdnd00an1n02x5 FILLER_236_1230 ();
 b15zdnd11an1n64x5 FILLER_236_1277 ();
 b15zdnd11an1n64x5 FILLER_236_1341 ();
 b15zdnd11an1n64x5 FILLER_236_1405 ();
 b15zdnd11an1n64x5 FILLER_236_1469 ();
 b15zdnd11an1n64x5 FILLER_236_1533 ();
 b15zdnd11an1n64x5 FILLER_236_1597 ();
 b15zdnd11an1n64x5 FILLER_236_1661 ();
 b15zdnd11an1n64x5 FILLER_236_1725 ();
 b15zdnd11an1n64x5 FILLER_236_1789 ();
 b15zdnd11an1n64x5 FILLER_236_1853 ();
 b15zdnd11an1n64x5 FILLER_236_1917 ();
 b15zdnd11an1n64x5 FILLER_236_1981 ();
 b15zdnd11an1n64x5 FILLER_236_2045 ();
 b15zdnd11an1n32x5 FILLER_236_2109 ();
 b15zdnd11an1n08x5 FILLER_236_2141 ();
 b15zdnd11an1n04x5 FILLER_236_2149 ();
 b15zdnd00an1n01x5 FILLER_236_2153 ();
 b15zdnd11an1n64x5 FILLER_236_2162 ();
 b15zdnd11an1n32x5 FILLER_236_2226 ();
 b15zdnd11an1n16x5 FILLER_236_2258 ();
 b15zdnd00an1n02x5 FILLER_236_2274 ();
 b15zdnd11an1n64x5 FILLER_237_0 ();
 b15zdnd11an1n64x5 FILLER_237_64 ();
 b15zdnd11an1n64x5 FILLER_237_128 ();
 b15zdnd11an1n64x5 FILLER_237_192 ();
 b15zdnd11an1n64x5 FILLER_237_256 ();
 b15zdnd11an1n64x5 FILLER_237_320 ();
 b15zdnd11an1n64x5 FILLER_237_384 ();
 b15zdnd11an1n64x5 FILLER_237_448 ();
 b15zdnd11an1n64x5 FILLER_237_512 ();
 b15zdnd11an1n64x5 FILLER_237_576 ();
 b15zdnd11an1n64x5 FILLER_237_640 ();
 b15zdnd11an1n64x5 FILLER_237_704 ();
 b15zdnd11an1n64x5 FILLER_237_768 ();
 b15zdnd11an1n64x5 FILLER_237_832 ();
 b15zdnd11an1n64x5 FILLER_237_896 ();
 b15zdnd11an1n64x5 FILLER_237_960 ();
 b15zdnd11an1n64x5 FILLER_237_1024 ();
 b15zdnd11an1n64x5 FILLER_237_1088 ();
 b15zdnd11an1n64x5 FILLER_237_1152 ();
 b15zdnd11an1n08x5 FILLER_237_1216 ();
 b15zdnd11an1n04x5 FILLER_237_1224 ();
 b15zdnd11an1n04x5 FILLER_237_1245 ();
 b15zdnd11an1n64x5 FILLER_237_1263 ();
 b15zdnd11an1n64x5 FILLER_237_1327 ();
 b15zdnd11an1n64x5 FILLER_237_1391 ();
 b15zdnd11an1n64x5 FILLER_237_1455 ();
 b15zdnd11an1n64x5 FILLER_237_1519 ();
 b15zdnd11an1n64x5 FILLER_237_1583 ();
 b15zdnd11an1n64x5 FILLER_237_1647 ();
 b15zdnd11an1n64x5 FILLER_237_1711 ();
 b15zdnd11an1n64x5 FILLER_237_1775 ();
 b15zdnd11an1n64x5 FILLER_237_1839 ();
 b15zdnd11an1n64x5 FILLER_237_1903 ();
 b15zdnd11an1n64x5 FILLER_237_1967 ();
 b15zdnd11an1n64x5 FILLER_237_2031 ();
 b15zdnd11an1n64x5 FILLER_237_2095 ();
 b15zdnd11an1n64x5 FILLER_237_2159 ();
 b15zdnd11an1n32x5 FILLER_237_2223 ();
 b15zdnd11an1n16x5 FILLER_237_2255 ();
 b15zdnd11an1n08x5 FILLER_237_2271 ();
 b15zdnd11an1n04x5 FILLER_237_2279 ();
 b15zdnd00an1n01x5 FILLER_237_2283 ();
 b15zdnd11an1n64x5 FILLER_238_8 ();
 b15zdnd11an1n64x5 FILLER_238_72 ();
 b15zdnd11an1n64x5 FILLER_238_136 ();
 b15zdnd11an1n64x5 FILLER_238_200 ();
 b15zdnd11an1n64x5 FILLER_238_264 ();
 b15zdnd11an1n64x5 FILLER_238_328 ();
 b15zdnd11an1n64x5 FILLER_238_392 ();
 b15zdnd11an1n64x5 FILLER_238_456 ();
 b15zdnd11an1n64x5 FILLER_238_520 ();
 b15zdnd11an1n64x5 FILLER_238_584 ();
 b15zdnd11an1n64x5 FILLER_238_648 ();
 b15zdnd11an1n04x5 FILLER_238_712 ();
 b15zdnd00an1n02x5 FILLER_238_716 ();
 b15zdnd11an1n64x5 FILLER_238_726 ();
 b15zdnd11an1n64x5 FILLER_238_790 ();
 b15zdnd11an1n64x5 FILLER_238_854 ();
 b15zdnd11an1n64x5 FILLER_238_918 ();
 b15zdnd11an1n64x5 FILLER_238_982 ();
 b15zdnd11an1n64x5 FILLER_238_1046 ();
 b15zdnd11an1n16x5 FILLER_238_1110 ();
 b15zdnd11an1n08x5 FILLER_238_1126 ();
 b15zdnd11an1n04x5 FILLER_238_1134 ();
 b15zdnd00an1n02x5 FILLER_238_1138 ();
 b15zdnd00an1n01x5 FILLER_238_1140 ();
 b15zdnd11an1n64x5 FILLER_238_1157 ();
 b15zdnd11an1n64x5 FILLER_238_1221 ();
 b15zdnd11an1n64x5 FILLER_238_1285 ();
 b15zdnd11an1n64x5 FILLER_238_1349 ();
 b15zdnd11an1n64x5 FILLER_238_1413 ();
 b15zdnd11an1n64x5 FILLER_238_1477 ();
 b15zdnd11an1n64x5 FILLER_238_1541 ();
 b15zdnd11an1n64x5 FILLER_238_1605 ();
 b15zdnd11an1n64x5 FILLER_238_1669 ();
 b15zdnd11an1n64x5 FILLER_238_1733 ();
 b15zdnd11an1n64x5 FILLER_238_1797 ();
 b15zdnd11an1n64x5 FILLER_238_1861 ();
 b15zdnd11an1n64x5 FILLER_238_1925 ();
 b15zdnd11an1n64x5 FILLER_238_1989 ();
 b15zdnd11an1n64x5 FILLER_238_2053 ();
 b15zdnd11an1n32x5 FILLER_238_2117 ();
 b15zdnd11an1n04x5 FILLER_238_2149 ();
 b15zdnd00an1n01x5 FILLER_238_2153 ();
 b15zdnd11an1n64x5 FILLER_238_2162 ();
 b15zdnd11an1n32x5 FILLER_238_2226 ();
 b15zdnd11an1n16x5 FILLER_238_2258 ();
 b15zdnd00an1n02x5 FILLER_238_2274 ();
 b15zdnd11an1n64x5 FILLER_239_0 ();
 b15zdnd11an1n64x5 FILLER_239_64 ();
 b15zdnd11an1n64x5 FILLER_239_128 ();
 b15zdnd11an1n64x5 FILLER_239_192 ();
 b15zdnd11an1n64x5 FILLER_239_256 ();
 b15zdnd11an1n64x5 FILLER_239_320 ();
 b15zdnd11an1n64x5 FILLER_239_384 ();
 b15zdnd11an1n64x5 FILLER_239_448 ();
 b15zdnd11an1n64x5 FILLER_239_512 ();
 b15zdnd11an1n64x5 FILLER_239_576 ();
 b15zdnd11an1n64x5 FILLER_239_640 ();
 b15zdnd11an1n64x5 FILLER_239_704 ();
 b15zdnd11an1n64x5 FILLER_239_768 ();
 b15zdnd11an1n64x5 FILLER_239_832 ();
 b15zdnd11an1n64x5 FILLER_239_896 ();
 b15zdnd11an1n64x5 FILLER_239_960 ();
 b15zdnd11an1n64x5 FILLER_239_1024 ();
 b15zdnd11an1n64x5 FILLER_239_1088 ();
 b15zdnd11an1n64x5 FILLER_239_1152 ();
 b15zdnd11an1n64x5 FILLER_239_1216 ();
 b15zdnd11an1n64x5 FILLER_239_1280 ();
 b15zdnd11an1n64x5 FILLER_239_1344 ();
 b15zdnd11an1n64x5 FILLER_239_1408 ();
 b15zdnd11an1n64x5 FILLER_239_1472 ();
 b15zdnd11an1n64x5 FILLER_239_1536 ();
 b15zdnd11an1n64x5 FILLER_239_1600 ();
 b15zdnd11an1n64x5 FILLER_239_1664 ();
 b15zdnd11an1n64x5 FILLER_239_1728 ();
 b15zdnd11an1n64x5 FILLER_239_1792 ();
 b15zdnd11an1n64x5 FILLER_239_1856 ();
 b15zdnd11an1n64x5 FILLER_239_1920 ();
 b15zdnd11an1n64x5 FILLER_239_1984 ();
 b15zdnd11an1n64x5 FILLER_239_2048 ();
 b15zdnd11an1n64x5 FILLER_239_2112 ();
 b15zdnd11an1n64x5 FILLER_239_2176 ();
 b15zdnd11an1n32x5 FILLER_239_2240 ();
 b15zdnd11an1n08x5 FILLER_239_2272 ();
 b15zdnd11an1n04x5 FILLER_239_2280 ();
 b15zdnd11an1n64x5 FILLER_240_8 ();
 b15zdnd11an1n64x5 FILLER_240_72 ();
 b15zdnd11an1n64x5 FILLER_240_136 ();
 b15zdnd11an1n64x5 FILLER_240_200 ();
 b15zdnd11an1n64x5 FILLER_240_264 ();
 b15zdnd11an1n64x5 FILLER_240_328 ();
 b15zdnd11an1n64x5 FILLER_240_392 ();
 b15zdnd11an1n64x5 FILLER_240_456 ();
 b15zdnd11an1n64x5 FILLER_240_520 ();
 b15zdnd11an1n32x5 FILLER_240_584 ();
 b15zdnd11an1n16x5 FILLER_240_616 ();
 b15zdnd11an1n08x5 FILLER_240_632 ();
 b15zdnd00an1n01x5 FILLER_240_640 ();
 b15zdnd11an1n64x5 FILLER_240_652 ();
 b15zdnd00an1n02x5 FILLER_240_716 ();
 b15zdnd11an1n64x5 FILLER_240_726 ();
 b15zdnd11an1n64x5 FILLER_240_790 ();
 b15zdnd11an1n64x5 FILLER_240_854 ();
 b15zdnd11an1n64x5 FILLER_240_918 ();
 b15zdnd11an1n64x5 FILLER_240_982 ();
 b15zdnd11an1n64x5 FILLER_240_1046 ();
 b15zdnd11an1n64x5 FILLER_240_1110 ();
 b15zdnd11an1n64x5 FILLER_240_1174 ();
 b15zdnd11an1n64x5 FILLER_240_1238 ();
 b15zdnd11an1n64x5 FILLER_240_1302 ();
 b15zdnd11an1n64x5 FILLER_240_1366 ();
 b15zdnd11an1n64x5 FILLER_240_1430 ();
 b15zdnd11an1n64x5 FILLER_240_1494 ();
 b15zdnd11an1n64x5 FILLER_240_1558 ();
 b15zdnd11an1n64x5 FILLER_240_1622 ();
 b15zdnd11an1n64x5 FILLER_240_1686 ();
 b15zdnd11an1n64x5 FILLER_240_1750 ();
 b15zdnd11an1n64x5 FILLER_240_1814 ();
 b15zdnd11an1n64x5 FILLER_240_1878 ();
 b15zdnd11an1n64x5 FILLER_240_1942 ();
 b15zdnd11an1n64x5 FILLER_240_2006 ();
 b15zdnd11an1n64x5 FILLER_240_2070 ();
 b15zdnd11an1n16x5 FILLER_240_2134 ();
 b15zdnd11an1n04x5 FILLER_240_2150 ();
 b15zdnd11an1n64x5 FILLER_240_2162 ();
 b15zdnd11an1n32x5 FILLER_240_2226 ();
 b15zdnd11an1n16x5 FILLER_240_2258 ();
 b15zdnd00an1n02x5 FILLER_240_2274 ();
 b15zdnd11an1n64x5 FILLER_241_0 ();
 b15zdnd11an1n64x5 FILLER_241_64 ();
 b15zdnd11an1n64x5 FILLER_241_128 ();
 b15zdnd11an1n64x5 FILLER_241_192 ();
 b15zdnd11an1n64x5 FILLER_241_256 ();
 b15zdnd11an1n64x5 FILLER_241_320 ();
 b15zdnd11an1n64x5 FILLER_241_384 ();
 b15zdnd11an1n64x5 FILLER_241_448 ();
 b15zdnd11an1n64x5 FILLER_241_512 ();
 b15zdnd11an1n64x5 FILLER_241_576 ();
 b15zdnd11an1n64x5 FILLER_241_640 ();
 b15zdnd11an1n64x5 FILLER_241_704 ();
 b15zdnd11an1n64x5 FILLER_241_768 ();
 b15zdnd11an1n64x5 FILLER_241_832 ();
 b15zdnd11an1n64x5 FILLER_241_896 ();
 b15zdnd11an1n64x5 FILLER_241_960 ();
 b15zdnd11an1n64x5 FILLER_241_1024 ();
 b15zdnd11an1n64x5 FILLER_241_1088 ();
 b15zdnd11an1n64x5 FILLER_241_1152 ();
 b15zdnd11an1n64x5 FILLER_241_1216 ();
 b15zdnd11an1n64x5 FILLER_241_1280 ();
 b15zdnd11an1n64x5 FILLER_241_1344 ();
 b15zdnd11an1n64x5 FILLER_241_1408 ();
 b15zdnd11an1n64x5 FILLER_241_1472 ();
 b15zdnd11an1n64x5 FILLER_241_1536 ();
 b15zdnd11an1n64x5 FILLER_241_1600 ();
 b15zdnd11an1n64x5 FILLER_241_1664 ();
 b15zdnd11an1n64x5 FILLER_241_1728 ();
 b15zdnd11an1n64x5 FILLER_241_1792 ();
 b15zdnd11an1n64x5 FILLER_241_1856 ();
 b15zdnd11an1n64x5 FILLER_241_1920 ();
 b15zdnd11an1n64x5 FILLER_241_1984 ();
 b15zdnd11an1n64x5 FILLER_241_2048 ();
 b15zdnd11an1n64x5 FILLER_241_2112 ();
 b15zdnd11an1n64x5 FILLER_241_2176 ();
 b15zdnd11an1n32x5 FILLER_241_2240 ();
 b15zdnd11an1n08x5 FILLER_241_2272 ();
 b15zdnd11an1n04x5 FILLER_241_2280 ();
 b15zdnd11an1n64x5 FILLER_242_8 ();
 b15zdnd11an1n64x5 FILLER_242_72 ();
 b15zdnd11an1n64x5 FILLER_242_136 ();
 b15zdnd11an1n64x5 FILLER_242_200 ();
 b15zdnd11an1n64x5 FILLER_242_264 ();
 b15zdnd11an1n64x5 FILLER_242_328 ();
 b15zdnd11an1n64x5 FILLER_242_392 ();
 b15zdnd11an1n64x5 FILLER_242_456 ();
 b15zdnd11an1n64x5 FILLER_242_520 ();
 b15zdnd11an1n64x5 FILLER_242_584 ();
 b15zdnd11an1n64x5 FILLER_242_648 ();
 b15zdnd11an1n04x5 FILLER_242_712 ();
 b15zdnd00an1n02x5 FILLER_242_716 ();
 b15zdnd11an1n64x5 FILLER_242_726 ();
 b15zdnd11an1n64x5 FILLER_242_790 ();
 b15zdnd11an1n64x5 FILLER_242_854 ();
 b15zdnd11an1n64x5 FILLER_242_918 ();
 b15zdnd11an1n32x5 FILLER_242_982 ();
 b15zdnd11an1n16x5 FILLER_242_1014 ();
 b15zdnd11an1n08x5 FILLER_242_1030 ();
 b15zdnd11an1n04x5 FILLER_242_1038 ();
 b15zdnd11an1n64x5 FILLER_242_1058 ();
 b15zdnd11an1n64x5 FILLER_242_1122 ();
 b15zdnd11an1n64x5 FILLER_242_1186 ();
 b15zdnd11an1n64x5 FILLER_242_1250 ();
 b15zdnd11an1n64x5 FILLER_242_1314 ();
 b15zdnd11an1n64x5 FILLER_242_1378 ();
 b15zdnd11an1n64x5 FILLER_242_1442 ();
 b15zdnd11an1n64x5 FILLER_242_1506 ();
 b15zdnd11an1n64x5 FILLER_242_1570 ();
 b15zdnd11an1n64x5 FILLER_242_1634 ();
 b15zdnd11an1n64x5 FILLER_242_1698 ();
 b15zdnd11an1n64x5 FILLER_242_1762 ();
 b15zdnd11an1n64x5 FILLER_242_1826 ();
 b15zdnd11an1n64x5 FILLER_242_1890 ();
 b15zdnd11an1n64x5 FILLER_242_1954 ();
 b15zdnd11an1n64x5 FILLER_242_2018 ();
 b15zdnd11an1n64x5 FILLER_242_2082 ();
 b15zdnd11an1n08x5 FILLER_242_2146 ();
 b15zdnd11an1n64x5 FILLER_242_2162 ();
 b15zdnd11an1n32x5 FILLER_242_2226 ();
 b15zdnd11an1n16x5 FILLER_242_2258 ();
 b15zdnd00an1n02x5 FILLER_242_2274 ();
 b15zdnd11an1n64x5 FILLER_243_0 ();
 b15zdnd11an1n64x5 FILLER_243_64 ();
 b15zdnd11an1n64x5 FILLER_243_128 ();
 b15zdnd11an1n64x5 FILLER_243_192 ();
 b15zdnd11an1n64x5 FILLER_243_256 ();
 b15zdnd11an1n64x5 FILLER_243_320 ();
 b15zdnd11an1n64x5 FILLER_243_384 ();
 b15zdnd11an1n64x5 FILLER_243_448 ();
 b15zdnd11an1n64x5 FILLER_243_512 ();
 b15zdnd11an1n64x5 FILLER_243_576 ();
 b15zdnd11an1n64x5 FILLER_243_640 ();
 b15zdnd11an1n64x5 FILLER_243_704 ();
 b15zdnd11an1n64x5 FILLER_243_768 ();
 b15zdnd11an1n64x5 FILLER_243_832 ();
 b15zdnd11an1n32x5 FILLER_243_896 ();
 b15zdnd11an1n08x5 FILLER_243_928 ();
 b15zdnd11an1n04x5 FILLER_243_936 ();
 b15zdnd00an1n02x5 FILLER_243_940 ();
 b15zdnd11an1n64x5 FILLER_243_958 ();
 b15zdnd11an1n64x5 FILLER_243_1022 ();
 b15zdnd11an1n64x5 FILLER_243_1086 ();
 b15zdnd11an1n64x5 FILLER_243_1150 ();
 b15zdnd11an1n64x5 FILLER_243_1214 ();
 b15zdnd11an1n64x5 FILLER_243_1278 ();
 b15zdnd11an1n64x5 FILLER_243_1342 ();
 b15zdnd11an1n64x5 FILLER_243_1406 ();
 b15zdnd11an1n64x5 FILLER_243_1470 ();
 b15zdnd11an1n64x5 FILLER_243_1534 ();
 b15zdnd11an1n64x5 FILLER_243_1598 ();
 b15zdnd11an1n64x5 FILLER_243_1662 ();
 b15zdnd11an1n64x5 FILLER_243_1726 ();
 b15zdnd11an1n64x5 FILLER_243_1790 ();
 b15zdnd11an1n64x5 FILLER_243_1854 ();
 b15zdnd11an1n64x5 FILLER_243_1918 ();
 b15zdnd11an1n64x5 FILLER_243_1982 ();
 b15zdnd11an1n64x5 FILLER_243_2046 ();
 b15zdnd11an1n64x5 FILLER_243_2110 ();
 b15zdnd11an1n64x5 FILLER_243_2174 ();
 b15zdnd11an1n32x5 FILLER_243_2238 ();
 b15zdnd11an1n08x5 FILLER_243_2270 ();
 b15zdnd11an1n04x5 FILLER_243_2278 ();
 b15zdnd00an1n02x5 FILLER_243_2282 ();
 b15zdnd11an1n64x5 FILLER_244_8 ();
 b15zdnd11an1n64x5 FILLER_244_72 ();
 b15zdnd11an1n64x5 FILLER_244_136 ();
 b15zdnd11an1n64x5 FILLER_244_200 ();
 b15zdnd11an1n64x5 FILLER_244_264 ();
 b15zdnd11an1n64x5 FILLER_244_328 ();
 b15zdnd11an1n64x5 FILLER_244_392 ();
 b15zdnd11an1n64x5 FILLER_244_456 ();
 b15zdnd11an1n64x5 FILLER_244_520 ();
 b15zdnd11an1n64x5 FILLER_244_584 ();
 b15zdnd11an1n64x5 FILLER_244_648 ();
 b15zdnd11an1n04x5 FILLER_244_712 ();
 b15zdnd00an1n02x5 FILLER_244_716 ();
 b15zdnd11an1n64x5 FILLER_244_726 ();
 b15zdnd11an1n64x5 FILLER_244_790 ();
 b15zdnd11an1n64x5 FILLER_244_854 ();
 b15zdnd11an1n64x5 FILLER_244_918 ();
 b15zdnd11an1n64x5 FILLER_244_982 ();
 b15zdnd11an1n64x5 FILLER_244_1046 ();
 b15zdnd11an1n64x5 FILLER_244_1110 ();
 b15zdnd11an1n64x5 FILLER_244_1174 ();
 b15zdnd11an1n64x5 FILLER_244_1238 ();
 b15zdnd11an1n64x5 FILLER_244_1302 ();
 b15zdnd11an1n64x5 FILLER_244_1366 ();
 b15zdnd11an1n64x5 FILLER_244_1430 ();
 b15zdnd11an1n64x5 FILLER_244_1494 ();
 b15zdnd11an1n64x5 FILLER_244_1558 ();
 b15zdnd11an1n64x5 FILLER_244_1622 ();
 b15zdnd11an1n64x5 FILLER_244_1686 ();
 b15zdnd11an1n64x5 FILLER_244_1750 ();
 b15zdnd11an1n64x5 FILLER_244_1814 ();
 b15zdnd11an1n64x5 FILLER_244_1878 ();
 b15zdnd11an1n64x5 FILLER_244_1942 ();
 b15zdnd11an1n64x5 FILLER_244_2006 ();
 b15zdnd11an1n64x5 FILLER_244_2070 ();
 b15zdnd11an1n16x5 FILLER_244_2134 ();
 b15zdnd11an1n04x5 FILLER_244_2150 ();
 b15zdnd11an1n64x5 FILLER_244_2162 ();
 b15zdnd11an1n32x5 FILLER_244_2226 ();
 b15zdnd11an1n16x5 FILLER_244_2258 ();
 b15zdnd00an1n02x5 FILLER_244_2274 ();
 b15zdnd11an1n64x5 FILLER_245_0 ();
 b15zdnd11an1n64x5 FILLER_245_64 ();
 b15zdnd11an1n64x5 FILLER_245_128 ();
 b15zdnd11an1n64x5 FILLER_245_192 ();
 b15zdnd11an1n64x5 FILLER_245_256 ();
 b15zdnd11an1n64x5 FILLER_245_320 ();
 b15zdnd11an1n64x5 FILLER_245_384 ();
 b15zdnd11an1n64x5 FILLER_245_448 ();
 b15zdnd11an1n64x5 FILLER_245_512 ();
 b15zdnd11an1n64x5 FILLER_245_576 ();
 b15zdnd11an1n64x5 FILLER_245_640 ();
 b15zdnd11an1n64x5 FILLER_245_704 ();
 b15zdnd11an1n64x5 FILLER_245_768 ();
 b15zdnd11an1n64x5 FILLER_245_832 ();
 b15zdnd11an1n64x5 FILLER_245_896 ();
 b15zdnd11an1n64x5 FILLER_245_960 ();
 b15zdnd11an1n16x5 FILLER_245_1024 ();
 b15zdnd11an1n08x5 FILLER_245_1040 ();
 b15zdnd00an1n02x5 FILLER_245_1048 ();
 b15zdnd11an1n64x5 FILLER_245_1092 ();
 b15zdnd11an1n64x5 FILLER_245_1156 ();
 b15zdnd11an1n64x5 FILLER_245_1220 ();
 b15zdnd11an1n64x5 FILLER_245_1284 ();
 b15zdnd11an1n64x5 FILLER_245_1348 ();
 b15zdnd11an1n64x5 FILLER_245_1412 ();
 b15zdnd11an1n64x5 FILLER_245_1476 ();
 b15zdnd11an1n64x5 FILLER_245_1540 ();
 b15zdnd11an1n64x5 FILLER_245_1604 ();
 b15zdnd11an1n64x5 FILLER_245_1668 ();
 b15zdnd11an1n64x5 FILLER_245_1732 ();
 b15zdnd11an1n64x5 FILLER_245_1796 ();
 b15zdnd11an1n64x5 FILLER_245_1860 ();
 b15zdnd11an1n64x5 FILLER_245_1924 ();
 b15zdnd11an1n64x5 FILLER_245_1988 ();
 b15zdnd11an1n64x5 FILLER_245_2052 ();
 b15zdnd11an1n64x5 FILLER_245_2116 ();
 b15zdnd11an1n64x5 FILLER_245_2180 ();
 b15zdnd11an1n32x5 FILLER_245_2244 ();
 b15zdnd11an1n08x5 FILLER_245_2276 ();
 b15zdnd11an1n64x5 FILLER_246_8 ();
 b15zdnd11an1n64x5 FILLER_246_72 ();
 b15zdnd11an1n64x5 FILLER_246_136 ();
 b15zdnd11an1n64x5 FILLER_246_200 ();
 b15zdnd11an1n64x5 FILLER_246_264 ();
 b15zdnd11an1n64x5 FILLER_246_328 ();
 b15zdnd11an1n64x5 FILLER_246_392 ();
 b15zdnd11an1n64x5 FILLER_246_456 ();
 b15zdnd11an1n64x5 FILLER_246_520 ();
 b15zdnd11an1n64x5 FILLER_246_584 ();
 b15zdnd11an1n64x5 FILLER_246_648 ();
 b15zdnd11an1n04x5 FILLER_246_712 ();
 b15zdnd00an1n02x5 FILLER_246_716 ();
 b15zdnd11an1n64x5 FILLER_246_726 ();
 b15zdnd11an1n64x5 FILLER_246_790 ();
 b15zdnd11an1n64x5 FILLER_246_854 ();
 b15zdnd11an1n64x5 FILLER_246_918 ();
 b15zdnd11an1n64x5 FILLER_246_982 ();
 b15zdnd11an1n64x5 FILLER_246_1046 ();
 b15zdnd11an1n64x5 FILLER_246_1110 ();
 b15zdnd11an1n64x5 FILLER_246_1174 ();
 b15zdnd11an1n64x5 FILLER_246_1238 ();
 b15zdnd11an1n64x5 FILLER_246_1302 ();
 b15zdnd11an1n64x5 FILLER_246_1366 ();
 b15zdnd11an1n64x5 FILLER_246_1430 ();
 b15zdnd11an1n64x5 FILLER_246_1494 ();
 b15zdnd11an1n64x5 FILLER_246_1558 ();
 b15zdnd11an1n64x5 FILLER_246_1622 ();
 b15zdnd11an1n64x5 FILLER_246_1686 ();
 b15zdnd11an1n64x5 FILLER_246_1750 ();
 b15zdnd11an1n64x5 FILLER_246_1814 ();
 b15zdnd11an1n64x5 FILLER_246_1878 ();
 b15zdnd11an1n64x5 FILLER_246_1942 ();
 b15zdnd11an1n64x5 FILLER_246_2006 ();
 b15zdnd11an1n64x5 FILLER_246_2070 ();
 b15zdnd11an1n16x5 FILLER_246_2134 ();
 b15zdnd11an1n04x5 FILLER_246_2150 ();
 b15zdnd11an1n64x5 FILLER_246_2162 ();
 b15zdnd11an1n32x5 FILLER_246_2226 ();
 b15zdnd11an1n16x5 FILLER_246_2258 ();
 b15zdnd00an1n02x5 FILLER_246_2274 ();
 b15zdnd11an1n64x5 FILLER_247_0 ();
 b15zdnd11an1n64x5 FILLER_247_64 ();
 b15zdnd11an1n64x5 FILLER_247_128 ();
 b15zdnd11an1n64x5 FILLER_247_192 ();
 b15zdnd11an1n64x5 FILLER_247_256 ();
 b15zdnd11an1n64x5 FILLER_247_320 ();
 b15zdnd11an1n64x5 FILLER_247_384 ();
 b15zdnd11an1n64x5 FILLER_247_448 ();
 b15zdnd11an1n64x5 FILLER_247_512 ();
 b15zdnd11an1n64x5 FILLER_247_576 ();
 b15zdnd11an1n64x5 FILLER_247_640 ();
 b15zdnd11an1n64x5 FILLER_247_704 ();
 b15zdnd11an1n64x5 FILLER_247_768 ();
 b15zdnd11an1n64x5 FILLER_247_832 ();
 b15zdnd11an1n64x5 FILLER_247_896 ();
 b15zdnd11an1n64x5 FILLER_247_960 ();
 b15zdnd11an1n64x5 FILLER_247_1024 ();
 b15zdnd11an1n64x5 FILLER_247_1088 ();
 b15zdnd11an1n64x5 FILLER_247_1152 ();
 b15zdnd11an1n64x5 FILLER_247_1216 ();
 b15zdnd11an1n64x5 FILLER_247_1280 ();
 b15zdnd11an1n64x5 FILLER_247_1344 ();
 b15zdnd11an1n64x5 FILLER_247_1408 ();
 b15zdnd11an1n64x5 FILLER_247_1472 ();
 b15zdnd11an1n64x5 FILLER_247_1536 ();
 b15zdnd11an1n64x5 FILLER_247_1600 ();
 b15zdnd11an1n64x5 FILLER_247_1664 ();
 b15zdnd11an1n64x5 FILLER_247_1728 ();
 b15zdnd11an1n64x5 FILLER_247_1792 ();
 b15zdnd11an1n64x5 FILLER_247_1856 ();
 b15zdnd11an1n64x5 FILLER_247_1920 ();
 b15zdnd11an1n64x5 FILLER_247_1984 ();
 b15zdnd11an1n64x5 FILLER_247_2048 ();
 b15zdnd11an1n64x5 FILLER_247_2112 ();
 b15zdnd11an1n64x5 FILLER_247_2176 ();
 b15zdnd11an1n32x5 FILLER_247_2240 ();
 b15zdnd11an1n08x5 FILLER_247_2272 ();
 b15zdnd11an1n04x5 FILLER_247_2280 ();
 b15zdnd11an1n64x5 FILLER_248_8 ();
 b15zdnd11an1n64x5 FILLER_248_72 ();
 b15zdnd11an1n64x5 FILLER_248_136 ();
 b15zdnd11an1n64x5 FILLER_248_200 ();
 b15zdnd11an1n64x5 FILLER_248_264 ();
 b15zdnd11an1n64x5 FILLER_248_328 ();
 b15zdnd11an1n64x5 FILLER_248_392 ();
 b15zdnd11an1n64x5 FILLER_248_456 ();
 b15zdnd11an1n64x5 FILLER_248_520 ();
 b15zdnd11an1n64x5 FILLER_248_584 ();
 b15zdnd11an1n64x5 FILLER_248_648 ();
 b15zdnd11an1n04x5 FILLER_248_712 ();
 b15zdnd00an1n02x5 FILLER_248_716 ();
 b15zdnd11an1n64x5 FILLER_248_726 ();
 b15zdnd11an1n64x5 FILLER_248_790 ();
 b15zdnd11an1n64x5 FILLER_248_854 ();
 b15zdnd11an1n64x5 FILLER_248_918 ();
 b15zdnd11an1n64x5 FILLER_248_982 ();
 b15zdnd11an1n64x5 FILLER_248_1046 ();
 b15zdnd11an1n64x5 FILLER_248_1110 ();
 b15zdnd11an1n64x5 FILLER_248_1174 ();
 b15zdnd11an1n64x5 FILLER_248_1238 ();
 b15zdnd11an1n64x5 FILLER_248_1302 ();
 b15zdnd11an1n64x5 FILLER_248_1366 ();
 b15zdnd11an1n64x5 FILLER_248_1430 ();
 b15zdnd11an1n64x5 FILLER_248_1494 ();
 b15zdnd11an1n64x5 FILLER_248_1558 ();
 b15zdnd11an1n64x5 FILLER_248_1622 ();
 b15zdnd11an1n64x5 FILLER_248_1686 ();
 b15zdnd11an1n64x5 FILLER_248_1750 ();
 b15zdnd11an1n64x5 FILLER_248_1814 ();
 b15zdnd11an1n64x5 FILLER_248_1878 ();
 b15zdnd11an1n64x5 FILLER_248_1942 ();
 b15zdnd11an1n64x5 FILLER_248_2006 ();
 b15zdnd11an1n64x5 FILLER_248_2070 ();
 b15zdnd11an1n16x5 FILLER_248_2134 ();
 b15zdnd11an1n04x5 FILLER_248_2150 ();
 b15zdnd11an1n64x5 FILLER_248_2162 ();
 b15zdnd11an1n32x5 FILLER_248_2226 ();
 b15zdnd11an1n16x5 FILLER_248_2258 ();
 b15zdnd00an1n02x5 FILLER_248_2274 ();
 b15zdnd11an1n64x5 FILLER_249_0 ();
 b15zdnd11an1n64x5 FILLER_249_64 ();
 b15zdnd11an1n64x5 FILLER_249_128 ();
 b15zdnd11an1n64x5 FILLER_249_192 ();
 b15zdnd11an1n64x5 FILLER_249_256 ();
 b15zdnd11an1n64x5 FILLER_249_320 ();
 b15zdnd11an1n64x5 FILLER_249_384 ();
 b15zdnd11an1n64x5 FILLER_249_448 ();
 b15zdnd11an1n64x5 FILLER_249_512 ();
 b15zdnd11an1n64x5 FILLER_249_576 ();
 b15zdnd11an1n64x5 FILLER_249_640 ();
 b15zdnd11an1n64x5 FILLER_249_704 ();
 b15zdnd11an1n64x5 FILLER_249_768 ();
 b15zdnd11an1n64x5 FILLER_249_832 ();
 b15zdnd11an1n64x5 FILLER_249_896 ();
 b15zdnd11an1n64x5 FILLER_249_960 ();
 b15zdnd11an1n64x5 FILLER_249_1024 ();
 b15zdnd11an1n64x5 FILLER_249_1088 ();
 b15zdnd11an1n64x5 FILLER_249_1152 ();
 b15zdnd11an1n64x5 FILLER_249_1216 ();
 b15zdnd11an1n64x5 FILLER_249_1280 ();
 b15zdnd11an1n64x5 FILLER_249_1344 ();
 b15zdnd11an1n64x5 FILLER_249_1408 ();
 b15zdnd11an1n64x5 FILLER_249_1472 ();
 b15zdnd11an1n64x5 FILLER_249_1536 ();
 b15zdnd11an1n64x5 FILLER_249_1600 ();
 b15zdnd11an1n64x5 FILLER_249_1664 ();
 b15zdnd11an1n64x5 FILLER_249_1728 ();
 b15zdnd11an1n64x5 FILLER_249_1792 ();
 b15zdnd11an1n64x5 FILLER_249_1856 ();
 b15zdnd11an1n64x5 FILLER_249_1920 ();
 b15zdnd11an1n64x5 FILLER_249_1984 ();
 b15zdnd11an1n64x5 FILLER_249_2048 ();
 b15zdnd11an1n64x5 FILLER_249_2112 ();
 b15zdnd11an1n64x5 FILLER_249_2176 ();
 b15zdnd11an1n32x5 FILLER_249_2240 ();
 b15zdnd11an1n08x5 FILLER_249_2272 ();
 b15zdnd11an1n04x5 FILLER_249_2280 ();
 b15zdnd11an1n64x5 FILLER_250_8 ();
 b15zdnd11an1n64x5 FILLER_250_72 ();
 b15zdnd11an1n64x5 FILLER_250_136 ();
 b15zdnd11an1n64x5 FILLER_250_200 ();
 b15zdnd11an1n64x5 FILLER_250_264 ();
 b15zdnd11an1n64x5 FILLER_250_328 ();
 b15zdnd11an1n64x5 FILLER_250_392 ();
 b15zdnd11an1n64x5 FILLER_250_456 ();
 b15zdnd11an1n64x5 FILLER_250_520 ();
 b15zdnd11an1n64x5 FILLER_250_584 ();
 b15zdnd11an1n64x5 FILLER_250_648 ();
 b15zdnd11an1n04x5 FILLER_250_712 ();
 b15zdnd00an1n02x5 FILLER_250_716 ();
 b15zdnd11an1n64x5 FILLER_250_726 ();
 b15zdnd11an1n64x5 FILLER_250_790 ();
 b15zdnd11an1n64x5 FILLER_250_854 ();
 b15zdnd11an1n64x5 FILLER_250_918 ();
 b15zdnd11an1n64x5 FILLER_250_982 ();
 b15zdnd11an1n64x5 FILLER_250_1046 ();
 b15zdnd11an1n64x5 FILLER_250_1110 ();
 b15zdnd11an1n64x5 FILLER_250_1174 ();
 b15zdnd11an1n64x5 FILLER_250_1238 ();
 b15zdnd11an1n64x5 FILLER_250_1302 ();
 b15zdnd11an1n64x5 FILLER_250_1366 ();
 b15zdnd11an1n64x5 FILLER_250_1430 ();
 b15zdnd11an1n64x5 FILLER_250_1494 ();
 b15zdnd11an1n64x5 FILLER_250_1558 ();
 b15zdnd11an1n64x5 FILLER_250_1622 ();
 b15zdnd11an1n64x5 FILLER_250_1686 ();
 b15zdnd11an1n64x5 FILLER_250_1750 ();
 b15zdnd11an1n64x5 FILLER_250_1814 ();
 b15zdnd11an1n64x5 FILLER_250_1878 ();
 b15zdnd11an1n64x5 FILLER_250_1942 ();
 b15zdnd11an1n64x5 FILLER_250_2006 ();
 b15zdnd11an1n64x5 FILLER_250_2070 ();
 b15zdnd11an1n16x5 FILLER_250_2134 ();
 b15zdnd11an1n04x5 FILLER_250_2150 ();
 b15zdnd11an1n64x5 FILLER_250_2162 ();
 b15zdnd11an1n32x5 FILLER_250_2226 ();
 b15zdnd11an1n16x5 FILLER_250_2258 ();
 b15zdnd00an1n02x5 FILLER_250_2274 ();
 b15zdnd11an1n64x5 FILLER_251_0 ();
 b15zdnd11an1n64x5 FILLER_251_64 ();
 b15zdnd11an1n64x5 FILLER_251_128 ();
 b15zdnd11an1n64x5 FILLER_251_192 ();
 b15zdnd11an1n64x5 FILLER_251_256 ();
 b15zdnd11an1n64x5 FILLER_251_320 ();
 b15zdnd11an1n64x5 FILLER_251_384 ();
 b15zdnd11an1n64x5 FILLER_251_448 ();
 b15zdnd11an1n64x5 FILLER_251_512 ();
 b15zdnd11an1n64x5 FILLER_251_576 ();
 b15zdnd11an1n64x5 FILLER_251_640 ();
 b15zdnd11an1n64x5 FILLER_251_704 ();
 b15zdnd11an1n64x5 FILLER_251_768 ();
 b15zdnd11an1n64x5 FILLER_251_832 ();
 b15zdnd11an1n64x5 FILLER_251_896 ();
 b15zdnd11an1n64x5 FILLER_251_960 ();
 b15zdnd11an1n64x5 FILLER_251_1024 ();
 b15zdnd11an1n64x5 FILLER_251_1088 ();
 b15zdnd11an1n64x5 FILLER_251_1152 ();
 b15zdnd11an1n64x5 FILLER_251_1216 ();
 b15zdnd11an1n64x5 FILLER_251_1280 ();
 b15zdnd11an1n64x5 FILLER_251_1344 ();
 b15zdnd11an1n64x5 FILLER_251_1408 ();
 b15zdnd11an1n64x5 FILLER_251_1472 ();
 b15zdnd11an1n64x5 FILLER_251_1536 ();
 b15zdnd11an1n64x5 FILLER_251_1600 ();
 b15zdnd11an1n64x5 FILLER_251_1664 ();
 b15zdnd11an1n64x5 FILLER_251_1728 ();
 b15zdnd11an1n64x5 FILLER_251_1792 ();
 b15zdnd11an1n64x5 FILLER_251_1856 ();
 b15zdnd11an1n64x5 FILLER_251_1920 ();
 b15zdnd11an1n64x5 FILLER_251_1984 ();
 b15zdnd11an1n64x5 FILLER_251_2048 ();
 b15zdnd11an1n64x5 FILLER_251_2112 ();
 b15zdnd11an1n64x5 FILLER_251_2176 ();
 b15zdnd11an1n32x5 FILLER_251_2240 ();
 b15zdnd11an1n08x5 FILLER_251_2272 ();
 b15zdnd11an1n04x5 FILLER_251_2280 ();
 b15zdnd11an1n64x5 FILLER_252_8 ();
 b15zdnd11an1n64x5 FILLER_252_72 ();
 b15zdnd11an1n64x5 FILLER_252_136 ();
 b15zdnd11an1n64x5 FILLER_252_200 ();
 b15zdnd11an1n64x5 FILLER_252_264 ();
 b15zdnd11an1n64x5 FILLER_252_328 ();
 b15zdnd11an1n64x5 FILLER_252_392 ();
 b15zdnd11an1n64x5 FILLER_252_456 ();
 b15zdnd11an1n64x5 FILLER_252_520 ();
 b15zdnd11an1n64x5 FILLER_252_584 ();
 b15zdnd11an1n64x5 FILLER_252_648 ();
 b15zdnd11an1n04x5 FILLER_252_712 ();
 b15zdnd00an1n02x5 FILLER_252_716 ();
 b15zdnd11an1n64x5 FILLER_252_726 ();
 b15zdnd11an1n64x5 FILLER_252_790 ();
 b15zdnd11an1n64x5 FILLER_252_854 ();
 b15zdnd11an1n64x5 FILLER_252_918 ();
 b15zdnd11an1n64x5 FILLER_252_982 ();
 b15zdnd11an1n64x5 FILLER_252_1046 ();
 b15zdnd11an1n64x5 FILLER_252_1110 ();
 b15zdnd11an1n64x5 FILLER_252_1174 ();
 b15zdnd11an1n64x5 FILLER_252_1238 ();
 b15zdnd11an1n64x5 FILLER_252_1302 ();
 b15zdnd11an1n64x5 FILLER_252_1366 ();
 b15zdnd11an1n64x5 FILLER_252_1430 ();
 b15zdnd11an1n64x5 FILLER_252_1494 ();
 b15zdnd11an1n64x5 FILLER_252_1558 ();
 b15zdnd11an1n64x5 FILLER_252_1622 ();
 b15zdnd11an1n64x5 FILLER_252_1686 ();
 b15zdnd11an1n64x5 FILLER_252_1750 ();
 b15zdnd11an1n64x5 FILLER_252_1814 ();
 b15zdnd11an1n64x5 FILLER_252_1878 ();
 b15zdnd11an1n64x5 FILLER_252_1942 ();
 b15zdnd11an1n64x5 FILLER_252_2006 ();
 b15zdnd11an1n64x5 FILLER_252_2070 ();
 b15zdnd11an1n16x5 FILLER_252_2134 ();
 b15zdnd11an1n04x5 FILLER_252_2150 ();
 b15zdnd11an1n64x5 FILLER_252_2162 ();
 b15zdnd11an1n32x5 FILLER_252_2226 ();
 b15zdnd11an1n16x5 FILLER_252_2258 ();
 b15zdnd00an1n02x5 FILLER_252_2274 ();
 b15zdnd11an1n64x5 FILLER_253_0 ();
 b15zdnd11an1n64x5 FILLER_253_64 ();
 b15zdnd11an1n64x5 FILLER_253_128 ();
 b15zdnd11an1n64x5 FILLER_253_192 ();
 b15zdnd11an1n64x5 FILLER_253_256 ();
 b15zdnd11an1n64x5 FILLER_253_320 ();
 b15zdnd11an1n64x5 FILLER_253_384 ();
 b15zdnd11an1n64x5 FILLER_253_448 ();
 b15zdnd11an1n64x5 FILLER_253_512 ();
 b15zdnd11an1n64x5 FILLER_253_576 ();
 b15zdnd11an1n64x5 FILLER_253_640 ();
 b15zdnd11an1n64x5 FILLER_253_704 ();
 b15zdnd11an1n64x5 FILLER_253_768 ();
 b15zdnd11an1n64x5 FILLER_253_832 ();
 b15zdnd11an1n64x5 FILLER_253_896 ();
 b15zdnd11an1n64x5 FILLER_253_960 ();
 b15zdnd11an1n64x5 FILLER_253_1024 ();
 b15zdnd11an1n64x5 FILLER_253_1088 ();
 b15zdnd11an1n64x5 FILLER_253_1152 ();
 b15zdnd11an1n64x5 FILLER_253_1216 ();
 b15zdnd11an1n64x5 FILLER_253_1280 ();
 b15zdnd11an1n64x5 FILLER_253_1344 ();
 b15zdnd11an1n64x5 FILLER_253_1408 ();
 b15zdnd11an1n64x5 FILLER_253_1472 ();
 b15zdnd11an1n64x5 FILLER_253_1536 ();
 b15zdnd11an1n64x5 FILLER_253_1600 ();
 b15zdnd11an1n64x5 FILLER_253_1664 ();
 b15zdnd11an1n64x5 FILLER_253_1728 ();
 b15zdnd11an1n64x5 FILLER_253_1792 ();
 b15zdnd11an1n64x5 FILLER_253_1856 ();
 b15zdnd11an1n64x5 FILLER_253_1920 ();
 b15zdnd11an1n64x5 FILLER_253_1984 ();
 b15zdnd11an1n64x5 FILLER_253_2048 ();
 b15zdnd11an1n64x5 FILLER_253_2112 ();
 b15zdnd11an1n64x5 FILLER_253_2176 ();
 b15zdnd11an1n32x5 FILLER_253_2240 ();
 b15zdnd11an1n08x5 FILLER_253_2272 ();
 b15zdnd11an1n04x5 FILLER_253_2280 ();
 b15zdnd11an1n64x5 FILLER_254_8 ();
 b15zdnd11an1n64x5 FILLER_254_72 ();
 b15zdnd11an1n64x5 FILLER_254_136 ();
 b15zdnd11an1n64x5 FILLER_254_200 ();
 b15zdnd11an1n64x5 FILLER_254_264 ();
 b15zdnd11an1n64x5 FILLER_254_328 ();
 b15zdnd11an1n64x5 FILLER_254_392 ();
 b15zdnd11an1n64x5 FILLER_254_456 ();
 b15zdnd11an1n64x5 FILLER_254_520 ();
 b15zdnd11an1n64x5 FILLER_254_584 ();
 b15zdnd11an1n64x5 FILLER_254_648 ();
 b15zdnd11an1n04x5 FILLER_254_712 ();
 b15zdnd00an1n02x5 FILLER_254_716 ();
 b15zdnd11an1n64x5 FILLER_254_726 ();
 b15zdnd11an1n64x5 FILLER_254_790 ();
 b15zdnd11an1n64x5 FILLER_254_854 ();
 b15zdnd11an1n64x5 FILLER_254_918 ();
 b15zdnd11an1n64x5 FILLER_254_982 ();
 b15zdnd11an1n64x5 FILLER_254_1046 ();
 b15zdnd11an1n64x5 FILLER_254_1110 ();
 b15zdnd11an1n64x5 FILLER_254_1174 ();
 b15zdnd11an1n64x5 FILLER_254_1238 ();
 b15zdnd11an1n64x5 FILLER_254_1302 ();
 b15zdnd11an1n64x5 FILLER_254_1366 ();
 b15zdnd11an1n64x5 FILLER_254_1430 ();
 b15zdnd11an1n64x5 FILLER_254_1494 ();
 b15zdnd11an1n64x5 FILLER_254_1558 ();
 b15zdnd11an1n64x5 FILLER_254_1622 ();
 b15zdnd11an1n64x5 FILLER_254_1686 ();
 b15zdnd11an1n64x5 FILLER_254_1750 ();
 b15zdnd11an1n64x5 FILLER_254_1814 ();
 b15zdnd11an1n64x5 FILLER_254_1878 ();
 b15zdnd11an1n64x5 FILLER_254_1942 ();
 b15zdnd11an1n64x5 FILLER_254_2006 ();
 b15zdnd11an1n64x5 FILLER_254_2070 ();
 b15zdnd11an1n16x5 FILLER_254_2134 ();
 b15zdnd11an1n04x5 FILLER_254_2150 ();
 b15zdnd11an1n64x5 FILLER_254_2162 ();
 b15zdnd11an1n32x5 FILLER_254_2226 ();
 b15zdnd11an1n16x5 FILLER_254_2258 ();
 b15zdnd00an1n02x5 FILLER_254_2274 ();
 b15zdnd11an1n64x5 FILLER_255_0 ();
 b15zdnd11an1n64x5 FILLER_255_64 ();
 b15zdnd11an1n64x5 FILLER_255_128 ();
 b15zdnd11an1n64x5 FILLER_255_192 ();
 b15zdnd11an1n64x5 FILLER_255_256 ();
 b15zdnd11an1n64x5 FILLER_255_320 ();
 b15zdnd11an1n64x5 FILLER_255_384 ();
 b15zdnd11an1n64x5 FILLER_255_448 ();
 b15zdnd11an1n64x5 FILLER_255_512 ();
 b15zdnd11an1n64x5 FILLER_255_576 ();
 b15zdnd11an1n64x5 FILLER_255_640 ();
 b15zdnd11an1n64x5 FILLER_255_704 ();
 b15zdnd11an1n64x5 FILLER_255_768 ();
 b15zdnd11an1n64x5 FILLER_255_832 ();
 b15zdnd11an1n64x5 FILLER_255_896 ();
 b15zdnd11an1n64x5 FILLER_255_960 ();
 b15zdnd11an1n64x5 FILLER_255_1024 ();
 b15zdnd11an1n64x5 FILLER_255_1088 ();
 b15zdnd11an1n64x5 FILLER_255_1152 ();
 b15zdnd11an1n64x5 FILLER_255_1216 ();
 b15zdnd11an1n64x5 FILLER_255_1280 ();
 b15zdnd11an1n64x5 FILLER_255_1344 ();
 b15zdnd11an1n64x5 FILLER_255_1408 ();
 b15zdnd11an1n64x5 FILLER_255_1472 ();
 b15zdnd11an1n64x5 FILLER_255_1536 ();
 b15zdnd11an1n64x5 FILLER_255_1600 ();
 b15zdnd11an1n64x5 FILLER_255_1664 ();
 b15zdnd11an1n64x5 FILLER_255_1728 ();
 b15zdnd11an1n64x5 FILLER_255_1792 ();
 b15zdnd11an1n64x5 FILLER_255_1856 ();
 b15zdnd11an1n64x5 FILLER_255_1920 ();
 b15zdnd11an1n64x5 FILLER_255_1984 ();
 b15zdnd11an1n64x5 FILLER_255_2048 ();
 b15zdnd11an1n64x5 FILLER_255_2112 ();
 b15zdnd11an1n64x5 FILLER_255_2176 ();
 b15zdnd11an1n32x5 FILLER_255_2240 ();
 b15zdnd11an1n08x5 FILLER_255_2272 ();
 b15zdnd11an1n04x5 FILLER_255_2280 ();
 b15zdnd11an1n64x5 FILLER_256_8 ();
 b15zdnd11an1n64x5 FILLER_256_72 ();
 b15zdnd11an1n64x5 FILLER_256_136 ();
 b15zdnd11an1n64x5 FILLER_256_200 ();
 b15zdnd11an1n64x5 FILLER_256_264 ();
 b15zdnd11an1n64x5 FILLER_256_328 ();
 b15zdnd11an1n64x5 FILLER_256_392 ();
 b15zdnd11an1n64x5 FILLER_256_456 ();
 b15zdnd11an1n64x5 FILLER_256_520 ();
 b15zdnd11an1n64x5 FILLER_256_584 ();
 b15zdnd11an1n64x5 FILLER_256_648 ();
 b15zdnd11an1n04x5 FILLER_256_712 ();
 b15zdnd00an1n02x5 FILLER_256_716 ();
 b15zdnd11an1n64x5 FILLER_256_726 ();
 b15zdnd11an1n64x5 FILLER_256_790 ();
 b15zdnd11an1n64x5 FILLER_256_854 ();
 b15zdnd11an1n64x5 FILLER_256_918 ();
 b15zdnd11an1n64x5 FILLER_256_982 ();
 b15zdnd11an1n64x5 FILLER_256_1046 ();
 b15zdnd11an1n64x5 FILLER_256_1110 ();
 b15zdnd11an1n64x5 FILLER_256_1174 ();
 b15zdnd11an1n04x5 FILLER_256_1238 ();
 b15zdnd00an1n02x5 FILLER_256_1242 ();
 b15zdnd11an1n04x5 FILLER_256_1255 ();
 b15zdnd11an1n64x5 FILLER_256_1275 ();
 b15zdnd11an1n64x5 FILLER_256_1339 ();
 b15zdnd11an1n64x5 FILLER_256_1403 ();
 b15zdnd11an1n64x5 FILLER_256_1467 ();
 b15zdnd11an1n64x5 FILLER_256_1531 ();
 b15zdnd11an1n64x5 FILLER_256_1595 ();
 b15zdnd11an1n64x5 FILLER_256_1659 ();
 b15zdnd11an1n64x5 FILLER_256_1723 ();
 b15zdnd11an1n64x5 FILLER_256_1787 ();
 b15zdnd11an1n64x5 FILLER_256_1851 ();
 b15zdnd11an1n64x5 FILLER_256_1915 ();
 b15zdnd11an1n64x5 FILLER_256_1979 ();
 b15zdnd11an1n64x5 FILLER_256_2043 ();
 b15zdnd11an1n32x5 FILLER_256_2107 ();
 b15zdnd11an1n08x5 FILLER_256_2139 ();
 b15zdnd11an1n04x5 FILLER_256_2147 ();
 b15zdnd00an1n02x5 FILLER_256_2151 ();
 b15zdnd00an1n01x5 FILLER_256_2153 ();
 b15zdnd11an1n64x5 FILLER_256_2162 ();
 b15zdnd11an1n32x5 FILLER_256_2226 ();
 b15zdnd11an1n16x5 FILLER_256_2258 ();
 b15zdnd00an1n02x5 FILLER_256_2274 ();
 b15zdnd11an1n64x5 FILLER_257_0 ();
 b15zdnd11an1n64x5 FILLER_257_64 ();
 b15zdnd11an1n64x5 FILLER_257_128 ();
 b15zdnd11an1n64x5 FILLER_257_192 ();
 b15zdnd11an1n64x5 FILLER_257_256 ();
 b15zdnd11an1n64x5 FILLER_257_320 ();
 b15zdnd11an1n64x5 FILLER_257_384 ();
 b15zdnd11an1n64x5 FILLER_257_448 ();
 b15zdnd11an1n64x5 FILLER_257_512 ();
 b15zdnd11an1n64x5 FILLER_257_576 ();
 b15zdnd11an1n64x5 FILLER_257_640 ();
 b15zdnd11an1n64x5 FILLER_257_704 ();
 b15zdnd11an1n64x5 FILLER_257_768 ();
 b15zdnd11an1n64x5 FILLER_257_832 ();
 b15zdnd11an1n64x5 FILLER_257_896 ();
 b15zdnd11an1n64x5 FILLER_257_960 ();
 b15zdnd11an1n64x5 FILLER_257_1024 ();
 b15zdnd11an1n64x5 FILLER_257_1088 ();
 b15zdnd11an1n64x5 FILLER_257_1152 ();
 b15zdnd11an1n32x5 FILLER_257_1216 ();
 b15zdnd00an1n02x5 FILLER_257_1248 ();
 b15zdnd00an1n01x5 FILLER_257_1250 ();
 b15zdnd11an1n64x5 FILLER_257_1293 ();
 b15zdnd11an1n64x5 FILLER_257_1357 ();
 b15zdnd11an1n64x5 FILLER_257_1421 ();
 b15zdnd11an1n64x5 FILLER_257_1485 ();
 b15zdnd11an1n64x5 FILLER_257_1549 ();
 b15zdnd11an1n64x5 FILLER_257_1613 ();
 b15zdnd11an1n64x5 FILLER_257_1677 ();
 b15zdnd11an1n64x5 FILLER_257_1741 ();
 b15zdnd11an1n64x5 FILLER_257_1805 ();
 b15zdnd11an1n64x5 FILLER_257_1869 ();
 b15zdnd11an1n64x5 FILLER_257_1933 ();
 b15zdnd11an1n64x5 FILLER_257_1997 ();
 b15zdnd11an1n64x5 FILLER_257_2061 ();
 b15zdnd11an1n64x5 FILLER_257_2125 ();
 b15zdnd11an1n64x5 FILLER_257_2189 ();
 b15zdnd11an1n16x5 FILLER_257_2253 ();
 b15zdnd11an1n08x5 FILLER_257_2269 ();
 b15zdnd11an1n04x5 FILLER_257_2277 ();
 b15zdnd00an1n02x5 FILLER_257_2281 ();
 b15zdnd00an1n01x5 FILLER_257_2283 ();
 b15zdnd11an1n64x5 FILLER_258_8 ();
 b15zdnd11an1n64x5 FILLER_258_72 ();
 b15zdnd11an1n64x5 FILLER_258_136 ();
 b15zdnd11an1n64x5 FILLER_258_200 ();
 b15zdnd11an1n64x5 FILLER_258_264 ();
 b15zdnd11an1n64x5 FILLER_258_328 ();
 b15zdnd11an1n64x5 FILLER_258_392 ();
 b15zdnd11an1n64x5 FILLER_258_456 ();
 b15zdnd11an1n64x5 FILLER_258_520 ();
 b15zdnd11an1n64x5 FILLER_258_584 ();
 b15zdnd11an1n64x5 FILLER_258_648 ();
 b15zdnd11an1n04x5 FILLER_258_712 ();
 b15zdnd00an1n02x5 FILLER_258_716 ();
 b15zdnd11an1n64x5 FILLER_258_726 ();
 b15zdnd11an1n64x5 FILLER_258_790 ();
 b15zdnd11an1n64x5 FILLER_258_854 ();
 b15zdnd11an1n64x5 FILLER_258_918 ();
 b15zdnd11an1n64x5 FILLER_258_982 ();
 b15zdnd11an1n64x5 FILLER_258_1046 ();
 b15zdnd11an1n64x5 FILLER_258_1110 ();
 b15zdnd11an1n64x5 FILLER_258_1174 ();
 b15zdnd11an1n04x5 FILLER_258_1238 ();
 b15zdnd00an1n02x5 FILLER_258_1242 ();
 b15zdnd00an1n01x5 FILLER_258_1244 ();
 b15zdnd11an1n04x5 FILLER_258_1255 ();
 b15zdnd11an1n64x5 FILLER_258_1266 ();
 b15zdnd11an1n64x5 FILLER_258_1330 ();
 b15zdnd11an1n64x5 FILLER_258_1394 ();
 b15zdnd11an1n64x5 FILLER_258_1458 ();
 b15zdnd11an1n64x5 FILLER_258_1522 ();
 b15zdnd11an1n64x5 FILLER_258_1586 ();
 b15zdnd11an1n64x5 FILLER_258_1650 ();
 b15zdnd11an1n64x5 FILLER_258_1714 ();
 b15zdnd11an1n64x5 FILLER_258_1778 ();
 b15zdnd11an1n64x5 FILLER_258_1842 ();
 b15zdnd11an1n64x5 FILLER_258_1906 ();
 b15zdnd11an1n64x5 FILLER_258_1970 ();
 b15zdnd11an1n64x5 FILLER_258_2034 ();
 b15zdnd11an1n32x5 FILLER_258_2098 ();
 b15zdnd11an1n16x5 FILLER_258_2130 ();
 b15zdnd11an1n08x5 FILLER_258_2146 ();
 b15zdnd11an1n64x5 FILLER_258_2162 ();
 b15zdnd11an1n32x5 FILLER_258_2226 ();
 b15zdnd11an1n16x5 FILLER_258_2258 ();
 b15zdnd00an1n02x5 FILLER_258_2274 ();
 b15zdnd11an1n64x5 FILLER_259_0 ();
 b15zdnd11an1n64x5 FILLER_259_64 ();
 b15zdnd11an1n64x5 FILLER_259_128 ();
 b15zdnd11an1n64x5 FILLER_259_192 ();
 b15zdnd11an1n64x5 FILLER_259_256 ();
 b15zdnd11an1n64x5 FILLER_259_320 ();
 b15zdnd11an1n64x5 FILLER_259_384 ();
 b15zdnd11an1n64x5 FILLER_259_448 ();
 b15zdnd11an1n64x5 FILLER_259_512 ();
 b15zdnd11an1n64x5 FILLER_259_576 ();
 b15zdnd11an1n64x5 FILLER_259_640 ();
 b15zdnd11an1n64x5 FILLER_259_704 ();
 b15zdnd11an1n64x5 FILLER_259_768 ();
 b15zdnd11an1n64x5 FILLER_259_832 ();
 b15zdnd11an1n64x5 FILLER_259_896 ();
 b15zdnd11an1n64x5 FILLER_259_960 ();
 b15zdnd11an1n64x5 FILLER_259_1024 ();
 b15zdnd11an1n64x5 FILLER_259_1088 ();
 b15zdnd11an1n64x5 FILLER_259_1152 ();
 b15zdnd11an1n64x5 FILLER_259_1216 ();
 b15zdnd11an1n64x5 FILLER_259_1280 ();
 b15zdnd11an1n64x5 FILLER_259_1344 ();
 b15zdnd11an1n64x5 FILLER_259_1408 ();
 b15zdnd11an1n64x5 FILLER_259_1472 ();
 b15zdnd11an1n64x5 FILLER_259_1536 ();
 b15zdnd11an1n64x5 FILLER_259_1600 ();
 b15zdnd11an1n64x5 FILLER_259_1664 ();
 b15zdnd11an1n64x5 FILLER_259_1728 ();
 b15zdnd11an1n64x5 FILLER_259_1792 ();
 b15zdnd11an1n64x5 FILLER_259_1856 ();
 b15zdnd11an1n64x5 FILLER_259_1920 ();
 b15zdnd11an1n64x5 FILLER_259_1984 ();
 b15zdnd11an1n64x5 FILLER_259_2048 ();
 b15zdnd11an1n64x5 FILLER_259_2112 ();
 b15zdnd11an1n64x5 FILLER_259_2176 ();
 b15zdnd11an1n32x5 FILLER_259_2240 ();
 b15zdnd11an1n08x5 FILLER_259_2272 ();
 b15zdnd11an1n04x5 FILLER_259_2280 ();
 b15zdnd11an1n64x5 FILLER_260_8 ();
 b15zdnd11an1n64x5 FILLER_260_72 ();
 b15zdnd11an1n64x5 FILLER_260_136 ();
 b15zdnd11an1n64x5 FILLER_260_200 ();
 b15zdnd11an1n64x5 FILLER_260_264 ();
 b15zdnd11an1n64x5 FILLER_260_328 ();
 b15zdnd11an1n64x5 FILLER_260_392 ();
 b15zdnd11an1n64x5 FILLER_260_456 ();
 b15zdnd11an1n64x5 FILLER_260_520 ();
 b15zdnd11an1n64x5 FILLER_260_584 ();
 b15zdnd11an1n64x5 FILLER_260_648 ();
 b15zdnd11an1n04x5 FILLER_260_712 ();
 b15zdnd00an1n02x5 FILLER_260_716 ();
 b15zdnd11an1n64x5 FILLER_260_726 ();
 b15zdnd11an1n64x5 FILLER_260_790 ();
 b15zdnd11an1n64x5 FILLER_260_854 ();
 b15zdnd11an1n64x5 FILLER_260_918 ();
 b15zdnd11an1n64x5 FILLER_260_982 ();
 b15zdnd11an1n64x5 FILLER_260_1046 ();
 b15zdnd11an1n64x5 FILLER_260_1110 ();
 b15zdnd11an1n64x5 FILLER_260_1174 ();
 b15zdnd11an1n64x5 FILLER_260_1238 ();
 b15zdnd11an1n64x5 FILLER_260_1302 ();
 b15zdnd11an1n64x5 FILLER_260_1366 ();
 b15zdnd11an1n64x5 FILLER_260_1430 ();
 b15zdnd11an1n64x5 FILLER_260_1494 ();
 b15zdnd11an1n64x5 FILLER_260_1558 ();
 b15zdnd11an1n64x5 FILLER_260_1622 ();
 b15zdnd11an1n64x5 FILLER_260_1686 ();
 b15zdnd11an1n64x5 FILLER_260_1750 ();
 b15zdnd11an1n64x5 FILLER_260_1814 ();
 b15zdnd11an1n64x5 FILLER_260_1878 ();
 b15zdnd11an1n64x5 FILLER_260_1942 ();
 b15zdnd11an1n64x5 FILLER_260_2006 ();
 b15zdnd11an1n64x5 FILLER_260_2070 ();
 b15zdnd11an1n16x5 FILLER_260_2134 ();
 b15zdnd11an1n04x5 FILLER_260_2150 ();
 b15zdnd11an1n64x5 FILLER_260_2162 ();
 b15zdnd11an1n32x5 FILLER_260_2226 ();
 b15zdnd11an1n16x5 FILLER_260_2258 ();
 b15zdnd00an1n02x5 FILLER_260_2274 ();
 b15zdnd11an1n64x5 FILLER_261_0 ();
 b15zdnd11an1n64x5 FILLER_261_64 ();
 b15zdnd11an1n64x5 FILLER_261_128 ();
 b15zdnd11an1n64x5 FILLER_261_192 ();
 b15zdnd11an1n64x5 FILLER_261_256 ();
 b15zdnd11an1n64x5 FILLER_261_320 ();
 b15zdnd11an1n64x5 FILLER_261_384 ();
 b15zdnd11an1n64x5 FILLER_261_448 ();
 b15zdnd11an1n64x5 FILLER_261_512 ();
 b15zdnd11an1n64x5 FILLER_261_576 ();
 b15zdnd11an1n64x5 FILLER_261_640 ();
 b15zdnd11an1n64x5 FILLER_261_704 ();
 b15zdnd11an1n64x5 FILLER_261_768 ();
 b15zdnd11an1n64x5 FILLER_261_832 ();
 b15zdnd11an1n64x5 FILLER_261_896 ();
 b15zdnd11an1n64x5 FILLER_261_960 ();
 b15zdnd11an1n64x5 FILLER_261_1024 ();
 b15zdnd11an1n64x5 FILLER_261_1088 ();
 b15zdnd11an1n64x5 FILLER_261_1152 ();
 b15zdnd11an1n64x5 FILLER_261_1216 ();
 b15zdnd11an1n64x5 FILLER_261_1280 ();
 b15zdnd11an1n64x5 FILLER_261_1344 ();
 b15zdnd11an1n64x5 FILLER_261_1408 ();
 b15zdnd11an1n64x5 FILLER_261_1472 ();
 b15zdnd11an1n64x5 FILLER_261_1536 ();
 b15zdnd11an1n64x5 FILLER_261_1600 ();
 b15zdnd11an1n64x5 FILLER_261_1664 ();
 b15zdnd11an1n64x5 FILLER_261_1728 ();
 b15zdnd11an1n64x5 FILLER_261_1792 ();
 b15zdnd11an1n64x5 FILLER_261_1856 ();
 b15zdnd11an1n64x5 FILLER_261_1920 ();
 b15zdnd11an1n64x5 FILLER_261_1984 ();
 b15zdnd11an1n64x5 FILLER_261_2048 ();
 b15zdnd11an1n16x5 FILLER_261_2112 ();
 b15zdnd11an1n08x5 FILLER_261_2128 ();
 b15zdnd11an1n04x5 FILLER_261_2136 ();
 b15zdnd00an1n02x5 FILLER_261_2140 ();
 b15zdnd00an1n01x5 FILLER_261_2142 ();
 b15zdnd11an1n64x5 FILLER_261_2159 ();
 b15zdnd11an1n32x5 FILLER_261_2223 ();
 b15zdnd11an1n16x5 FILLER_261_2255 ();
 b15zdnd11an1n08x5 FILLER_261_2271 ();
 b15zdnd11an1n04x5 FILLER_261_2279 ();
 b15zdnd00an1n01x5 FILLER_261_2283 ();
 b15zdnd11an1n64x5 FILLER_262_8 ();
 b15zdnd11an1n64x5 FILLER_262_72 ();
 b15zdnd11an1n64x5 FILLER_262_136 ();
 b15zdnd11an1n64x5 FILLER_262_200 ();
 b15zdnd11an1n64x5 FILLER_262_264 ();
 b15zdnd11an1n64x5 FILLER_262_328 ();
 b15zdnd11an1n64x5 FILLER_262_392 ();
 b15zdnd11an1n64x5 FILLER_262_456 ();
 b15zdnd11an1n64x5 FILLER_262_520 ();
 b15zdnd11an1n64x5 FILLER_262_584 ();
 b15zdnd11an1n64x5 FILLER_262_648 ();
 b15zdnd11an1n04x5 FILLER_262_712 ();
 b15zdnd00an1n02x5 FILLER_262_716 ();
 b15zdnd11an1n64x5 FILLER_262_726 ();
 b15zdnd11an1n64x5 FILLER_262_790 ();
 b15zdnd11an1n64x5 FILLER_262_854 ();
 b15zdnd11an1n64x5 FILLER_262_918 ();
 b15zdnd11an1n64x5 FILLER_262_982 ();
 b15zdnd11an1n64x5 FILLER_262_1046 ();
 b15zdnd11an1n64x5 FILLER_262_1110 ();
 b15zdnd11an1n64x5 FILLER_262_1174 ();
 b15zdnd11an1n64x5 FILLER_262_1238 ();
 b15zdnd11an1n64x5 FILLER_262_1302 ();
 b15zdnd11an1n64x5 FILLER_262_1366 ();
 b15zdnd11an1n64x5 FILLER_262_1430 ();
 b15zdnd11an1n64x5 FILLER_262_1494 ();
 b15zdnd11an1n64x5 FILLER_262_1558 ();
 b15zdnd11an1n64x5 FILLER_262_1622 ();
 b15zdnd11an1n64x5 FILLER_262_1686 ();
 b15zdnd11an1n64x5 FILLER_262_1750 ();
 b15zdnd11an1n64x5 FILLER_262_1814 ();
 b15zdnd11an1n64x5 FILLER_262_1878 ();
 b15zdnd11an1n64x5 FILLER_262_1942 ();
 b15zdnd11an1n64x5 FILLER_262_2006 ();
 b15zdnd11an1n64x5 FILLER_262_2070 ();
 b15zdnd11an1n16x5 FILLER_262_2134 ();
 b15zdnd11an1n04x5 FILLER_262_2150 ();
 b15zdnd11an1n64x5 FILLER_262_2162 ();
 b15zdnd11an1n32x5 FILLER_262_2226 ();
 b15zdnd11an1n16x5 FILLER_262_2258 ();
 b15zdnd00an1n02x5 FILLER_262_2274 ();
 b15zdnd11an1n64x5 FILLER_263_0 ();
 b15zdnd11an1n64x5 FILLER_263_64 ();
 b15zdnd11an1n64x5 FILLER_263_128 ();
 b15zdnd11an1n64x5 FILLER_263_192 ();
 b15zdnd11an1n64x5 FILLER_263_256 ();
 b15zdnd11an1n64x5 FILLER_263_320 ();
 b15zdnd11an1n64x5 FILLER_263_384 ();
 b15zdnd11an1n64x5 FILLER_263_448 ();
 b15zdnd11an1n64x5 FILLER_263_512 ();
 b15zdnd11an1n64x5 FILLER_263_576 ();
 b15zdnd11an1n64x5 FILLER_263_640 ();
 b15zdnd11an1n64x5 FILLER_263_704 ();
 b15zdnd11an1n64x5 FILLER_263_768 ();
 b15zdnd11an1n64x5 FILLER_263_832 ();
 b15zdnd11an1n64x5 FILLER_263_896 ();
 b15zdnd11an1n64x5 FILLER_263_960 ();
 b15zdnd11an1n64x5 FILLER_263_1024 ();
 b15zdnd11an1n64x5 FILLER_263_1088 ();
 b15zdnd11an1n64x5 FILLER_263_1152 ();
 b15zdnd11an1n64x5 FILLER_263_1216 ();
 b15zdnd11an1n64x5 FILLER_263_1280 ();
 b15zdnd11an1n64x5 FILLER_263_1344 ();
 b15zdnd11an1n64x5 FILLER_263_1408 ();
 b15zdnd11an1n64x5 FILLER_263_1472 ();
 b15zdnd11an1n64x5 FILLER_263_1536 ();
 b15zdnd11an1n64x5 FILLER_263_1600 ();
 b15zdnd11an1n64x5 FILLER_263_1664 ();
 b15zdnd11an1n64x5 FILLER_263_1728 ();
 b15zdnd11an1n64x5 FILLER_263_1792 ();
 b15zdnd11an1n64x5 FILLER_263_1856 ();
 b15zdnd11an1n64x5 FILLER_263_1920 ();
 b15zdnd11an1n64x5 FILLER_263_1984 ();
 b15zdnd11an1n64x5 FILLER_263_2048 ();
 b15zdnd11an1n64x5 FILLER_263_2112 ();
 b15zdnd11an1n64x5 FILLER_263_2176 ();
 b15zdnd11an1n32x5 FILLER_263_2240 ();
 b15zdnd11an1n08x5 FILLER_263_2272 ();
 b15zdnd11an1n04x5 FILLER_263_2280 ();
 b15zdnd11an1n64x5 FILLER_264_8 ();
 b15zdnd11an1n64x5 FILLER_264_72 ();
 b15zdnd11an1n64x5 FILLER_264_136 ();
 b15zdnd11an1n64x5 FILLER_264_200 ();
 b15zdnd11an1n64x5 FILLER_264_264 ();
 b15zdnd11an1n64x5 FILLER_264_328 ();
 b15zdnd11an1n64x5 FILLER_264_392 ();
 b15zdnd11an1n64x5 FILLER_264_456 ();
 b15zdnd11an1n64x5 FILLER_264_520 ();
 b15zdnd11an1n64x5 FILLER_264_584 ();
 b15zdnd11an1n64x5 FILLER_264_648 ();
 b15zdnd11an1n04x5 FILLER_264_712 ();
 b15zdnd00an1n02x5 FILLER_264_716 ();
 b15zdnd11an1n64x5 FILLER_264_726 ();
 b15zdnd11an1n64x5 FILLER_264_790 ();
 b15zdnd11an1n64x5 FILLER_264_854 ();
 b15zdnd11an1n64x5 FILLER_264_918 ();
 b15zdnd11an1n64x5 FILLER_264_982 ();
 b15zdnd11an1n64x5 FILLER_264_1046 ();
 b15zdnd11an1n64x5 FILLER_264_1110 ();
 b15zdnd11an1n64x5 FILLER_264_1174 ();
 b15zdnd11an1n64x5 FILLER_264_1238 ();
 b15zdnd11an1n64x5 FILLER_264_1302 ();
 b15zdnd11an1n64x5 FILLER_264_1366 ();
 b15zdnd11an1n64x5 FILLER_264_1430 ();
 b15zdnd11an1n64x5 FILLER_264_1494 ();
 b15zdnd11an1n64x5 FILLER_264_1558 ();
 b15zdnd11an1n64x5 FILLER_264_1622 ();
 b15zdnd11an1n64x5 FILLER_264_1686 ();
 b15zdnd11an1n64x5 FILLER_264_1750 ();
 b15zdnd11an1n64x5 FILLER_264_1814 ();
 b15zdnd11an1n64x5 FILLER_264_1878 ();
 b15zdnd11an1n64x5 FILLER_264_1942 ();
 b15zdnd11an1n64x5 FILLER_264_2006 ();
 b15zdnd11an1n64x5 FILLER_264_2070 ();
 b15zdnd11an1n16x5 FILLER_264_2134 ();
 b15zdnd11an1n04x5 FILLER_264_2150 ();
 b15zdnd11an1n64x5 FILLER_264_2162 ();
 b15zdnd11an1n32x5 FILLER_264_2226 ();
 b15zdnd11an1n16x5 FILLER_264_2258 ();
 b15zdnd00an1n02x5 FILLER_264_2274 ();
 b15zdnd11an1n64x5 FILLER_265_0 ();
 b15zdnd11an1n64x5 FILLER_265_64 ();
 b15zdnd11an1n64x5 FILLER_265_128 ();
 b15zdnd11an1n64x5 FILLER_265_192 ();
 b15zdnd11an1n64x5 FILLER_265_256 ();
 b15zdnd11an1n64x5 FILLER_265_320 ();
 b15zdnd11an1n64x5 FILLER_265_384 ();
 b15zdnd11an1n64x5 FILLER_265_448 ();
 b15zdnd11an1n64x5 FILLER_265_512 ();
 b15zdnd11an1n64x5 FILLER_265_576 ();
 b15zdnd11an1n64x5 FILLER_265_640 ();
 b15zdnd11an1n64x5 FILLER_265_704 ();
 b15zdnd11an1n64x5 FILLER_265_768 ();
 b15zdnd11an1n64x5 FILLER_265_832 ();
 b15zdnd11an1n64x5 FILLER_265_896 ();
 b15zdnd11an1n64x5 FILLER_265_960 ();
 b15zdnd11an1n64x5 FILLER_265_1024 ();
 b15zdnd11an1n64x5 FILLER_265_1088 ();
 b15zdnd11an1n64x5 FILLER_265_1152 ();
 b15zdnd11an1n64x5 FILLER_265_1216 ();
 b15zdnd11an1n64x5 FILLER_265_1280 ();
 b15zdnd11an1n64x5 FILLER_265_1344 ();
 b15zdnd11an1n64x5 FILLER_265_1408 ();
 b15zdnd11an1n64x5 FILLER_265_1472 ();
 b15zdnd11an1n64x5 FILLER_265_1536 ();
 b15zdnd11an1n64x5 FILLER_265_1600 ();
 b15zdnd11an1n64x5 FILLER_265_1664 ();
 b15zdnd11an1n64x5 FILLER_265_1728 ();
 b15zdnd11an1n64x5 FILLER_265_1792 ();
 b15zdnd11an1n64x5 FILLER_265_1856 ();
 b15zdnd11an1n64x5 FILLER_265_1920 ();
 b15zdnd11an1n64x5 FILLER_265_1984 ();
 b15zdnd11an1n64x5 FILLER_265_2048 ();
 b15zdnd11an1n64x5 FILLER_265_2112 ();
 b15zdnd11an1n64x5 FILLER_265_2176 ();
 b15zdnd11an1n32x5 FILLER_265_2240 ();
 b15zdnd11an1n08x5 FILLER_265_2272 ();
 b15zdnd11an1n04x5 FILLER_265_2280 ();
 b15zdnd11an1n64x5 FILLER_266_8 ();
 b15zdnd11an1n64x5 FILLER_266_72 ();
 b15zdnd11an1n64x5 FILLER_266_136 ();
 b15zdnd11an1n64x5 FILLER_266_200 ();
 b15zdnd11an1n64x5 FILLER_266_264 ();
 b15zdnd11an1n64x5 FILLER_266_328 ();
 b15zdnd11an1n64x5 FILLER_266_392 ();
 b15zdnd11an1n64x5 FILLER_266_456 ();
 b15zdnd11an1n64x5 FILLER_266_520 ();
 b15zdnd11an1n64x5 FILLER_266_584 ();
 b15zdnd11an1n64x5 FILLER_266_648 ();
 b15zdnd11an1n04x5 FILLER_266_712 ();
 b15zdnd00an1n02x5 FILLER_266_716 ();
 b15zdnd11an1n64x5 FILLER_266_726 ();
 b15zdnd11an1n64x5 FILLER_266_790 ();
 b15zdnd11an1n64x5 FILLER_266_854 ();
 b15zdnd11an1n64x5 FILLER_266_918 ();
 b15zdnd11an1n64x5 FILLER_266_982 ();
 b15zdnd11an1n64x5 FILLER_266_1046 ();
 b15zdnd11an1n64x5 FILLER_266_1110 ();
 b15zdnd11an1n64x5 FILLER_266_1174 ();
 b15zdnd11an1n64x5 FILLER_266_1238 ();
 b15zdnd11an1n64x5 FILLER_266_1302 ();
 b15zdnd11an1n64x5 FILLER_266_1366 ();
 b15zdnd11an1n64x5 FILLER_266_1430 ();
 b15zdnd11an1n64x5 FILLER_266_1494 ();
 b15zdnd11an1n64x5 FILLER_266_1558 ();
 b15zdnd11an1n16x5 FILLER_266_1622 ();
 b15zdnd00an1n02x5 FILLER_266_1638 ();
 b15zdnd11an1n04x5 FILLER_266_1651 ();
 b15zdnd11an1n64x5 FILLER_266_1661 ();
 b15zdnd11an1n64x5 FILLER_266_1725 ();
 b15zdnd11an1n64x5 FILLER_266_1789 ();
 b15zdnd11an1n64x5 FILLER_266_1853 ();
 b15zdnd11an1n64x5 FILLER_266_1917 ();
 b15zdnd11an1n64x5 FILLER_266_1981 ();
 b15zdnd11an1n64x5 FILLER_266_2045 ();
 b15zdnd11an1n32x5 FILLER_266_2109 ();
 b15zdnd11an1n08x5 FILLER_266_2141 ();
 b15zdnd11an1n04x5 FILLER_266_2149 ();
 b15zdnd00an1n01x5 FILLER_266_2153 ();
 b15zdnd11an1n64x5 FILLER_266_2162 ();
 b15zdnd11an1n32x5 FILLER_266_2226 ();
 b15zdnd11an1n16x5 FILLER_266_2258 ();
 b15zdnd00an1n02x5 FILLER_266_2274 ();
 b15zdnd11an1n64x5 FILLER_267_0 ();
 b15zdnd11an1n64x5 FILLER_267_64 ();
 b15zdnd11an1n64x5 FILLER_267_128 ();
 b15zdnd11an1n64x5 FILLER_267_192 ();
 b15zdnd11an1n64x5 FILLER_267_256 ();
 b15zdnd11an1n64x5 FILLER_267_320 ();
 b15zdnd11an1n64x5 FILLER_267_384 ();
 b15zdnd11an1n64x5 FILLER_267_448 ();
 b15zdnd11an1n64x5 FILLER_267_512 ();
 b15zdnd11an1n64x5 FILLER_267_576 ();
 b15zdnd11an1n64x5 FILLER_267_640 ();
 b15zdnd11an1n64x5 FILLER_267_704 ();
 b15zdnd11an1n64x5 FILLER_267_768 ();
 b15zdnd11an1n64x5 FILLER_267_832 ();
 b15zdnd11an1n64x5 FILLER_267_896 ();
 b15zdnd11an1n64x5 FILLER_267_960 ();
 b15zdnd11an1n64x5 FILLER_267_1024 ();
 b15zdnd11an1n64x5 FILLER_267_1088 ();
 b15zdnd11an1n64x5 FILLER_267_1152 ();
 b15zdnd11an1n64x5 FILLER_267_1216 ();
 b15zdnd11an1n64x5 FILLER_267_1280 ();
 b15zdnd11an1n64x5 FILLER_267_1344 ();
 b15zdnd11an1n64x5 FILLER_267_1408 ();
 b15zdnd11an1n64x5 FILLER_267_1472 ();
 b15zdnd11an1n64x5 FILLER_267_1536 ();
 b15zdnd11an1n64x5 FILLER_267_1600 ();
 b15zdnd11an1n64x5 FILLER_267_1664 ();
 b15zdnd11an1n64x5 FILLER_267_1728 ();
 b15zdnd11an1n64x5 FILLER_267_1792 ();
 b15zdnd11an1n64x5 FILLER_267_1856 ();
 b15zdnd11an1n64x5 FILLER_267_1920 ();
 b15zdnd11an1n64x5 FILLER_267_1984 ();
 b15zdnd11an1n64x5 FILLER_267_2048 ();
 b15zdnd11an1n64x5 FILLER_267_2112 ();
 b15zdnd11an1n64x5 FILLER_267_2176 ();
 b15zdnd11an1n32x5 FILLER_267_2240 ();
 b15zdnd11an1n08x5 FILLER_267_2272 ();
 b15zdnd11an1n04x5 FILLER_267_2280 ();
 b15zdnd11an1n64x5 FILLER_268_8 ();
 b15zdnd11an1n64x5 FILLER_268_72 ();
 b15zdnd11an1n64x5 FILLER_268_136 ();
 b15zdnd11an1n64x5 FILLER_268_200 ();
 b15zdnd11an1n64x5 FILLER_268_264 ();
 b15zdnd11an1n64x5 FILLER_268_328 ();
 b15zdnd11an1n64x5 FILLER_268_392 ();
 b15zdnd11an1n64x5 FILLER_268_456 ();
 b15zdnd11an1n64x5 FILLER_268_520 ();
 b15zdnd11an1n64x5 FILLER_268_584 ();
 b15zdnd11an1n64x5 FILLER_268_648 ();
 b15zdnd11an1n04x5 FILLER_268_712 ();
 b15zdnd00an1n02x5 FILLER_268_716 ();
 b15zdnd11an1n64x5 FILLER_268_726 ();
 b15zdnd11an1n64x5 FILLER_268_790 ();
 b15zdnd11an1n64x5 FILLER_268_854 ();
 b15zdnd11an1n64x5 FILLER_268_918 ();
 b15zdnd11an1n64x5 FILLER_268_982 ();
 b15zdnd11an1n64x5 FILLER_268_1046 ();
 b15zdnd11an1n64x5 FILLER_268_1110 ();
 b15zdnd11an1n64x5 FILLER_268_1174 ();
 b15zdnd11an1n64x5 FILLER_268_1238 ();
 b15zdnd11an1n64x5 FILLER_268_1302 ();
 b15zdnd11an1n64x5 FILLER_268_1366 ();
 b15zdnd11an1n64x5 FILLER_268_1430 ();
 b15zdnd11an1n64x5 FILLER_268_1494 ();
 b15zdnd11an1n64x5 FILLER_268_1558 ();
 b15zdnd11an1n64x5 FILLER_268_1622 ();
 b15zdnd11an1n64x5 FILLER_268_1686 ();
 b15zdnd11an1n64x5 FILLER_268_1750 ();
 b15zdnd11an1n64x5 FILLER_268_1814 ();
 b15zdnd11an1n64x5 FILLER_268_1878 ();
 b15zdnd11an1n64x5 FILLER_268_1942 ();
 b15zdnd11an1n64x5 FILLER_268_2006 ();
 b15zdnd11an1n64x5 FILLER_268_2070 ();
 b15zdnd11an1n16x5 FILLER_268_2134 ();
 b15zdnd11an1n04x5 FILLER_268_2150 ();
 b15zdnd11an1n64x5 FILLER_268_2162 ();
 b15zdnd11an1n32x5 FILLER_268_2226 ();
 b15zdnd11an1n16x5 FILLER_268_2258 ();
 b15zdnd00an1n02x5 FILLER_268_2274 ();
 b15zdnd11an1n64x5 FILLER_269_0 ();
 b15zdnd11an1n64x5 FILLER_269_64 ();
 b15zdnd11an1n64x5 FILLER_269_128 ();
 b15zdnd11an1n64x5 FILLER_269_192 ();
 b15zdnd11an1n64x5 FILLER_269_256 ();
 b15zdnd11an1n64x5 FILLER_269_320 ();
 b15zdnd11an1n64x5 FILLER_269_384 ();
 b15zdnd11an1n64x5 FILLER_269_448 ();
 b15zdnd11an1n64x5 FILLER_269_512 ();
 b15zdnd11an1n64x5 FILLER_269_576 ();
 b15zdnd11an1n64x5 FILLER_269_640 ();
 b15zdnd11an1n64x5 FILLER_269_704 ();
 b15zdnd11an1n64x5 FILLER_269_768 ();
 b15zdnd11an1n64x5 FILLER_269_832 ();
 b15zdnd11an1n64x5 FILLER_269_896 ();
 b15zdnd11an1n64x5 FILLER_269_960 ();
 b15zdnd11an1n64x5 FILLER_269_1024 ();
 b15zdnd11an1n64x5 FILLER_269_1088 ();
 b15zdnd11an1n64x5 FILLER_269_1152 ();
 b15zdnd11an1n64x5 FILLER_269_1216 ();
 b15zdnd11an1n64x5 FILLER_269_1280 ();
 b15zdnd11an1n64x5 FILLER_269_1344 ();
 b15zdnd11an1n64x5 FILLER_269_1408 ();
 b15zdnd11an1n64x5 FILLER_269_1472 ();
 b15zdnd11an1n64x5 FILLER_269_1536 ();
 b15zdnd11an1n64x5 FILLER_269_1600 ();
 b15zdnd11an1n64x5 FILLER_269_1664 ();
 b15zdnd11an1n64x5 FILLER_269_1728 ();
 b15zdnd11an1n64x5 FILLER_269_1792 ();
 b15zdnd11an1n64x5 FILLER_269_1856 ();
 b15zdnd11an1n64x5 FILLER_269_1920 ();
 b15zdnd11an1n64x5 FILLER_269_1984 ();
 b15zdnd11an1n64x5 FILLER_269_2048 ();
 b15zdnd11an1n64x5 FILLER_269_2112 ();
 b15zdnd11an1n64x5 FILLER_269_2176 ();
 b15zdnd11an1n32x5 FILLER_269_2240 ();
 b15zdnd11an1n08x5 FILLER_269_2272 ();
 b15zdnd11an1n04x5 FILLER_269_2280 ();
 b15zdnd11an1n64x5 FILLER_270_8 ();
 b15zdnd11an1n64x5 FILLER_270_72 ();
 b15zdnd11an1n64x5 FILLER_270_136 ();
 b15zdnd11an1n64x5 FILLER_270_200 ();
 b15zdnd11an1n64x5 FILLER_270_264 ();
 b15zdnd11an1n64x5 FILLER_270_328 ();
 b15zdnd11an1n64x5 FILLER_270_392 ();
 b15zdnd11an1n64x5 FILLER_270_456 ();
 b15zdnd11an1n64x5 FILLER_270_520 ();
 b15zdnd11an1n64x5 FILLER_270_584 ();
 b15zdnd11an1n64x5 FILLER_270_648 ();
 b15zdnd11an1n04x5 FILLER_270_712 ();
 b15zdnd00an1n02x5 FILLER_270_716 ();
 b15zdnd11an1n64x5 FILLER_270_726 ();
 b15zdnd11an1n64x5 FILLER_270_790 ();
 b15zdnd11an1n64x5 FILLER_270_854 ();
 b15zdnd11an1n64x5 FILLER_270_918 ();
 b15zdnd11an1n64x5 FILLER_270_982 ();
 b15zdnd11an1n64x5 FILLER_270_1046 ();
 b15zdnd11an1n64x5 FILLER_270_1110 ();
 b15zdnd11an1n64x5 FILLER_270_1174 ();
 b15zdnd11an1n64x5 FILLER_270_1238 ();
 b15zdnd11an1n64x5 FILLER_270_1302 ();
 b15zdnd11an1n64x5 FILLER_270_1366 ();
 b15zdnd11an1n64x5 FILLER_270_1430 ();
 b15zdnd11an1n64x5 FILLER_270_1494 ();
 b15zdnd11an1n64x5 FILLER_270_1558 ();
 b15zdnd11an1n64x5 FILLER_270_1622 ();
 b15zdnd11an1n64x5 FILLER_270_1686 ();
 b15zdnd11an1n64x5 FILLER_270_1750 ();
 b15zdnd11an1n64x5 FILLER_270_1814 ();
 b15zdnd11an1n64x5 FILLER_270_1878 ();
 b15zdnd11an1n64x5 FILLER_270_1942 ();
 b15zdnd11an1n64x5 FILLER_270_2006 ();
 b15zdnd11an1n64x5 FILLER_270_2070 ();
 b15zdnd11an1n16x5 FILLER_270_2134 ();
 b15zdnd11an1n04x5 FILLER_270_2150 ();
 b15zdnd11an1n64x5 FILLER_270_2162 ();
 b15zdnd11an1n32x5 FILLER_270_2226 ();
 b15zdnd11an1n16x5 FILLER_270_2258 ();
 b15zdnd00an1n02x5 FILLER_270_2274 ();
 b15zdnd11an1n64x5 FILLER_271_0 ();
 b15zdnd11an1n64x5 FILLER_271_64 ();
 b15zdnd11an1n64x5 FILLER_271_128 ();
 b15zdnd11an1n64x5 FILLER_271_192 ();
 b15zdnd11an1n64x5 FILLER_271_256 ();
 b15zdnd11an1n64x5 FILLER_271_320 ();
 b15zdnd11an1n64x5 FILLER_271_384 ();
 b15zdnd11an1n64x5 FILLER_271_448 ();
 b15zdnd11an1n64x5 FILLER_271_512 ();
 b15zdnd11an1n64x5 FILLER_271_576 ();
 b15zdnd11an1n64x5 FILLER_271_640 ();
 b15zdnd11an1n64x5 FILLER_271_704 ();
 b15zdnd11an1n64x5 FILLER_271_768 ();
 b15zdnd11an1n64x5 FILLER_271_832 ();
 b15zdnd11an1n64x5 FILLER_271_896 ();
 b15zdnd11an1n64x5 FILLER_271_960 ();
 b15zdnd11an1n64x5 FILLER_271_1024 ();
 b15zdnd11an1n64x5 FILLER_271_1088 ();
 b15zdnd11an1n64x5 FILLER_271_1152 ();
 b15zdnd11an1n64x5 FILLER_271_1216 ();
 b15zdnd11an1n64x5 FILLER_271_1280 ();
 b15zdnd11an1n64x5 FILLER_271_1344 ();
 b15zdnd11an1n64x5 FILLER_271_1408 ();
 b15zdnd11an1n64x5 FILLER_271_1472 ();
 b15zdnd11an1n64x5 FILLER_271_1536 ();
 b15zdnd11an1n64x5 FILLER_271_1600 ();
 b15zdnd11an1n64x5 FILLER_271_1664 ();
 b15zdnd11an1n64x5 FILLER_271_1728 ();
 b15zdnd11an1n64x5 FILLER_271_1792 ();
 b15zdnd11an1n64x5 FILLER_271_1856 ();
 b15zdnd11an1n64x5 FILLER_271_1920 ();
 b15zdnd11an1n64x5 FILLER_271_1984 ();
 b15zdnd11an1n64x5 FILLER_271_2048 ();
 b15zdnd11an1n64x5 FILLER_271_2112 ();
 b15zdnd11an1n64x5 FILLER_271_2176 ();
 b15zdnd11an1n32x5 FILLER_271_2240 ();
 b15zdnd11an1n08x5 FILLER_271_2272 ();
 b15zdnd11an1n04x5 FILLER_271_2280 ();
 b15zdnd11an1n64x5 FILLER_272_8 ();
 b15zdnd11an1n64x5 FILLER_272_72 ();
 b15zdnd11an1n64x5 FILLER_272_136 ();
 b15zdnd11an1n64x5 FILLER_272_200 ();
 b15zdnd11an1n64x5 FILLER_272_264 ();
 b15zdnd11an1n64x5 FILLER_272_328 ();
 b15zdnd11an1n64x5 FILLER_272_392 ();
 b15zdnd11an1n64x5 FILLER_272_456 ();
 b15zdnd11an1n64x5 FILLER_272_520 ();
 b15zdnd11an1n64x5 FILLER_272_584 ();
 b15zdnd11an1n64x5 FILLER_272_648 ();
 b15zdnd11an1n04x5 FILLER_272_712 ();
 b15zdnd00an1n02x5 FILLER_272_716 ();
 b15zdnd11an1n64x5 FILLER_272_726 ();
 b15zdnd11an1n64x5 FILLER_272_790 ();
 b15zdnd11an1n64x5 FILLER_272_854 ();
 b15zdnd11an1n64x5 FILLER_272_918 ();
 b15zdnd11an1n64x5 FILLER_272_982 ();
 b15zdnd11an1n64x5 FILLER_272_1046 ();
 b15zdnd11an1n64x5 FILLER_272_1110 ();
 b15zdnd11an1n64x5 FILLER_272_1174 ();
 b15zdnd11an1n64x5 FILLER_272_1238 ();
 b15zdnd11an1n64x5 FILLER_272_1302 ();
 b15zdnd11an1n64x5 FILLER_272_1366 ();
 b15zdnd11an1n64x5 FILLER_272_1430 ();
 b15zdnd11an1n64x5 FILLER_272_1494 ();
 b15zdnd11an1n64x5 FILLER_272_1558 ();
 b15zdnd11an1n64x5 FILLER_272_1622 ();
 b15zdnd11an1n64x5 FILLER_272_1686 ();
 b15zdnd11an1n64x5 FILLER_272_1750 ();
 b15zdnd11an1n64x5 FILLER_272_1814 ();
 b15zdnd11an1n64x5 FILLER_272_1878 ();
 b15zdnd11an1n64x5 FILLER_272_1942 ();
 b15zdnd11an1n64x5 FILLER_272_2006 ();
 b15zdnd11an1n64x5 FILLER_272_2070 ();
 b15zdnd11an1n16x5 FILLER_272_2134 ();
 b15zdnd11an1n04x5 FILLER_272_2150 ();
 b15zdnd11an1n64x5 FILLER_272_2162 ();
 b15zdnd11an1n32x5 FILLER_272_2226 ();
 b15zdnd11an1n16x5 FILLER_272_2258 ();
 b15zdnd00an1n02x5 FILLER_272_2274 ();
 b15zdnd11an1n64x5 FILLER_273_0 ();
 b15zdnd11an1n64x5 FILLER_273_64 ();
 b15zdnd11an1n64x5 FILLER_273_128 ();
 b15zdnd11an1n64x5 FILLER_273_192 ();
 b15zdnd11an1n64x5 FILLER_273_256 ();
 b15zdnd11an1n64x5 FILLER_273_320 ();
 b15zdnd11an1n64x5 FILLER_273_384 ();
 b15zdnd11an1n64x5 FILLER_273_448 ();
 b15zdnd11an1n64x5 FILLER_273_512 ();
 b15zdnd11an1n64x5 FILLER_273_576 ();
 b15zdnd11an1n64x5 FILLER_273_640 ();
 b15zdnd11an1n64x5 FILLER_273_704 ();
 b15zdnd11an1n64x5 FILLER_273_768 ();
 b15zdnd11an1n64x5 FILLER_273_832 ();
 b15zdnd11an1n64x5 FILLER_273_896 ();
 b15zdnd11an1n64x5 FILLER_273_960 ();
 b15zdnd11an1n64x5 FILLER_273_1024 ();
 b15zdnd11an1n64x5 FILLER_273_1088 ();
 b15zdnd11an1n64x5 FILLER_273_1152 ();
 b15zdnd11an1n64x5 FILLER_273_1216 ();
 b15zdnd11an1n64x5 FILLER_273_1280 ();
 b15zdnd11an1n64x5 FILLER_273_1344 ();
 b15zdnd11an1n64x5 FILLER_273_1408 ();
 b15zdnd11an1n64x5 FILLER_273_1472 ();
 b15zdnd11an1n64x5 FILLER_273_1536 ();
 b15zdnd11an1n64x5 FILLER_273_1600 ();
 b15zdnd11an1n64x5 FILLER_273_1664 ();
 b15zdnd11an1n64x5 FILLER_273_1728 ();
 b15zdnd11an1n64x5 FILLER_273_1792 ();
 b15zdnd11an1n64x5 FILLER_273_1856 ();
 b15zdnd11an1n64x5 FILLER_273_1920 ();
 b15zdnd11an1n64x5 FILLER_273_1984 ();
 b15zdnd11an1n64x5 FILLER_273_2048 ();
 b15zdnd11an1n64x5 FILLER_273_2112 ();
 b15zdnd11an1n64x5 FILLER_273_2176 ();
 b15zdnd11an1n32x5 FILLER_273_2240 ();
 b15zdnd11an1n08x5 FILLER_273_2272 ();
 b15zdnd11an1n04x5 FILLER_273_2280 ();
 b15zdnd11an1n64x5 FILLER_274_8 ();
 b15zdnd11an1n64x5 FILLER_274_72 ();
 b15zdnd11an1n64x5 FILLER_274_136 ();
 b15zdnd11an1n64x5 FILLER_274_200 ();
 b15zdnd11an1n64x5 FILLER_274_264 ();
 b15zdnd11an1n64x5 FILLER_274_328 ();
 b15zdnd11an1n64x5 FILLER_274_392 ();
 b15zdnd11an1n64x5 FILLER_274_456 ();
 b15zdnd11an1n64x5 FILLER_274_520 ();
 b15zdnd11an1n64x5 FILLER_274_584 ();
 b15zdnd11an1n64x5 FILLER_274_648 ();
 b15zdnd11an1n04x5 FILLER_274_712 ();
 b15zdnd00an1n02x5 FILLER_274_716 ();
 b15zdnd11an1n64x5 FILLER_274_726 ();
 b15zdnd11an1n64x5 FILLER_274_790 ();
 b15zdnd11an1n64x5 FILLER_274_854 ();
 b15zdnd11an1n64x5 FILLER_274_918 ();
 b15zdnd11an1n64x5 FILLER_274_982 ();
 b15zdnd11an1n64x5 FILLER_274_1046 ();
 b15zdnd11an1n64x5 FILLER_274_1110 ();
 b15zdnd11an1n64x5 FILLER_274_1174 ();
 b15zdnd11an1n64x5 FILLER_274_1238 ();
 b15zdnd11an1n64x5 FILLER_274_1302 ();
 b15zdnd11an1n64x5 FILLER_274_1366 ();
 b15zdnd11an1n64x5 FILLER_274_1430 ();
 b15zdnd11an1n64x5 FILLER_274_1494 ();
 b15zdnd11an1n64x5 FILLER_274_1558 ();
 b15zdnd11an1n64x5 FILLER_274_1622 ();
 b15zdnd11an1n64x5 FILLER_274_1686 ();
 b15zdnd11an1n64x5 FILLER_274_1750 ();
 b15zdnd11an1n64x5 FILLER_274_1814 ();
 b15zdnd11an1n64x5 FILLER_274_1878 ();
 b15zdnd11an1n64x5 FILLER_274_1942 ();
 b15zdnd11an1n64x5 FILLER_274_2006 ();
 b15zdnd11an1n64x5 FILLER_274_2070 ();
 b15zdnd11an1n16x5 FILLER_274_2134 ();
 b15zdnd11an1n04x5 FILLER_274_2150 ();
 b15zdnd11an1n64x5 FILLER_274_2162 ();
 b15zdnd11an1n32x5 FILLER_274_2226 ();
 b15zdnd11an1n16x5 FILLER_274_2258 ();
 b15zdnd00an1n02x5 FILLER_274_2274 ();
 b15zdnd11an1n64x5 FILLER_275_0 ();
 b15zdnd11an1n64x5 FILLER_275_64 ();
 b15zdnd11an1n64x5 FILLER_275_128 ();
 b15zdnd11an1n64x5 FILLER_275_192 ();
 b15zdnd11an1n64x5 FILLER_275_256 ();
 b15zdnd11an1n64x5 FILLER_275_320 ();
 b15zdnd11an1n64x5 FILLER_275_384 ();
 b15zdnd11an1n64x5 FILLER_275_448 ();
 b15zdnd11an1n64x5 FILLER_275_512 ();
 b15zdnd11an1n64x5 FILLER_275_576 ();
 b15zdnd11an1n64x5 FILLER_275_640 ();
 b15zdnd11an1n64x5 FILLER_275_704 ();
 b15zdnd11an1n64x5 FILLER_275_768 ();
 b15zdnd11an1n64x5 FILLER_275_832 ();
 b15zdnd11an1n64x5 FILLER_275_896 ();
 b15zdnd11an1n64x5 FILLER_275_960 ();
 b15zdnd11an1n64x5 FILLER_275_1024 ();
 b15zdnd11an1n64x5 FILLER_275_1088 ();
 b15zdnd11an1n64x5 FILLER_275_1152 ();
 b15zdnd11an1n64x5 FILLER_275_1216 ();
 b15zdnd11an1n64x5 FILLER_275_1280 ();
 b15zdnd11an1n64x5 FILLER_275_1344 ();
 b15zdnd11an1n64x5 FILLER_275_1408 ();
 b15zdnd11an1n64x5 FILLER_275_1472 ();
 b15zdnd11an1n64x5 FILLER_275_1536 ();
 b15zdnd11an1n64x5 FILLER_275_1600 ();
 b15zdnd11an1n64x5 FILLER_275_1664 ();
 b15zdnd11an1n64x5 FILLER_275_1728 ();
 b15zdnd11an1n64x5 FILLER_275_1792 ();
 b15zdnd11an1n64x5 FILLER_275_1856 ();
 b15zdnd11an1n64x5 FILLER_275_1920 ();
 b15zdnd11an1n64x5 FILLER_275_1984 ();
 b15zdnd11an1n64x5 FILLER_275_2048 ();
 b15zdnd11an1n64x5 FILLER_275_2112 ();
 b15zdnd11an1n64x5 FILLER_275_2176 ();
 b15zdnd11an1n32x5 FILLER_275_2240 ();
 b15zdnd11an1n08x5 FILLER_275_2272 ();
 b15zdnd11an1n04x5 FILLER_275_2280 ();
 b15zdnd11an1n64x5 FILLER_276_8 ();
 b15zdnd11an1n64x5 FILLER_276_72 ();
 b15zdnd11an1n64x5 FILLER_276_136 ();
 b15zdnd11an1n64x5 FILLER_276_200 ();
 b15zdnd11an1n64x5 FILLER_276_264 ();
 b15zdnd11an1n64x5 FILLER_276_328 ();
 b15zdnd11an1n64x5 FILLER_276_392 ();
 b15zdnd11an1n64x5 FILLER_276_456 ();
 b15zdnd11an1n64x5 FILLER_276_520 ();
 b15zdnd11an1n64x5 FILLER_276_584 ();
 b15zdnd11an1n64x5 FILLER_276_648 ();
 b15zdnd11an1n04x5 FILLER_276_712 ();
 b15zdnd00an1n02x5 FILLER_276_716 ();
 b15zdnd11an1n64x5 FILLER_276_726 ();
 b15zdnd11an1n64x5 FILLER_276_790 ();
 b15zdnd11an1n64x5 FILLER_276_854 ();
 b15zdnd11an1n64x5 FILLER_276_918 ();
 b15zdnd11an1n64x5 FILLER_276_982 ();
 b15zdnd11an1n64x5 FILLER_276_1046 ();
 b15zdnd11an1n64x5 FILLER_276_1110 ();
 b15zdnd11an1n64x5 FILLER_276_1174 ();
 b15zdnd11an1n64x5 FILLER_276_1238 ();
 b15zdnd11an1n64x5 FILLER_276_1302 ();
 b15zdnd11an1n64x5 FILLER_276_1366 ();
 b15zdnd11an1n64x5 FILLER_276_1430 ();
 b15zdnd11an1n64x5 FILLER_276_1494 ();
 b15zdnd11an1n64x5 FILLER_276_1558 ();
 b15zdnd11an1n64x5 FILLER_276_1622 ();
 b15zdnd11an1n64x5 FILLER_276_1686 ();
 b15zdnd11an1n64x5 FILLER_276_1750 ();
 b15zdnd11an1n64x5 FILLER_276_1814 ();
 b15zdnd11an1n64x5 FILLER_276_1878 ();
 b15zdnd11an1n64x5 FILLER_276_1942 ();
 b15zdnd11an1n64x5 FILLER_276_2006 ();
 b15zdnd11an1n64x5 FILLER_276_2070 ();
 b15zdnd11an1n16x5 FILLER_276_2134 ();
 b15zdnd11an1n04x5 FILLER_276_2150 ();
 b15zdnd11an1n64x5 FILLER_276_2162 ();
 b15zdnd11an1n32x5 FILLER_276_2226 ();
 b15zdnd11an1n16x5 FILLER_276_2258 ();
 b15zdnd00an1n02x5 FILLER_276_2274 ();
 b15zdnd11an1n64x5 FILLER_277_0 ();
 b15zdnd11an1n64x5 FILLER_277_64 ();
 b15zdnd11an1n64x5 FILLER_277_128 ();
 b15zdnd11an1n64x5 FILLER_277_192 ();
 b15zdnd11an1n64x5 FILLER_277_256 ();
 b15zdnd11an1n64x5 FILLER_277_320 ();
 b15zdnd11an1n64x5 FILLER_277_384 ();
 b15zdnd11an1n64x5 FILLER_277_448 ();
 b15zdnd11an1n64x5 FILLER_277_512 ();
 b15zdnd11an1n64x5 FILLER_277_576 ();
 b15zdnd11an1n64x5 FILLER_277_640 ();
 b15zdnd11an1n64x5 FILLER_277_704 ();
 b15zdnd11an1n64x5 FILLER_277_768 ();
 b15zdnd11an1n64x5 FILLER_277_832 ();
 b15zdnd11an1n64x5 FILLER_277_896 ();
 b15zdnd11an1n64x5 FILLER_277_960 ();
 b15zdnd11an1n64x5 FILLER_277_1024 ();
 b15zdnd11an1n64x5 FILLER_277_1088 ();
 b15zdnd11an1n64x5 FILLER_277_1152 ();
 b15zdnd11an1n64x5 FILLER_277_1216 ();
 b15zdnd11an1n64x5 FILLER_277_1280 ();
 b15zdnd11an1n64x5 FILLER_277_1344 ();
 b15zdnd11an1n64x5 FILLER_277_1408 ();
 b15zdnd11an1n64x5 FILLER_277_1472 ();
 b15zdnd11an1n64x5 FILLER_277_1536 ();
 b15zdnd11an1n64x5 FILLER_277_1600 ();
 b15zdnd11an1n64x5 FILLER_277_1664 ();
 b15zdnd11an1n64x5 FILLER_277_1728 ();
 b15zdnd11an1n64x5 FILLER_277_1792 ();
 b15zdnd11an1n64x5 FILLER_277_1856 ();
 b15zdnd11an1n64x5 FILLER_277_1920 ();
 b15zdnd11an1n64x5 FILLER_277_1984 ();
 b15zdnd11an1n64x5 FILLER_277_2048 ();
 b15zdnd11an1n64x5 FILLER_277_2112 ();
 b15zdnd11an1n64x5 FILLER_277_2176 ();
 b15zdnd11an1n32x5 FILLER_277_2240 ();
 b15zdnd11an1n08x5 FILLER_277_2272 ();
 b15zdnd11an1n04x5 FILLER_277_2280 ();
 b15zdnd11an1n64x5 FILLER_278_8 ();
 b15zdnd11an1n64x5 FILLER_278_72 ();
 b15zdnd11an1n64x5 FILLER_278_136 ();
 b15zdnd11an1n64x5 FILLER_278_200 ();
 b15zdnd11an1n64x5 FILLER_278_264 ();
 b15zdnd11an1n64x5 FILLER_278_328 ();
 b15zdnd11an1n64x5 FILLER_278_392 ();
 b15zdnd11an1n64x5 FILLER_278_456 ();
 b15zdnd11an1n64x5 FILLER_278_520 ();
 b15zdnd11an1n64x5 FILLER_278_584 ();
 b15zdnd11an1n64x5 FILLER_278_648 ();
 b15zdnd11an1n04x5 FILLER_278_712 ();
 b15zdnd00an1n02x5 FILLER_278_716 ();
 b15zdnd11an1n64x5 FILLER_278_726 ();
 b15zdnd11an1n64x5 FILLER_278_790 ();
 b15zdnd11an1n64x5 FILLER_278_854 ();
 b15zdnd11an1n64x5 FILLER_278_918 ();
 b15zdnd11an1n64x5 FILLER_278_982 ();
 b15zdnd11an1n64x5 FILLER_278_1046 ();
 b15zdnd11an1n64x5 FILLER_278_1110 ();
 b15zdnd11an1n64x5 FILLER_278_1174 ();
 b15zdnd11an1n64x5 FILLER_278_1238 ();
 b15zdnd11an1n64x5 FILLER_278_1302 ();
 b15zdnd11an1n64x5 FILLER_278_1366 ();
 b15zdnd11an1n64x5 FILLER_278_1430 ();
 b15zdnd11an1n64x5 FILLER_278_1494 ();
 b15zdnd11an1n64x5 FILLER_278_1558 ();
 b15zdnd11an1n64x5 FILLER_278_1622 ();
 b15zdnd11an1n64x5 FILLER_278_1686 ();
 b15zdnd11an1n64x5 FILLER_278_1750 ();
 b15zdnd11an1n64x5 FILLER_278_1814 ();
 b15zdnd11an1n64x5 FILLER_278_1878 ();
 b15zdnd11an1n64x5 FILLER_278_1942 ();
 b15zdnd11an1n64x5 FILLER_278_2006 ();
 b15zdnd11an1n64x5 FILLER_278_2070 ();
 b15zdnd11an1n16x5 FILLER_278_2134 ();
 b15zdnd11an1n04x5 FILLER_278_2150 ();
 b15zdnd11an1n64x5 FILLER_278_2162 ();
 b15zdnd11an1n32x5 FILLER_278_2226 ();
 b15zdnd11an1n16x5 FILLER_278_2258 ();
 b15zdnd00an1n02x5 FILLER_278_2274 ();
 b15zdnd11an1n64x5 FILLER_279_0 ();
 b15zdnd11an1n64x5 FILLER_279_64 ();
 b15zdnd11an1n64x5 FILLER_279_128 ();
 b15zdnd11an1n64x5 FILLER_279_192 ();
 b15zdnd11an1n64x5 FILLER_279_256 ();
 b15zdnd11an1n64x5 FILLER_279_320 ();
 b15zdnd11an1n64x5 FILLER_279_384 ();
 b15zdnd11an1n64x5 FILLER_279_448 ();
 b15zdnd11an1n64x5 FILLER_279_512 ();
 b15zdnd11an1n64x5 FILLER_279_576 ();
 b15zdnd11an1n64x5 FILLER_279_640 ();
 b15zdnd11an1n64x5 FILLER_279_704 ();
 b15zdnd11an1n64x5 FILLER_279_768 ();
 b15zdnd11an1n64x5 FILLER_279_832 ();
 b15zdnd11an1n64x5 FILLER_279_896 ();
 b15zdnd11an1n64x5 FILLER_279_960 ();
 b15zdnd11an1n64x5 FILLER_279_1024 ();
 b15zdnd11an1n64x5 FILLER_279_1088 ();
 b15zdnd11an1n64x5 FILLER_279_1152 ();
 b15zdnd11an1n64x5 FILLER_279_1216 ();
 b15zdnd11an1n64x5 FILLER_279_1280 ();
 b15zdnd11an1n64x5 FILLER_279_1344 ();
 b15zdnd11an1n64x5 FILLER_279_1408 ();
 b15zdnd11an1n64x5 FILLER_279_1472 ();
 b15zdnd11an1n64x5 FILLER_279_1536 ();
 b15zdnd11an1n64x5 FILLER_279_1600 ();
 b15zdnd11an1n64x5 FILLER_279_1664 ();
 b15zdnd11an1n64x5 FILLER_279_1728 ();
 b15zdnd11an1n64x5 FILLER_279_1792 ();
 b15zdnd11an1n64x5 FILLER_279_1856 ();
 b15zdnd11an1n64x5 FILLER_279_1920 ();
 b15zdnd11an1n64x5 FILLER_279_1984 ();
 b15zdnd11an1n64x5 FILLER_279_2048 ();
 b15zdnd11an1n64x5 FILLER_279_2112 ();
 b15zdnd11an1n64x5 FILLER_279_2176 ();
 b15zdnd11an1n32x5 FILLER_279_2240 ();
 b15zdnd11an1n08x5 FILLER_279_2272 ();
 b15zdnd11an1n04x5 FILLER_279_2280 ();
 b15zdnd11an1n64x5 FILLER_280_8 ();
 b15zdnd11an1n64x5 FILLER_280_72 ();
 b15zdnd11an1n64x5 FILLER_280_136 ();
 b15zdnd11an1n64x5 FILLER_280_200 ();
 b15zdnd11an1n64x5 FILLER_280_264 ();
 b15zdnd11an1n64x5 FILLER_280_328 ();
 b15zdnd11an1n64x5 FILLER_280_392 ();
 b15zdnd11an1n64x5 FILLER_280_456 ();
 b15zdnd11an1n64x5 FILLER_280_520 ();
 b15zdnd11an1n64x5 FILLER_280_584 ();
 b15zdnd11an1n64x5 FILLER_280_648 ();
 b15zdnd11an1n04x5 FILLER_280_712 ();
 b15zdnd00an1n02x5 FILLER_280_716 ();
 b15zdnd11an1n64x5 FILLER_280_726 ();
 b15zdnd11an1n64x5 FILLER_280_790 ();
 b15zdnd11an1n64x5 FILLER_280_854 ();
 b15zdnd11an1n64x5 FILLER_280_918 ();
 b15zdnd11an1n64x5 FILLER_280_982 ();
 b15zdnd11an1n64x5 FILLER_280_1046 ();
 b15zdnd11an1n64x5 FILLER_280_1110 ();
 b15zdnd11an1n64x5 FILLER_280_1174 ();
 b15zdnd11an1n64x5 FILLER_280_1238 ();
 b15zdnd11an1n64x5 FILLER_280_1302 ();
 b15zdnd11an1n64x5 FILLER_280_1366 ();
 b15zdnd11an1n64x5 FILLER_280_1430 ();
 b15zdnd11an1n64x5 FILLER_280_1494 ();
 b15zdnd11an1n64x5 FILLER_280_1558 ();
 b15zdnd11an1n64x5 FILLER_280_1622 ();
 b15zdnd11an1n64x5 FILLER_280_1686 ();
 b15zdnd11an1n64x5 FILLER_280_1750 ();
 b15zdnd11an1n64x5 FILLER_280_1814 ();
 b15zdnd11an1n64x5 FILLER_280_1878 ();
 b15zdnd11an1n64x5 FILLER_280_1942 ();
 b15zdnd11an1n64x5 FILLER_280_2006 ();
 b15zdnd11an1n64x5 FILLER_280_2070 ();
 b15zdnd11an1n16x5 FILLER_280_2134 ();
 b15zdnd11an1n04x5 FILLER_280_2150 ();
 b15zdnd11an1n64x5 FILLER_280_2162 ();
 b15zdnd11an1n32x5 FILLER_280_2226 ();
 b15zdnd11an1n16x5 FILLER_280_2258 ();
 b15zdnd00an1n02x5 FILLER_280_2274 ();
 b15zdnd11an1n64x5 FILLER_281_0 ();
 b15zdnd11an1n64x5 FILLER_281_64 ();
 b15zdnd11an1n64x5 FILLER_281_128 ();
 b15zdnd11an1n64x5 FILLER_281_192 ();
 b15zdnd11an1n64x5 FILLER_281_256 ();
 b15zdnd11an1n64x5 FILLER_281_320 ();
 b15zdnd11an1n64x5 FILLER_281_384 ();
 b15zdnd11an1n64x5 FILLER_281_448 ();
 b15zdnd11an1n64x5 FILLER_281_512 ();
 b15zdnd11an1n64x5 FILLER_281_576 ();
 b15zdnd11an1n64x5 FILLER_281_640 ();
 b15zdnd11an1n64x5 FILLER_281_704 ();
 b15zdnd11an1n64x5 FILLER_281_768 ();
 b15zdnd11an1n64x5 FILLER_281_832 ();
 b15zdnd11an1n64x5 FILLER_281_896 ();
 b15zdnd11an1n64x5 FILLER_281_960 ();
 b15zdnd11an1n64x5 FILLER_281_1024 ();
 b15zdnd11an1n64x5 FILLER_281_1088 ();
 b15zdnd11an1n64x5 FILLER_281_1152 ();
 b15zdnd11an1n64x5 FILLER_281_1216 ();
 b15zdnd11an1n64x5 FILLER_281_1280 ();
 b15zdnd11an1n64x5 FILLER_281_1344 ();
 b15zdnd11an1n64x5 FILLER_281_1408 ();
 b15zdnd11an1n64x5 FILLER_281_1472 ();
 b15zdnd11an1n64x5 FILLER_281_1536 ();
 b15zdnd11an1n64x5 FILLER_281_1600 ();
 b15zdnd11an1n64x5 FILLER_281_1664 ();
 b15zdnd11an1n64x5 FILLER_281_1728 ();
 b15zdnd11an1n64x5 FILLER_281_1792 ();
 b15zdnd11an1n64x5 FILLER_281_1856 ();
 b15zdnd11an1n64x5 FILLER_281_1920 ();
 b15zdnd11an1n64x5 FILLER_281_1984 ();
 b15zdnd11an1n64x5 FILLER_281_2048 ();
 b15zdnd11an1n64x5 FILLER_281_2112 ();
 b15zdnd11an1n64x5 FILLER_281_2176 ();
 b15zdnd11an1n32x5 FILLER_281_2240 ();
 b15zdnd11an1n08x5 FILLER_281_2272 ();
 b15zdnd11an1n04x5 FILLER_281_2280 ();
 b15zdnd11an1n64x5 FILLER_282_8 ();
 b15zdnd11an1n64x5 FILLER_282_72 ();
 b15zdnd11an1n64x5 FILLER_282_136 ();
 b15zdnd11an1n64x5 FILLER_282_200 ();
 b15zdnd11an1n64x5 FILLER_282_264 ();
 b15zdnd11an1n64x5 FILLER_282_328 ();
 b15zdnd11an1n64x5 FILLER_282_392 ();
 b15zdnd11an1n64x5 FILLER_282_456 ();
 b15zdnd11an1n64x5 FILLER_282_520 ();
 b15zdnd11an1n64x5 FILLER_282_584 ();
 b15zdnd11an1n64x5 FILLER_282_648 ();
 b15zdnd11an1n04x5 FILLER_282_712 ();
 b15zdnd00an1n02x5 FILLER_282_716 ();
 b15zdnd11an1n64x5 FILLER_282_726 ();
 b15zdnd11an1n64x5 FILLER_282_790 ();
 b15zdnd11an1n64x5 FILLER_282_854 ();
 b15zdnd11an1n64x5 FILLER_282_918 ();
 b15zdnd11an1n64x5 FILLER_282_982 ();
 b15zdnd11an1n64x5 FILLER_282_1046 ();
 b15zdnd11an1n64x5 FILLER_282_1110 ();
 b15zdnd11an1n64x5 FILLER_282_1174 ();
 b15zdnd11an1n64x5 FILLER_282_1238 ();
 b15zdnd11an1n64x5 FILLER_282_1302 ();
 b15zdnd11an1n64x5 FILLER_282_1366 ();
 b15zdnd11an1n64x5 FILLER_282_1430 ();
 b15zdnd11an1n64x5 FILLER_282_1494 ();
 b15zdnd11an1n64x5 FILLER_282_1558 ();
 b15zdnd11an1n64x5 FILLER_282_1622 ();
 b15zdnd11an1n64x5 FILLER_282_1686 ();
 b15zdnd11an1n64x5 FILLER_282_1750 ();
 b15zdnd11an1n64x5 FILLER_282_1814 ();
 b15zdnd11an1n64x5 FILLER_282_1878 ();
 b15zdnd11an1n64x5 FILLER_282_1942 ();
 b15zdnd11an1n64x5 FILLER_282_2006 ();
 b15zdnd11an1n64x5 FILLER_282_2070 ();
 b15zdnd11an1n16x5 FILLER_282_2134 ();
 b15zdnd11an1n04x5 FILLER_282_2150 ();
 b15zdnd11an1n64x5 FILLER_282_2162 ();
 b15zdnd11an1n32x5 FILLER_282_2226 ();
 b15zdnd11an1n16x5 FILLER_282_2258 ();
 b15zdnd00an1n02x5 FILLER_282_2274 ();
 b15zdnd11an1n64x5 FILLER_283_0 ();
 b15zdnd11an1n64x5 FILLER_283_64 ();
 b15zdnd11an1n64x5 FILLER_283_128 ();
 b15zdnd11an1n64x5 FILLER_283_192 ();
 b15zdnd11an1n64x5 FILLER_283_256 ();
 b15zdnd11an1n64x5 FILLER_283_320 ();
 b15zdnd11an1n64x5 FILLER_283_384 ();
 b15zdnd11an1n64x5 FILLER_283_448 ();
 b15zdnd11an1n64x5 FILLER_283_512 ();
 b15zdnd11an1n64x5 FILLER_283_576 ();
 b15zdnd11an1n64x5 FILLER_283_640 ();
 b15zdnd11an1n64x5 FILLER_283_704 ();
 b15zdnd11an1n64x5 FILLER_283_768 ();
 b15zdnd11an1n64x5 FILLER_283_832 ();
 b15zdnd11an1n64x5 FILLER_283_896 ();
 b15zdnd11an1n64x5 FILLER_283_960 ();
 b15zdnd11an1n64x5 FILLER_283_1024 ();
 b15zdnd11an1n64x5 FILLER_283_1088 ();
 b15zdnd11an1n64x5 FILLER_283_1152 ();
 b15zdnd11an1n64x5 FILLER_283_1216 ();
 b15zdnd11an1n64x5 FILLER_283_1280 ();
 b15zdnd11an1n64x5 FILLER_283_1344 ();
 b15zdnd11an1n64x5 FILLER_283_1408 ();
 b15zdnd11an1n64x5 FILLER_283_1472 ();
 b15zdnd11an1n64x5 FILLER_283_1536 ();
 b15zdnd11an1n64x5 FILLER_283_1600 ();
 b15zdnd11an1n64x5 FILLER_283_1664 ();
 b15zdnd11an1n64x5 FILLER_283_1728 ();
 b15zdnd11an1n64x5 FILLER_283_1792 ();
 b15zdnd11an1n64x5 FILLER_283_1856 ();
 b15zdnd11an1n64x5 FILLER_283_1920 ();
 b15zdnd11an1n64x5 FILLER_283_1984 ();
 b15zdnd11an1n64x5 FILLER_283_2048 ();
 b15zdnd11an1n64x5 FILLER_283_2112 ();
 b15zdnd11an1n64x5 FILLER_283_2176 ();
 b15zdnd11an1n32x5 FILLER_283_2240 ();
 b15zdnd11an1n08x5 FILLER_283_2272 ();
 b15zdnd11an1n04x5 FILLER_283_2280 ();
 b15zdnd11an1n64x5 FILLER_284_8 ();
 b15zdnd11an1n64x5 FILLER_284_72 ();
 b15zdnd11an1n64x5 FILLER_284_136 ();
 b15zdnd11an1n64x5 FILLER_284_200 ();
 b15zdnd11an1n64x5 FILLER_284_264 ();
 b15zdnd11an1n64x5 FILLER_284_328 ();
 b15zdnd11an1n64x5 FILLER_284_392 ();
 b15zdnd11an1n64x5 FILLER_284_456 ();
 b15zdnd11an1n64x5 FILLER_284_520 ();
 b15zdnd11an1n64x5 FILLER_284_584 ();
 b15zdnd11an1n64x5 FILLER_284_648 ();
 b15zdnd11an1n04x5 FILLER_284_712 ();
 b15zdnd00an1n02x5 FILLER_284_716 ();
 b15zdnd11an1n64x5 FILLER_284_726 ();
 b15zdnd11an1n64x5 FILLER_284_790 ();
 b15zdnd11an1n64x5 FILLER_284_854 ();
 b15zdnd11an1n64x5 FILLER_284_918 ();
 b15zdnd11an1n64x5 FILLER_284_982 ();
 b15zdnd11an1n64x5 FILLER_284_1046 ();
 b15zdnd11an1n64x5 FILLER_284_1110 ();
 b15zdnd11an1n64x5 FILLER_284_1174 ();
 b15zdnd11an1n64x5 FILLER_284_1238 ();
 b15zdnd11an1n64x5 FILLER_284_1302 ();
 b15zdnd11an1n64x5 FILLER_284_1366 ();
 b15zdnd11an1n64x5 FILLER_284_1430 ();
 b15zdnd11an1n64x5 FILLER_284_1494 ();
 b15zdnd11an1n64x5 FILLER_284_1558 ();
 b15zdnd11an1n64x5 FILLER_284_1622 ();
 b15zdnd11an1n64x5 FILLER_284_1686 ();
 b15zdnd11an1n64x5 FILLER_284_1750 ();
 b15zdnd11an1n64x5 FILLER_284_1814 ();
 b15zdnd11an1n64x5 FILLER_284_1878 ();
 b15zdnd11an1n64x5 FILLER_284_1942 ();
 b15zdnd11an1n64x5 FILLER_284_2006 ();
 b15zdnd11an1n64x5 FILLER_284_2070 ();
 b15zdnd11an1n16x5 FILLER_284_2134 ();
 b15zdnd11an1n04x5 FILLER_284_2150 ();
 b15zdnd11an1n64x5 FILLER_284_2162 ();
 b15zdnd11an1n32x5 FILLER_284_2226 ();
 b15zdnd11an1n16x5 FILLER_284_2258 ();
 b15zdnd00an1n02x5 FILLER_284_2274 ();
 b15zdnd11an1n64x5 FILLER_285_0 ();
 b15zdnd11an1n64x5 FILLER_285_64 ();
 b15zdnd11an1n64x5 FILLER_285_128 ();
 b15zdnd11an1n64x5 FILLER_285_192 ();
 b15zdnd11an1n64x5 FILLER_285_256 ();
 b15zdnd11an1n64x5 FILLER_285_320 ();
 b15zdnd11an1n64x5 FILLER_285_384 ();
 b15zdnd11an1n64x5 FILLER_285_448 ();
 b15zdnd11an1n64x5 FILLER_285_512 ();
 b15zdnd11an1n64x5 FILLER_285_576 ();
 b15zdnd11an1n64x5 FILLER_285_640 ();
 b15zdnd11an1n64x5 FILLER_285_704 ();
 b15zdnd11an1n64x5 FILLER_285_768 ();
 b15zdnd11an1n64x5 FILLER_285_832 ();
 b15zdnd11an1n64x5 FILLER_285_896 ();
 b15zdnd11an1n64x5 FILLER_285_960 ();
 b15zdnd11an1n64x5 FILLER_285_1024 ();
 b15zdnd11an1n64x5 FILLER_285_1088 ();
 b15zdnd11an1n64x5 FILLER_285_1152 ();
 b15zdnd11an1n64x5 FILLER_285_1216 ();
 b15zdnd11an1n64x5 FILLER_285_1280 ();
 b15zdnd11an1n64x5 FILLER_285_1344 ();
 b15zdnd11an1n64x5 FILLER_285_1408 ();
 b15zdnd11an1n64x5 FILLER_285_1472 ();
 b15zdnd11an1n64x5 FILLER_285_1536 ();
 b15zdnd11an1n64x5 FILLER_285_1600 ();
 b15zdnd11an1n64x5 FILLER_285_1664 ();
 b15zdnd11an1n64x5 FILLER_285_1728 ();
 b15zdnd11an1n64x5 FILLER_285_1792 ();
 b15zdnd11an1n64x5 FILLER_285_1856 ();
 b15zdnd11an1n64x5 FILLER_285_1920 ();
 b15zdnd11an1n64x5 FILLER_285_1984 ();
 b15zdnd11an1n64x5 FILLER_285_2048 ();
 b15zdnd11an1n64x5 FILLER_285_2112 ();
 b15zdnd11an1n64x5 FILLER_285_2176 ();
 b15zdnd11an1n32x5 FILLER_285_2240 ();
 b15zdnd11an1n08x5 FILLER_285_2272 ();
 b15zdnd11an1n04x5 FILLER_285_2280 ();
 b15zdnd11an1n64x5 FILLER_286_8 ();
 b15zdnd11an1n64x5 FILLER_286_72 ();
 b15zdnd11an1n64x5 FILLER_286_136 ();
 b15zdnd11an1n64x5 FILLER_286_200 ();
 b15zdnd11an1n64x5 FILLER_286_264 ();
 b15zdnd11an1n64x5 FILLER_286_328 ();
 b15zdnd11an1n64x5 FILLER_286_392 ();
 b15zdnd11an1n64x5 FILLER_286_456 ();
 b15zdnd11an1n64x5 FILLER_286_520 ();
 b15zdnd11an1n64x5 FILLER_286_584 ();
 b15zdnd11an1n64x5 FILLER_286_648 ();
 b15zdnd11an1n04x5 FILLER_286_712 ();
 b15zdnd00an1n02x5 FILLER_286_716 ();
 b15zdnd11an1n64x5 FILLER_286_726 ();
 b15zdnd11an1n64x5 FILLER_286_790 ();
 b15zdnd11an1n64x5 FILLER_286_854 ();
 b15zdnd11an1n64x5 FILLER_286_918 ();
 b15zdnd11an1n64x5 FILLER_286_982 ();
 b15zdnd11an1n64x5 FILLER_286_1046 ();
 b15zdnd11an1n64x5 FILLER_286_1110 ();
 b15zdnd11an1n64x5 FILLER_286_1174 ();
 b15zdnd11an1n64x5 FILLER_286_1238 ();
 b15zdnd11an1n64x5 FILLER_286_1302 ();
 b15zdnd11an1n64x5 FILLER_286_1366 ();
 b15zdnd11an1n64x5 FILLER_286_1430 ();
 b15zdnd11an1n64x5 FILLER_286_1494 ();
 b15zdnd11an1n64x5 FILLER_286_1558 ();
 b15zdnd11an1n64x5 FILLER_286_1622 ();
 b15zdnd11an1n64x5 FILLER_286_1686 ();
 b15zdnd11an1n64x5 FILLER_286_1750 ();
 b15zdnd11an1n64x5 FILLER_286_1814 ();
 b15zdnd11an1n64x5 FILLER_286_1878 ();
 b15zdnd11an1n64x5 FILLER_286_1942 ();
 b15zdnd11an1n64x5 FILLER_286_2006 ();
 b15zdnd11an1n64x5 FILLER_286_2070 ();
 b15zdnd11an1n16x5 FILLER_286_2134 ();
 b15zdnd11an1n04x5 FILLER_286_2150 ();
 b15zdnd11an1n64x5 FILLER_286_2162 ();
 b15zdnd11an1n32x5 FILLER_286_2226 ();
 b15zdnd11an1n16x5 FILLER_286_2258 ();
 b15zdnd00an1n02x5 FILLER_286_2274 ();
 b15zdnd11an1n64x5 FILLER_287_0 ();
 b15zdnd11an1n64x5 FILLER_287_64 ();
 b15zdnd11an1n64x5 FILLER_287_128 ();
 b15zdnd11an1n64x5 FILLER_287_192 ();
 b15zdnd11an1n64x5 FILLER_287_256 ();
 b15zdnd11an1n64x5 FILLER_287_320 ();
 b15zdnd11an1n64x5 FILLER_287_384 ();
 b15zdnd11an1n64x5 FILLER_287_448 ();
 b15zdnd11an1n64x5 FILLER_287_512 ();
 b15zdnd11an1n64x5 FILLER_287_576 ();
 b15zdnd11an1n64x5 FILLER_287_640 ();
 b15zdnd11an1n64x5 FILLER_287_704 ();
 b15zdnd11an1n64x5 FILLER_287_768 ();
 b15zdnd11an1n64x5 FILLER_287_832 ();
 b15zdnd11an1n64x5 FILLER_287_896 ();
 b15zdnd11an1n64x5 FILLER_287_960 ();
 b15zdnd11an1n64x5 FILLER_287_1024 ();
 b15zdnd11an1n64x5 FILLER_287_1088 ();
 b15zdnd11an1n64x5 FILLER_287_1152 ();
 b15zdnd11an1n64x5 FILLER_287_1216 ();
 b15zdnd11an1n64x5 FILLER_287_1280 ();
 b15zdnd11an1n64x5 FILLER_287_1344 ();
 b15zdnd11an1n64x5 FILLER_287_1408 ();
 b15zdnd11an1n64x5 FILLER_287_1472 ();
 b15zdnd11an1n64x5 FILLER_287_1536 ();
 b15zdnd11an1n64x5 FILLER_287_1600 ();
 b15zdnd11an1n64x5 FILLER_287_1664 ();
 b15zdnd11an1n64x5 FILLER_287_1728 ();
 b15zdnd11an1n64x5 FILLER_287_1792 ();
 b15zdnd11an1n64x5 FILLER_287_1856 ();
 b15zdnd11an1n64x5 FILLER_287_1920 ();
 b15zdnd11an1n64x5 FILLER_287_1984 ();
 b15zdnd11an1n64x5 FILLER_287_2048 ();
 b15zdnd11an1n64x5 FILLER_287_2112 ();
 b15zdnd11an1n64x5 FILLER_287_2176 ();
 b15zdnd11an1n32x5 FILLER_287_2240 ();
 b15zdnd11an1n08x5 FILLER_287_2272 ();
 b15zdnd11an1n04x5 FILLER_287_2280 ();
 b15zdnd11an1n64x5 FILLER_288_8 ();
 b15zdnd11an1n64x5 FILLER_288_72 ();
 b15zdnd11an1n64x5 FILLER_288_136 ();
 b15zdnd11an1n64x5 FILLER_288_200 ();
 b15zdnd11an1n64x5 FILLER_288_264 ();
 b15zdnd11an1n64x5 FILLER_288_328 ();
 b15zdnd11an1n64x5 FILLER_288_392 ();
 b15zdnd11an1n64x5 FILLER_288_456 ();
 b15zdnd11an1n64x5 FILLER_288_520 ();
 b15zdnd11an1n64x5 FILLER_288_584 ();
 b15zdnd11an1n64x5 FILLER_288_648 ();
 b15zdnd11an1n04x5 FILLER_288_712 ();
 b15zdnd00an1n02x5 FILLER_288_716 ();
 b15zdnd11an1n64x5 FILLER_288_726 ();
 b15zdnd11an1n64x5 FILLER_288_790 ();
 b15zdnd11an1n64x5 FILLER_288_854 ();
 b15zdnd11an1n64x5 FILLER_288_918 ();
 b15zdnd11an1n64x5 FILLER_288_982 ();
 b15zdnd11an1n64x5 FILLER_288_1046 ();
 b15zdnd11an1n64x5 FILLER_288_1110 ();
 b15zdnd11an1n64x5 FILLER_288_1174 ();
 b15zdnd11an1n64x5 FILLER_288_1238 ();
 b15zdnd11an1n64x5 FILLER_288_1302 ();
 b15zdnd11an1n64x5 FILLER_288_1366 ();
 b15zdnd11an1n64x5 FILLER_288_1430 ();
 b15zdnd11an1n64x5 FILLER_288_1494 ();
 b15zdnd11an1n64x5 FILLER_288_1558 ();
 b15zdnd11an1n64x5 FILLER_288_1622 ();
 b15zdnd11an1n64x5 FILLER_288_1686 ();
 b15zdnd11an1n64x5 FILLER_288_1750 ();
 b15zdnd11an1n64x5 FILLER_288_1814 ();
 b15zdnd11an1n64x5 FILLER_288_1878 ();
 b15zdnd11an1n64x5 FILLER_288_1942 ();
 b15zdnd11an1n64x5 FILLER_288_2006 ();
 b15zdnd11an1n64x5 FILLER_288_2070 ();
 b15zdnd11an1n16x5 FILLER_288_2134 ();
 b15zdnd11an1n04x5 FILLER_288_2150 ();
 b15zdnd11an1n64x5 FILLER_288_2162 ();
 b15zdnd11an1n32x5 FILLER_288_2226 ();
 b15zdnd11an1n16x5 FILLER_288_2258 ();
 b15zdnd00an1n02x5 FILLER_288_2274 ();
 b15zdnd11an1n64x5 FILLER_289_0 ();
 b15zdnd11an1n64x5 FILLER_289_64 ();
 b15zdnd11an1n64x5 FILLER_289_128 ();
 b15zdnd11an1n64x5 FILLER_289_192 ();
 b15zdnd11an1n64x5 FILLER_289_256 ();
 b15zdnd11an1n64x5 FILLER_289_320 ();
 b15zdnd11an1n64x5 FILLER_289_384 ();
 b15zdnd11an1n64x5 FILLER_289_448 ();
 b15zdnd11an1n64x5 FILLER_289_512 ();
 b15zdnd11an1n64x5 FILLER_289_576 ();
 b15zdnd11an1n64x5 FILLER_289_640 ();
 b15zdnd11an1n64x5 FILLER_289_704 ();
 b15zdnd11an1n64x5 FILLER_289_768 ();
 b15zdnd11an1n64x5 FILLER_289_832 ();
 b15zdnd11an1n64x5 FILLER_289_896 ();
 b15zdnd11an1n64x5 FILLER_289_960 ();
 b15zdnd11an1n64x5 FILLER_289_1024 ();
 b15zdnd11an1n64x5 FILLER_289_1088 ();
 b15zdnd11an1n64x5 FILLER_289_1152 ();
 b15zdnd11an1n64x5 FILLER_289_1216 ();
 b15zdnd11an1n64x5 FILLER_289_1280 ();
 b15zdnd11an1n64x5 FILLER_289_1344 ();
 b15zdnd11an1n64x5 FILLER_289_1408 ();
 b15zdnd11an1n64x5 FILLER_289_1472 ();
 b15zdnd11an1n64x5 FILLER_289_1536 ();
 b15zdnd11an1n64x5 FILLER_289_1600 ();
 b15zdnd11an1n64x5 FILLER_289_1664 ();
 b15zdnd11an1n64x5 FILLER_289_1728 ();
 b15zdnd11an1n64x5 FILLER_289_1792 ();
 b15zdnd11an1n64x5 FILLER_289_1856 ();
 b15zdnd11an1n64x5 FILLER_289_1920 ();
 b15zdnd11an1n64x5 FILLER_289_1984 ();
 b15zdnd11an1n64x5 FILLER_289_2048 ();
 b15zdnd11an1n64x5 FILLER_289_2112 ();
 b15zdnd11an1n64x5 FILLER_289_2176 ();
 b15zdnd11an1n32x5 FILLER_289_2240 ();
 b15zdnd11an1n08x5 FILLER_289_2272 ();
 b15zdnd11an1n04x5 FILLER_289_2280 ();
 b15zdnd11an1n64x5 FILLER_290_8 ();
 b15zdnd11an1n64x5 FILLER_290_72 ();
 b15zdnd11an1n64x5 FILLER_290_136 ();
 b15zdnd11an1n64x5 FILLER_290_200 ();
 b15zdnd11an1n64x5 FILLER_290_264 ();
 b15zdnd11an1n64x5 FILLER_290_328 ();
 b15zdnd11an1n64x5 FILLER_290_392 ();
 b15zdnd11an1n64x5 FILLER_290_456 ();
 b15zdnd11an1n64x5 FILLER_290_520 ();
 b15zdnd11an1n64x5 FILLER_290_584 ();
 b15zdnd11an1n64x5 FILLER_290_648 ();
 b15zdnd11an1n04x5 FILLER_290_712 ();
 b15zdnd00an1n02x5 FILLER_290_716 ();
 b15zdnd11an1n64x5 FILLER_290_726 ();
 b15zdnd11an1n64x5 FILLER_290_790 ();
 b15zdnd11an1n64x5 FILLER_290_854 ();
 b15zdnd11an1n64x5 FILLER_290_918 ();
 b15zdnd11an1n64x5 FILLER_290_982 ();
 b15zdnd11an1n64x5 FILLER_290_1046 ();
 b15zdnd11an1n64x5 FILLER_290_1110 ();
 b15zdnd11an1n64x5 FILLER_290_1174 ();
 b15zdnd11an1n64x5 FILLER_290_1238 ();
 b15zdnd11an1n64x5 FILLER_290_1302 ();
 b15zdnd11an1n64x5 FILLER_290_1366 ();
 b15zdnd11an1n64x5 FILLER_290_1430 ();
 b15zdnd11an1n64x5 FILLER_290_1494 ();
 b15zdnd11an1n64x5 FILLER_290_1558 ();
 b15zdnd11an1n64x5 FILLER_290_1622 ();
 b15zdnd11an1n64x5 FILLER_290_1686 ();
 b15zdnd11an1n64x5 FILLER_290_1750 ();
 b15zdnd11an1n64x5 FILLER_290_1814 ();
 b15zdnd11an1n64x5 FILLER_290_1878 ();
 b15zdnd11an1n64x5 FILLER_290_1942 ();
 b15zdnd11an1n64x5 FILLER_290_2006 ();
 b15zdnd11an1n64x5 FILLER_290_2070 ();
 b15zdnd11an1n16x5 FILLER_290_2134 ();
 b15zdnd11an1n04x5 FILLER_290_2150 ();
 b15zdnd11an1n64x5 FILLER_290_2162 ();
 b15zdnd11an1n32x5 FILLER_290_2226 ();
 b15zdnd11an1n16x5 FILLER_290_2258 ();
 b15zdnd00an1n02x5 FILLER_290_2274 ();
 b15zdnd11an1n64x5 FILLER_291_0 ();
 b15zdnd11an1n64x5 FILLER_291_64 ();
 b15zdnd11an1n64x5 FILLER_291_128 ();
 b15zdnd11an1n64x5 FILLER_291_192 ();
 b15zdnd11an1n64x5 FILLER_291_256 ();
 b15zdnd11an1n64x5 FILLER_291_320 ();
 b15zdnd11an1n64x5 FILLER_291_384 ();
 b15zdnd11an1n64x5 FILLER_291_448 ();
 b15zdnd11an1n64x5 FILLER_291_512 ();
 b15zdnd11an1n64x5 FILLER_291_576 ();
 b15zdnd11an1n64x5 FILLER_291_640 ();
 b15zdnd11an1n64x5 FILLER_291_704 ();
 b15zdnd11an1n64x5 FILLER_291_768 ();
 b15zdnd11an1n64x5 FILLER_291_832 ();
 b15zdnd11an1n64x5 FILLER_291_896 ();
 b15zdnd11an1n64x5 FILLER_291_960 ();
 b15zdnd11an1n64x5 FILLER_291_1024 ();
 b15zdnd11an1n64x5 FILLER_291_1088 ();
 b15zdnd11an1n64x5 FILLER_291_1152 ();
 b15zdnd11an1n64x5 FILLER_291_1216 ();
 b15zdnd11an1n64x5 FILLER_291_1280 ();
 b15zdnd11an1n64x5 FILLER_291_1344 ();
 b15zdnd11an1n64x5 FILLER_291_1408 ();
 b15zdnd11an1n64x5 FILLER_291_1472 ();
 b15zdnd11an1n64x5 FILLER_291_1536 ();
 b15zdnd11an1n64x5 FILLER_291_1600 ();
 b15zdnd11an1n64x5 FILLER_291_1664 ();
 b15zdnd11an1n64x5 FILLER_291_1728 ();
 b15zdnd11an1n64x5 FILLER_291_1792 ();
 b15zdnd11an1n64x5 FILLER_291_1856 ();
 b15zdnd11an1n64x5 FILLER_291_1920 ();
 b15zdnd11an1n64x5 FILLER_291_1984 ();
 b15zdnd11an1n64x5 FILLER_291_2048 ();
 b15zdnd11an1n64x5 FILLER_291_2112 ();
 b15zdnd11an1n64x5 FILLER_291_2176 ();
 b15zdnd11an1n32x5 FILLER_291_2240 ();
 b15zdnd11an1n08x5 FILLER_291_2272 ();
 b15zdnd11an1n04x5 FILLER_291_2280 ();
 b15zdnd11an1n64x5 FILLER_292_8 ();
 b15zdnd11an1n64x5 FILLER_292_72 ();
 b15zdnd11an1n64x5 FILLER_292_136 ();
 b15zdnd11an1n64x5 FILLER_292_200 ();
 b15zdnd11an1n64x5 FILLER_292_264 ();
 b15zdnd11an1n64x5 FILLER_292_328 ();
 b15zdnd11an1n64x5 FILLER_292_392 ();
 b15zdnd11an1n64x5 FILLER_292_456 ();
 b15zdnd11an1n64x5 FILLER_292_520 ();
 b15zdnd11an1n64x5 FILLER_292_584 ();
 b15zdnd11an1n64x5 FILLER_292_648 ();
 b15zdnd11an1n04x5 FILLER_292_712 ();
 b15zdnd00an1n02x5 FILLER_292_716 ();
 b15zdnd11an1n64x5 FILLER_292_726 ();
 b15zdnd11an1n64x5 FILLER_292_790 ();
 b15zdnd11an1n64x5 FILLER_292_854 ();
 b15zdnd11an1n64x5 FILLER_292_918 ();
 b15zdnd11an1n64x5 FILLER_292_982 ();
 b15zdnd11an1n64x5 FILLER_292_1046 ();
 b15zdnd11an1n64x5 FILLER_292_1110 ();
 b15zdnd11an1n64x5 FILLER_292_1174 ();
 b15zdnd11an1n64x5 FILLER_292_1238 ();
 b15zdnd11an1n64x5 FILLER_292_1302 ();
 b15zdnd11an1n64x5 FILLER_292_1366 ();
 b15zdnd11an1n64x5 FILLER_292_1430 ();
 b15zdnd11an1n64x5 FILLER_292_1494 ();
 b15zdnd11an1n64x5 FILLER_292_1558 ();
 b15zdnd11an1n64x5 FILLER_292_1622 ();
 b15zdnd11an1n64x5 FILLER_292_1686 ();
 b15zdnd11an1n64x5 FILLER_292_1750 ();
 b15zdnd11an1n64x5 FILLER_292_1814 ();
 b15zdnd11an1n64x5 FILLER_292_1878 ();
 b15zdnd11an1n64x5 FILLER_292_1942 ();
 b15zdnd11an1n64x5 FILLER_292_2006 ();
 b15zdnd11an1n64x5 FILLER_292_2070 ();
 b15zdnd11an1n16x5 FILLER_292_2134 ();
 b15zdnd11an1n04x5 FILLER_292_2150 ();
 b15zdnd11an1n64x5 FILLER_292_2162 ();
 b15zdnd11an1n32x5 FILLER_292_2226 ();
 b15zdnd11an1n16x5 FILLER_292_2258 ();
 b15zdnd00an1n02x5 FILLER_292_2274 ();
 b15zdnd11an1n64x5 FILLER_293_0 ();
 b15zdnd11an1n64x5 FILLER_293_64 ();
 b15zdnd11an1n64x5 FILLER_293_128 ();
 b15zdnd11an1n64x5 FILLER_293_192 ();
 b15zdnd11an1n64x5 FILLER_293_256 ();
 b15zdnd11an1n64x5 FILLER_293_320 ();
 b15zdnd11an1n64x5 FILLER_293_384 ();
 b15zdnd11an1n64x5 FILLER_293_448 ();
 b15zdnd11an1n64x5 FILLER_293_512 ();
 b15zdnd11an1n64x5 FILLER_293_576 ();
 b15zdnd11an1n64x5 FILLER_293_640 ();
 b15zdnd11an1n64x5 FILLER_293_704 ();
 b15zdnd11an1n64x5 FILLER_293_768 ();
 b15zdnd11an1n64x5 FILLER_293_832 ();
 b15zdnd11an1n64x5 FILLER_293_896 ();
 b15zdnd11an1n64x5 FILLER_293_960 ();
 b15zdnd11an1n64x5 FILLER_293_1024 ();
 b15zdnd11an1n64x5 FILLER_293_1088 ();
 b15zdnd11an1n64x5 FILLER_293_1152 ();
 b15zdnd11an1n64x5 FILLER_293_1216 ();
 b15zdnd11an1n64x5 FILLER_293_1280 ();
 b15zdnd11an1n64x5 FILLER_293_1344 ();
 b15zdnd11an1n64x5 FILLER_293_1408 ();
 b15zdnd11an1n64x5 FILLER_293_1472 ();
 b15zdnd11an1n64x5 FILLER_293_1536 ();
 b15zdnd11an1n64x5 FILLER_293_1600 ();
 b15zdnd11an1n64x5 FILLER_293_1664 ();
 b15zdnd11an1n64x5 FILLER_293_1728 ();
 b15zdnd11an1n64x5 FILLER_293_1792 ();
 b15zdnd11an1n64x5 FILLER_293_1856 ();
 b15zdnd11an1n64x5 FILLER_293_1920 ();
 b15zdnd11an1n64x5 FILLER_293_1984 ();
 b15zdnd11an1n64x5 FILLER_293_2048 ();
 b15zdnd11an1n64x5 FILLER_293_2112 ();
 b15zdnd11an1n64x5 FILLER_293_2176 ();
 b15zdnd11an1n32x5 FILLER_293_2240 ();
 b15zdnd11an1n08x5 FILLER_293_2272 ();
 b15zdnd11an1n04x5 FILLER_293_2280 ();
 b15zdnd11an1n64x5 FILLER_294_8 ();
 b15zdnd11an1n64x5 FILLER_294_72 ();
 b15zdnd11an1n64x5 FILLER_294_136 ();
 b15zdnd11an1n64x5 FILLER_294_200 ();
 b15zdnd11an1n64x5 FILLER_294_264 ();
 b15zdnd11an1n64x5 FILLER_294_328 ();
 b15zdnd11an1n64x5 FILLER_294_392 ();
 b15zdnd11an1n64x5 FILLER_294_456 ();
 b15zdnd11an1n64x5 FILLER_294_520 ();
 b15zdnd11an1n64x5 FILLER_294_584 ();
 b15zdnd11an1n64x5 FILLER_294_648 ();
 b15zdnd11an1n04x5 FILLER_294_712 ();
 b15zdnd00an1n02x5 FILLER_294_716 ();
 b15zdnd11an1n64x5 FILLER_294_726 ();
 b15zdnd11an1n64x5 FILLER_294_790 ();
 b15zdnd11an1n64x5 FILLER_294_854 ();
 b15zdnd11an1n64x5 FILLER_294_918 ();
 b15zdnd11an1n64x5 FILLER_294_982 ();
 b15zdnd11an1n64x5 FILLER_294_1046 ();
 b15zdnd11an1n64x5 FILLER_294_1110 ();
 b15zdnd11an1n64x5 FILLER_294_1174 ();
 b15zdnd11an1n64x5 FILLER_294_1238 ();
 b15zdnd11an1n64x5 FILLER_294_1302 ();
 b15zdnd11an1n64x5 FILLER_294_1366 ();
 b15zdnd11an1n64x5 FILLER_294_1430 ();
 b15zdnd11an1n64x5 FILLER_294_1494 ();
 b15zdnd11an1n64x5 FILLER_294_1558 ();
 b15zdnd11an1n64x5 FILLER_294_1622 ();
 b15zdnd11an1n64x5 FILLER_294_1686 ();
 b15zdnd11an1n64x5 FILLER_294_1750 ();
 b15zdnd11an1n64x5 FILLER_294_1814 ();
 b15zdnd11an1n64x5 FILLER_294_1878 ();
 b15zdnd11an1n64x5 FILLER_294_1942 ();
 b15zdnd11an1n64x5 FILLER_294_2006 ();
 b15zdnd11an1n64x5 FILLER_294_2070 ();
 b15zdnd11an1n16x5 FILLER_294_2134 ();
 b15zdnd11an1n04x5 FILLER_294_2150 ();
 b15zdnd11an1n64x5 FILLER_294_2162 ();
 b15zdnd11an1n32x5 FILLER_294_2226 ();
 b15zdnd11an1n16x5 FILLER_294_2258 ();
 b15zdnd00an1n02x5 FILLER_294_2274 ();
 b15zdnd11an1n64x5 FILLER_295_0 ();
 b15zdnd11an1n64x5 FILLER_295_64 ();
 b15zdnd11an1n64x5 FILLER_295_128 ();
 b15zdnd11an1n64x5 FILLER_295_192 ();
 b15zdnd11an1n64x5 FILLER_295_256 ();
 b15zdnd11an1n64x5 FILLER_295_320 ();
 b15zdnd11an1n64x5 FILLER_295_384 ();
 b15zdnd11an1n64x5 FILLER_295_448 ();
 b15zdnd11an1n64x5 FILLER_295_512 ();
 b15zdnd11an1n64x5 FILLER_295_576 ();
 b15zdnd11an1n64x5 FILLER_295_640 ();
 b15zdnd11an1n64x5 FILLER_295_704 ();
 b15zdnd11an1n64x5 FILLER_295_768 ();
 b15zdnd11an1n64x5 FILLER_295_832 ();
 b15zdnd11an1n64x5 FILLER_295_896 ();
 b15zdnd11an1n64x5 FILLER_295_960 ();
 b15zdnd11an1n64x5 FILLER_295_1024 ();
 b15zdnd11an1n64x5 FILLER_295_1088 ();
 b15zdnd11an1n64x5 FILLER_295_1152 ();
 b15zdnd11an1n64x5 FILLER_295_1216 ();
 b15zdnd11an1n64x5 FILLER_295_1280 ();
 b15zdnd11an1n64x5 FILLER_295_1344 ();
 b15zdnd11an1n64x5 FILLER_295_1408 ();
 b15zdnd11an1n64x5 FILLER_295_1472 ();
 b15zdnd11an1n64x5 FILLER_295_1536 ();
 b15zdnd11an1n64x5 FILLER_295_1600 ();
 b15zdnd11an1n64x5 FILLER_295_1664 ();
 b15zdnd11an1n64x5 FILLER_295_1728 ();
 b15zdnd11an1n64x5 FILLER_295_1792 ();
 b15zdnd11an1n64x5 FILLER_295_1856 ();
 b15zdnd11an1n64x5 FILLER_295_1920 ();
 b15zdnd11an1n64x5 FILLER_295_1984 ();
 b15zdnd11an1n64x5 FILLER_295_2048 ();
 b15zdnd11an1n64x5 FILLER_295_2112 ();
 b15zdnd11an1n64x5 FILLER_295_2176 ();
 b15zdnd11an1n32x5 FILLER_295_2240 ();
 b15zdnd11an1n08x5 FILLER_295_2272 ();
 b15zdnd11an1n04x5 FILLER_295_2280 ();
 b15zdnd11an1n64x5 FILLER_296_8 ();
 b15zdnd11an1n64x5 FILLER_296_72 ();
 b15zdnd11an1n64x5 FILLER_296_136 ();
 b15zdnd11an1n64x5 FILLER_296_200 ();
 b15zdnd11an1n64x5 FILLER_296_264 ();
 b15zdnd11an1n64x5 FILLER_296_328 ();
 b15zdnd11an1n64x5 FILLER_296_392 ();
 b15zdnd11an1n64x5 FILLER_296_456 ();
 b15zdnd11an1n64x5 FILLER_296_520 ();
 b15zdnd11an1n64x5 FILLER_296_584 ();
 b15zdnd11an1n64x5 FILLER_296_648 ();
 b15zdnd11an1n04x5 FILLER_296_712 ();
 b15zdnd00an1n02x5 FILLER_296_716 ();
 b15zdnd11an1n64x5 FILLER_296_726 ();
 b15zdnd11an1n64x5 FILLER_296_790 ();
 b15zdnd11an1n64x5 FILLER_296_854 ();
 b15zdnd11an1n64x5 FILLER_296_918 ();
 b15zdnd11an1n64x5 FILLER_296_982 ();
 b15zdnd11an1n64x5 FILLER_296_1046 ();
 b15zdnd11an1n64x5 FILLER_296_1110 ();
 b15zdnd11an1n64x5 FILLER_296_1174 ();
 b15zdnd11an1n64x5 FILLER_296_1238 ();
 b15zdnd11an1n64x5 FILLER_296_1302 ();
 b15zdnd11an1n64x5 FILLER_296_1366 ();
 b15zdnd11an1n64x5 FILLER_296_1430 ();
 b15zdnd11an1n64x5 FILLER_296_1494 ();
 b15zdnd11an1n64x5 FILLER_296_1558 ();
 b15zdnd11an1n64x5 FILLER_296_1622 ();
 b15zdnd11an1n64x5 FILLER_296_1686 ();
 b15zdnd11an1n64x5 FILLER_296_1750 ();
 b15zdnd11an1n64x5 FILLER_296_1814 ();
 b15zdnd11an1n64x5 FILLER_296_1878 ();
 b15zdnd11an1n64x5 FILLER_296_1942 ();
 b15zdnd11an1n64x5 FILLER_296_2006 ();
 b15zdnd11an1n64x5 FILLER_296_2070 ();
 b15zdnd11an1n16x5 FILLER_296_2134 ();
 b15zdnd11an1n04x5 FILLER_296_2150 ();
 b15zdnd11an1n64x5 FILLER_296_2162 ();
 b15zdnd11an1n32x5 FILLER_296_2226 ();
 b15zdnd11an1n16x5 FILLER_296_2258 ();
 b15zdnd00an1n02x5 FILLER_296_2274 ();
 b15zdnd11an1n64x5 FILLER_297_0 ();
 b15zdnd11an1n64x5 FILLER_297_64 ();
 b15zdnd11an1n64x5 FILLER_297_128 ();
 b15zdnd11an1n64x5 FILLER_297_192 ();
 b15zdnd11an1n64x5 FILLER_297_256 ();
 b15zdnd11an1n64x5 FILLER_297_320 ();
 b15zdnd11an1n64x5 FILLER_297_384 ();
 b15zdnd11an1n64x5 FILLER_297_448 ();
 b15zdnd11an1n64x5 FILLER_297_512 ();
 b15zdnd11an1n64x5 FILLER_297_576 ();
 b15zdnd11an1n64x5 FILLER_297_640 ();
 b15zdnd11an1n64x5 FILLER_297_704 ();
 b15zdnd11an1n64x5 FILLER_297_768 ();
 b15zdnd11an1n64x5 FILLER_297_832 ();
 b15zdnd11an1n64x5 FILLER_297_896 ();
 b15zdnd11an1n64x5 FILLER_297_960 ();
 b15zdnd11an1n64x5 FILLER_297_1024 ();
 b15zdnd11an1n64x5 FILLER_297_1088 ();
 b15zdnd11an1n64x5 FILLER_297_1152 ();
 b15zdnd11an1n64x5 FILLER_297_1216 ();
 b15zdnd11an1n64x5 FILLER_297_1280 ();
 b15zdnd11an1n64x5 FILLER_297_1344 ();
 b15zdnd11an1n64x5 FILLER_297_1408 ();
 b15zdnd11an1n64x5 FILLER_297_1472 ();
 b15zdnd11an1n64x5 FILLER_297_1536 ();
 b15zdnd11an1n64x5 FILLER_297_1600 ();
 b15zdnd11an1n64x5 FILLER_297_1664 ();
 b15zdnd11an1n64x5 FILLER_297_1728 ();
 b15zdnd11an1n64x5 FILLER_297_1792 ();
 b15zdnd11an1n64x5 FILLER_297_1856 ();
 b15zdnd11an1n64x5 FILLER_297_1920 ();
 b15zdnd11an1n64x5 FILLER_297_1984 ();
 b15zdnd11an1n64x5 FILLER_297_2048 ();
 b15zdnd11an1n64x5 FILLER_297_2112 ();
 b15zdnd11an1n64x5 FILLER_297_2176 ();
 b15zdnd11an1n32x5 FILLER_297_2240 ();
 b15zdnd11an1n08x5 FILLER_297_2272 ();
 b15zdnd11an1n04x5 FILLER_297_2280 ();
 b15zdnd11an1n64x5 FILLER_298_8 ();
 b15zdnd11an1n64x5 FILLER_298_72 ();
 b15zdnd11an1n64x5 FILLER_298_136 ();
 b15zdnd11an1n64x5 FILLER_298_200 ();
 b15zdnd11an1n64x5 FILLER_298_264 ();
 b15zdnd11an1n64x5 FILLER_298_328 ();
 b15zdnd11an1n64x5 FILLER_298_392 ();
 b15zdnd11an1n64x5 FILLER_298_456 ();
 b15zdnd11an1n64x5 FILLER_298_520 ();
 b15zdnd11an1n64x5 FILLER_298_584 ();
 b15zdnd11an1n64x5 FILLER_298_648 ();
 b15zdnd11an1n04x5 FILLER_298_712 ();
 b15zdnd00an1n02x5 FILLER_298_716 ();
 b15zdnd11an1n64x5 FILLER_298_726 ();
 b15zdnd11an1n64x5 FILLER_298_790 ();
 b15zdnd11an1n64x5 FILLER_298_854 ();
 b15zdnd11an1n64x5 FILLER_298_918 ();
 b15zdnd11an1n64x5 FILLER_298_982 ();
 b15zdnd11an1n64x5 FILLER_298_1046 ();
 b15zdnd11an1n64x5 FILLER_298_1110 ();
 b15zdnd11an1n64x5 FILLER_298_1174 ();
 b15zdnd11an1n64x5 FILLER_298_1238 ();
 b15zdnd11an1n64x5 FILLER_298_1302 ();
 b15zdnd11an1n64x5 FILLER_298_1366 ();
 b15zdnd11an1n64x5 FILLER_298_1430 ();
 b15zdnd11an1n64x5 FILLER_298_1494 ();
 b15zdnd11an1n64x5 FILLER_298_1558 ();
 b15zdnd11an1n64x5 FILLER_298_1622 ();
 b15zdnd11an1n64x5 FILLER_298_1686 ();
 b15zdnd11an1n64x5 FILLER_298_1750 ();
 b15zdnd11an1n64x5 FILLER_298_1814 ();
 b15zdnd11an1n64x5 FILLER_298_1878 ();
 b15zdnd11an1n64x5 FILLER_298_1942 ();
 b15zdnd11an1n64x5 FILLER_298_2006 ();
 b15zdnd11an1n64x5 FILLER_298_2070 ();
 b15zdnd11an1n16x5 FILLER_298_2134 ();
 b15zdnd11an1n04x5 FILLER_298_2150 ();
 b15zdnd11an1n64x5 FILLER_298_2162 ();
 b15zdnd11an1n32x5 FILLER_298_2226 ();
 b15zdnd11an1n16x5 FILLER_298_2258 ();
 b15zdnd00an1n02x5 FILLER_298_2274 ();
 b15zdnd11an1n64x5 FILLER_299_0 ();
 b15zdnd11an1n64x5 FILLER_299_64 ();
 b15zdnd11an1n64x5 FILLER_299_128 ();
 b15zdnd11an1n64x5 FILLER_299_192 ();
 b15zdnd11an1n64x5 FILLER_299_256 ();
 b15zdnd11an1n64x5 FILLER_299_320 ();
 b15zdnd11an1n64x5 FILLER_299_384 ();
 b15zdnd11an1n64x5 FILLER_299_448 ();
 b15zdnd11an1n64x5 FILLER_299_512 ();
 b15zdnd11an1n64x5 FILLER_299_576 ();
 b15zdnd11an1n64x5 FILLER_299_640 ();
 b15zdnd11an1n64x5 FILLER_299_704 ();
 b15zdnd11an1n64x5 FILLER_299_768 ();
 b15zdnd11an1n64x5 FILLER_299_832 ();
 b15zdnd11an1n64x5 FILLER_299_896 ();
 b15zdnd11an1n64x5 FILLER_299_960 ();
 b15zdnd11an1n64x5 FILLER_299_1024 ();
 b15zdnd11an1n64x5 FILLER_299_1088 ();
 b15zdnd11an1n64x5 FILLER_299_1152 ();
 b15zdnd11an1n64x5 FILLER_299_1216 ();
 b15zdnd11an1n64x5 FILLER_299_1280 ();
 b15zdnd11an1n64x5 FILLER_299_1344 ();
 b15zdnd11an1n64x5 FILLER_299_1408 ();
 b15zdnd11an1n64x5 FILLER_299_1472 ();
 b15zdnd11an1n64x5 FILLER_299_1536 ();
 b15zdnd11an1n64x5 FILLER_299_1600 ();
 b15zdnd11an1n64x5 FILLER_299_1664 ();
 b15zdnd11an1n64x5 FILLER_299_1728 ();
 b15zdnd11an1n64x5 FILLER_299_1792 ();
 b15zdnd11an1n64x5 FILLER_299_1856 ();
 b15zdnd11an1n64x5 FILLER_299_1920 ();
 b15zdnd11an1n64x5 FILLER_299_1984 ();
 b15zdnd11an1n64x5 FILLER_299_2048 ();
 b15zdnd11an1n64x5 FILLER_299_2112 ();
 b15zdnd11an1n64x5 FILLER_299_2176 ();
 b15zdnd11an1n32x5 FILLER_299_2240 ();
 b15zdnd11an1n08x5 FILLER_299_2272 ();
 b15zdnd11an1n04x5 FILLER_299_2280 ();
 b15zdnd11an1n64x5 FILLER_300_8 ();
 b15zdnd11an1n64x5 FILLER_300_72 ();
 b15zdnd11an1n64x5 FILLER_300_136 ();
 b15zdnd11an1n64x5 FILLER_300_200 ();
 b15zdnd11an1n64x5 FILLER_300_264 ();
 b15zdnd11an1n64x5 FILLER_300_328 ();
 b15zdnd11an1n64x5 FILLER_300_392 ();
 b15zdnd11an1n64x5 FILLER_300_456 ();
 b15zdnd11an1n64x5 FILLER_300_520 ();
 b15zdnd11an1n64x5 FILLER_300_584 ();
 b15zdnd11an1n64x5 FILLER_300_648 ();
 b15zdnd11an1n04x5 FILLER_300_712 ();
 b15zdnd00an1n02x5 FILLER_300_716 ();
 b15zdnd11an1n64x5 FILLER_300_726 ();
 b15zdnd11an1n64x5 FILLER_300_790 ();
 b15zdnd11an1n64x5 FILLER_300_854 ();
 b15zdnd11an1n64x5 FILLER_300_918 ();
 b15zdnd11an1n64x5 FILLER_300_982 ();
 b15zdnd11an1n64x5 FILLER_300_1046 ();
 b15zdnd11an1n64x5 FILLER_300_1110 ();
 b15zdnd11an1n64x5 FILLER_300_1174 ();
 b15zdnd11an1n64x5 FILLER_300_1238 ();
 b15zdnd11an1n64x5 FILLER_300_1302 ();
 b15zdnd11an1n64x5 FILLER_300_1366 ();
 b15zdnd11an1n64x5 FILLER_300_1430 ();
 b15zdnd11an1n64x5 FILLER_300_1494 ();
 b15zdnd11an1n64x5 FILLER_300_1558 ();
 b15zdnd11an1n64x5 FILLER_300_1622 ();
 b15zdnd11an1n64x5 FILLER_300_1686 ();
 b15zdnd11an1n64x5 FILLER_300_1750 ();
 b15zdnd11an1n64x5 FILLER_300_1814 ();
 b15zdnd11an1n64x5 FILLER_300_1878 ();
 b15zdnd11an1n64x5 FILLER_300_1942 ();
 b15zdnd11an1n64x5 FILLER_300_2006 ();
 b15zdnd11an1n64x5 FILLER_300_2070 ();
 b15zdnd11an1n16x5 FILLER_300_2134 ();
 b15zdnd11an1n04x5 FILLER_300_2150 ();
 b15zdnd11an1n64x5 FILLER_300_2162 ();
 b15zdnd11an1n32x5 FILLER_300_2226 ();
 b15zdnd11an1n16x5 FILLER_300_2258 ();
 b15zdnd00an1n02x5 FILLER_300_2274 ();
 b15zdnd11an1n64x5 FILLER_301_0 ();
 b15zdnd11an1n64x5 FILLER_301_64 ();
 b15zdnd11an1n64x5 FILLER_301_128 ();
 b15zdnd11an1n64x5 FILLER_301_192 ();
 b15zdnd11an1n64x5 FILLER_301_256 ();
 b15zdnd11an1n64x5 FILLER_301_320 ();
 b15zdnd11an1n64x5 FILLER_301_384 ();
 b15zdnd11an1n64x5 FILLER_301_448 ();
 b15zdnd11an1n64x5 FILLER_301_512 ();
 b15zdnd11an1n64x5 FILLER_301_576 ();
 b15zdnd11an1n64x5 FILLER_301_640 ();
 b15zdnd11an1n64x5 FILLER_301_704 ();
 b15zdnd11an1n64x5 FILLER_301_768 ();
 b15zdnd11an1n64x5 FILLER_301_832 ();
 b15zdnd11an1n64x5 FILLER_301_896 ();
 b15zdnd11an1n64x5 FILLER_301_960 ();
 b15zdnd11an1n64x5 FILLER_301_1024 ();
 b15zdnd11an1n64x5 FILLER_301_1088 ();
 b15zdnd11an1n64x5 FILLER_301_1152 ();
 b15zdnd11an1n64x5 FILLER_301_1216 ();
 b15zdnd11an1n64x5 FILLER_301_1280 ();
 b15zdnd11an1n64x5 FILLER_301_1344 ();
 b15zdnd11an1n64x5 FILLER_301_1408 ();
 b15zdnd11an1n64x5 FILLER_301_1472 ();
 b15zdnd11an1n64x5 FILLER_301_1536 ();
 b15zdnd11an1n64x5 FILLER_301_1600 ();
 b15zdnd11an1n64x5 FILLER_301_1664 ();
 b15zdnd11an1n64x5 FILLER_301_1728 ();
 b15zdnd11an1n64x5 FILLER_301_1792 ();
 b15zdnd11an1n64x5 FILLER_301_1856 ();
 b15zdnd11an1n64x5 FILLER_301_1920 ();
 b15zdnd11an1n64x5 FILLER_301_1984 ();
 b15zdnd11an1n64x5 FILLER_301_2048 ();
 b15zdnd11an1n64x5 FILLER_301_2112 ();
 b15zdnd11an1n64x5 FILLER_301_2176 ();
 b15zdnd11an1n32x5 FILLER_301_2240 ();
 b15zdnd11an1n08x5 FILLER_301_2272 ();
 b15zdnd11an1n04x5 FILLER_301_2280 ();
 b15zdnd11an1n64x5 FILLER_302_8 ();
 b15zdnd11an1n64x5 FILLER_302_72 ();
 b15zdnd11an1n64x5 FILLER_302_136 ();
 b15zdnd11an1n64x5 FILLER_302_200 ();
 b15zdnd11an1n64x5 FILLER_302_264 ();
 b15zdnd11an1n64x5 FILLER_302_328 ();
 b15zdnd11an1n64x5 FILLER_302_392 ();
 b15zdnd11an1n64x5 FILLER_302_456 ();
 b15zdnd11an1n64x5 FILLER_302_520 ();
 b15zdnd11an1n64x5 FILLER_302_584 ();
 b15zdnd11an1n64x5 FILLER_302_648 ();
 b15zdnd11an1n04x5 FILLER_302_712 ();
 b15zdnd00an1n02x5 FILLER_302_716 ();
 b15zdnd11an1n64x5 FILLER_302_726 ();
 b15zdnd11an1n64x5 FILLER_302_790 ();
 b15zdnd11an1n64x5 FILLER_302_854 ();
 b15zdnd11an1n64x5 FILLER_302_918 ();
 b15zdnd11an1n64x5 FILLER_302_982 ();
 b15zdnd11an1n64x5 FILLER_302_1046 ();
 b15zdnd11an1n64x5 FILLER_302_1110 ();
 b15zdnd11an1n64x5 FILLER_302_1174 ();
 b15zdnd11an1n64x5 FILLER_302_1238 ();
 b15zdnd11an1n64x5 FILLER_302_1302 ();
 b15zdnd11an1n64x5 FILLER_302_1366 ();
 b15zdnd11an1n64x5 FILLER_302_1430 ();
 b15zdnd11an1n64x5 FILLER_302_1494 ();
 b15zdnd11an1n64x5 FILLER_302_1558 ();
 b15zdnd11an1n64x5 FILLER_302_1622 ();
 b15zdnd11an1n64x5 FILLER_302_1686 ();
 b15zdnd11an1n64x5 FILLER_302_1750 ();
 b15zdnd11an1n64x5 FILLER_302_1814 ();
 b15zdnd11an1n64x5 FILLER_302_1878 ();
 b15zdnd11an1n64x5 FILLER_302_1942 ();
 b15zdnd11an1n64x5 FILLER_302_2006 ();
 b15zdnd11an1n64x5 FILLER_302_2070 ();
 b15zdnd11an1n16x5 FILLER_302_2134 ();
 b15zdnd11an1n04x5 FILLER_302_2150 ();
 b15zdnd11an1n64x5 FILLER_302_2162 ();
 b15zdnd11an1n32x5 FILLER_302_2226 ();
 b15zdnd11an1n16x5 FILLER_302_2258 ();
 b15zdnd00an1n02x5 FILLER_302_2274 ();
 b15zdnd11an1n64x5 FILLER_303_0 ();
 b15zdnd11an1n64x5 FILLER_303_64 ();
 b15zdnd11an1n64x5 FILLER_303_128 ();
 b15zdnd11an1n64x5 FILLER_303_192 ();
 b15zdnd11an1n64x5 FILLER_303_256 ();
 b15zdnd11an1n64x5 FILLER_303_320 ();
 b15zdnd11an1n64x5 FILLER_303_384 ();
 b15zdnd11an1n64x5 FILLER_303_448 ();
 b15zdnd11an1n64x5 FILLER_303_512 ();
 b15zdnd11an1n64x5 FILLER_303_576 ();
 b15zdnd11an1n64x5 FILLER_303_640 ();
 b15zdnd11an1n64x5 FILLER_303_704 ();
 b15zdnd11an1n64x5 FILLER_303_768 ();
 b15zdnd11an1n64x5 FILLER_303_832 ();
 b15zdnd11an1n64x5 FILLER_303_896 ();
 b15zdnd11an1n64x5 FILLER_303_960 ();
 b15zdnd11an1n64x5 FILLER_303_1024 ();
 b15zdnd11an1n64x5 FILLER_303_1088 ();
 b15zdnd11an1n64x5 FILLER_303_1152 ();
 b15zdnd11an1n64x5 FILLER_303_1216 ();
 b15zdnd11an1n64x5 FILLER_303_1280 ();
 b15zdnd11an1n64x5 FILLER_303_1344 ();
 b15zdnd11an1n64x5 FILLER_303_1408 ();
 b15zdnd11an1n64x5 FILLER_303_1472 ();
 b15zdnd11an1n64x5 FILLER_303_1536 ();
 b15zdnd11an1n64x5 FILLER_303_1600 ();
 b15zdnd11an1n64x5 FILLER_303_1664 ();
 b15zdnd11an1n64x5 FILLER_303_1728 ();
 b15zdnd11an1n64x5 FILLER_303_1792 ();
 b15zdnd11an1n64x5 FILLER_303_1856 ();
 b15zdnd11an1n64x5 FILLER_303_1920 ();
 b15zdnd11an1n64x5 FILLER_303_1984 ();
 b15zdnd11an1n64x5 FILLER_303_2048 ();
 b15zdnd11an1n64x5 FILLER_303_2112 ();
 b15zdnd11an1n64x5 FILLER_303_2176 ();
 b15zdnd11an1n32x5 FILLER_303_2240 ();
 b15zdnd11an1n08x5 FILLER_303_2272 ();
 b15zdnd11an1n04x5 FILLER_303_2280 ();
 b15zdnd11an1n64x5 FILLER_304_8 ();
 b15zdnd11an1n64x5 FILLER_304_72 ();
 b15zdnd11an1n64x5 FILLER_304_136 ();
 b15zdnd11an1n64x5 FILLER_304_200 ();
 b15zdnd11an1n64x5 FILLER_304_264 ();
 b15zdnd11an1n64x5 FILLER_304_328 ();
 b15zdnd11an1n64x5 FILLER_304_392 ();
 b15zdnd11an1n64x5 FILLER_304_456 ();
 b15zdnd11an1n64x5 FILLER_304_520 ();
 b15zdnd11an1n64x5 FILLER_304_584 ();
 b15zdnd11an1n64x5 FILLER_304_648 ();
 b15zdnd11an1n04x5 FILLER_304_712 ();
 b15zdnd00an1n02x5 FILLER_304_716 ();
 b15zdnd11an1n64x5 FILLER_304_726 ();
 b15zdnd11an1n64x5 FILLER_304_790 ();
 b15zdnd11an1n64x5 FILLER_304_854 ();
 b15zdnd11an1n32x5 FILLER_304_918 ();
 b15zdnd11an1n16x5 FILLER_304_950 ();
 b15zdnd00an1n02x5 FILLER_304_966 ();
 b15zdnd11an1n64x5 FILLER_304_1010 ();
 b15zdnd11an1n64x5 FILLER_304_1074 ();
 b15zdnd11an1n64x5 FILLER_304_1138 ();
 b15zdnd11an1n64x5 FILLER_304_1202 ();
 b15zdnd11an1n64x5 FILLER_304_1266 ();
 b15zdnd11an1n64x5 FILLER_304_1330 ();
 b15zdnd11an1n64x5 FILLER_304_1394 ();
 b15zdnd11an1n64x5 FILLER_304_1458 ();
 b15zdnd11an1n64x5 FILLER_304_1522 ();
 b15zdnd11an1n64x5 FILLER_304_1586 ();
 b15zdnd11an1n64x5 FILLER_304_1650 ();
 b15zdnd11an1n64x5 FILLER_304_1714 ();
 b15zdnd11an1n64x5 FILLER_304_1778 ();
 b15zdnd11an1n64x5 FILLER_304_1842 ();
 b15zdnd11an1n64x5 FILLER_304_1906 ();
 b15zdnd11an1n64x5 FILLER_304_1970 ();
 b15zdnd11an1n64x5 FILLER_304_2034 ();
 b15zdnd11an1n32x5 FILLER_304_2098 ();
 b15zdnd11an1n16x5 FILLER_304_2130 ();
 b15zdnd11an1n08x5 FILLER_304_2146 ();
 b15zdnd11an1n64x5 FILLER_304_2162 ();
 b15zdnd11an1n32x5 FILLER_304_2226 ();
 b15zdnd11an1n16x5 FILLER_304_2258 ();
 b15zdnd00an1n02x5 FILLER_304_2274 ();
 b15zdnd11an1n64x5 FILLER_305_0 ();
 b15zdnd11an1n64x5 FILLER_305_64 ();
 b15zdnd11an1n64x5 FILLER_305_128 ();
 b15zdnd11an1n64x5 FILLER_305_192 ();
 b15zdnd11an1n64x5 FILLER_305_256 ();
 b15zdnd11an1n64x5 FILLER_305_320 ();
 b15zdnd11an1n64x5 FILLER_305_384 ();
 b15zdnd11an1n64x5 FILLER_305_448 ();
 b15zdnd11an1n64x5 FILLER_305_512 ();
 b15zdnd11an1n64x5 FILLER_305_576 ();
 b15zdnd11an1n64x5 FILLER_305_640 ();
 b15zdnd11an1n64x5 FILLER_305_704 ();
 b15zdnd11an1n64x5 FILLER_305_768 ();
 b15zdnd11an1n64x5 FILLER_305_832 ();
 b15zdnd11an1n64x5 FILLER_305_896 ();
 b15zdnd11an1n04x5 FILLER_305_960 ();
 b15zdnd11an1n64x5 FILLER_305_1006 ();
 b15zdnd11an1n64x5 FILLER_305_1070 ();
 b15zdnd11an1n64x5 FILLER_305_1134 ();
 b15zdnd11an1n64x5 FILLER_305_1198 ();
 b15zdnd11an1n64x5 FILLER_305_1262 ();
 b15zdnd11an1n64x5 FILLER_305_1326 ();
 b15zdnd11an1n64x5 FILLER_305_1390 ();
 b15zdnd11an1n64x5 FILLER_305_1454 ();
 b15zdnd11an1n64x5 FILLER_305_1518 ();
 b15zdnd11an1n64x5 FILLER_305_1582 ();
 b15zdnd11an1n64x5 FILLER_305_1646 ();
 b15zdnd11an1n64x5 FILLER_305_1710 ();
 b15zdnd11an1n64x5 FILLER_305_1774 ();
 b15zdnd11an1n64x5 FILLER_305_1838 ();
 b15zdnd11an1n64x5 FILLER_305_1902 ();
 b15zdnd11an1n64x5 FILLER_305_1966 ();
 b15zdnd11an1n64x5 FILLER_305_2030 ();
 b15zdnd11an1n64x5 FILLER_305_2094 ();
 b15zdnd11an1n64x5 FILLER_305_2158 ();
 b15zdnd11an1n32x5 FILLER_305_2222 ();
 b15zdnd11an1n16x5 FILLER_305_2254 ();
 b15zdnd11an1n08x5 FILLER_305_2270 ();
 b15zdnd11an1n04x5 FILLER_305_2278 ();
 b15zdnd00an1n02x5 FILLER_305_2282 ();
 b15zdnd11an1n64x5 FILLER_306_8 ();
 b15zdnd11an1n64x5 FILLER_306_72 ();
 b15zdnd11an1n64x5 FILLER_306_136 ();
 b15zdnd11an1n64x5 FILLER_306_200 ();
 b15zdnd11an1n64x5 FILLER_306_264 ();
 b15zdnd11an1n64x5 FILLER_306_328 ();
 b15zdnd11an1n64x5 FILLER_306_392 ();
 b15zdnd11an1n64x5 FILLER_306_456 ();
 b15zdnd11an1n64x5 FILLER_306_520 ();
 b15zdnd11an1n64x5 FILLER_306_584 ();
 b15zdnd11an1n64x5 FILLER_306_648 ();
 b15zdnd11an1n04x5 FILLER_306_712 ();
 b15zdnd00an1n02x5 FILLER_306_716 ();
 b15zdnd11an1n64x5 FILLER_306_726 ();
 b15zdnd11an1n32x5 FILLER_306_790 ();
 b15zdnd11an1n08x5 FILLER_306_822 ();
 b15zdnd00an1n02x5 FILLER_306_830 ();
 b15zdnd11an1n64x5 FILLER_306_874 ();
 b15zdnd11an1n32x5 FILLER_306_938 ();
 b15zdnd00an1n01x5 FILLER_306_970 ();
 b15zdnd11an1n64x5 FILLER_306_1013 ();
 b15zdnd11an1n64x5 FILLER_306_1077 ();
 b15zdnd11an1n64x5 FILLER_306_1141 ();
 b15zdnd11an1n64x5 FILLER_306_1205 ();
 b15zdnd11an1n64x5 FILLER_306_1269 ();
 b15zdnd11an1n64x5 FILLER_306_1333 ();
 b15zdnd11an1n64x5 FILLER_306_1397 ();
 b15zdnd11an1n64x5 FILLER_306_1461 ();
 b15zdnd11an1n64x5 FILLER_306_1525 ();
 b15zdnd11an1n64x5 FILLER_306_1589 ();
 b15zdnd11an1n64x5 FILLER_306_1653 ();
 b15zdnd11an1n64x5 FILLER_306_1717 ();
 b15zdnd11an1n64x5 FILLER_306_1781 ();
 b15zdnd11an1n64x5 FILLER_306_1845 ();
 b15zdnd11an1n64x5 FILLER_306_1909 ();
 b15zdnd11an1n64x5 FILLER_306_1973 ();
 b15zdnd11an1n64x5 FILLER_306_2037 ();
 b15zdnd11an1n32x5 FILLER_306_2101 ();
 b15zdnd11an1n16x5 FILLER_306_2133 ();
 b15zdnd11an1n04x5 FILLER_306_2149 ();
 b15zdnd00an1n01x5 FILLER_306_2153 ();
 b15zdnd11an1n64x5 FILLER_306_2162 ();
 b15zdnd11an1n32x5 FILLER_306_2226 ();
 b15zdnd11an1n16x5 FILLER_306_2258 ();
 b15zdnd00an1n02x5 FILLER_306_2274 ();
 b15zdnd11an1n64x5 FILLER_307_0 ();
 b15zdnd11an1n64x5 FILLER_307_64 ();
 b15zdnd11an1n64x5 FILLER_307_128 ();
 b15zdnd11an1n64x5 FILLER_307_192 ();
 b15zdnd11an1n64x5 FILLER_307_256 ();
 b15zdnd11an1n64x5 FILLER_307_320 ();
 b15zdnd11an1n64x5 FILLER_307_384 ();
 b15zdnd11an1n64x5 FILLER_307_448 ();
 b15zdnd11an1n64x5 FILLER_307_512 ();
 b15zdnd11an1n64x5 FILLER_307_576 ();
 b15zdnd11an1n64x5 FILLER_307_640 ();
 b15zdnd11an1n64x5 FILLER_307_704 ();
 b15zdnd11an1n64x5 FILLER_307_768 ();
 b15zdnd00an1n02x5 FILLER_307_832 ();
 b15zdnd11an1n64x5 FILLER_307_876 ();
 b15zdnd11an1n64x5 FILLER_307_940 ();
 b15zdnd11an1n64x5 FILLER_307_1004 ();
 b15zdnd11an1n64x5 FILLER_307_1068 ();
 b15zdnd11an1n64x5 FILLER_307_1132 ();
 b15zdnd11an1n64x5 FILLER_307_1196 ();
 b15zdnd11an1n64x5 FILLER_307_1260 ();
 b15zdnd11an1n64x5 FILLER_307_1324 ();
 b15zdnd11an1n64x5 FILLER_307_1388 ();
 b15zdnd11an1n64x5 FILLER_307_1452 ();
 b15zdnd11an1n64x5 FILLER_307_1516 ();
 b15zdnd11an1n64x5 FILLER_307_1580 ();
 b15zdnd11an1n64x5 FILLER_307_1644 ();
 b15zdnd11an1n64x5 FILLER_307_1708 ();
 b15zdnd11an1n64x5 FILLER_307_1772 ();
 b15zdnd11an1n64x5 FILLER_307_1836 ();
 b15zdnd11an1n64x5 FILLER_307_1900 ();
 b15zdnd11an1n64x5 FILLER_307_1964 ();
 b15zdnd11an1n64x5 FILLER_307_2028 ();
 b15zdnd11an1n64x5 FILLER_307_2092 ();
 b15zdnd11an1n64x5 FILLER_307_2156 ();
 b15zdnd11an1n64x5 FILLER_307_2220 ();
 b15zdnd11an1n64x5 FILLER_308_8 ();
 b15zdnd11an1n64x5 FILLER_308_72 ();
 b15zdnd11an1n64x5 FILLER_308_136 ();
 b15zdnd11an1n64x5 FILLER_308_200 ();
 b15zdnd11an1n64x5 FILLER_308_264 ();
 b15zdnd11an1n64x5 FILLER_308_328 ();
 b15zdnd11an1n64x5 FILLER_308_392 ();
 b15zdnd11an1n64x5 FILLER_308_456 ();
 b15zdnd11an1n64x5 FILLER_308_520 ();
 b15zdnd11an1n64x5 FILLER_308_584 ();
 b15zdnd11an1n64x5 FILLER_308_648 ();
 b15zdnd11an1n04x5 FILLER_308_712 ();
 b15zdnd00an1n02x5 FILLER_308_716 ();
 b15zdnd11an1n64x5 FILLER_308_726 ();
 b15zdnd11an1n32x5 FILLER_308_790 ();
 b15zdnd11an1n16x5 FILLER_308_822 ();
 b15zdnd00an1n01x5 FILLER_308_838 ();
 b15zdnd11an1n64x5 FILLER_308_881 ();
 b15zdnd11an1n64x5 FILLER_308_945 ();
 b15zdnd11an1n64x5 FILLER_308_1009 ();
 b15zdnd11an1n64x5 FILLER_308_1073 ();
 b15zdnd11an1n64x5 FILLER_308_1137 ();
 b15zdnd11an1n64x5 FILLER_308_1201 ();
 b15zdnd11an1n64x5 FILLER_308_1265 ();
 b15zdnd11an1n64x5 FILLER_308_1329 ();
 b15zdnd11an1n64x5 FILLER_308_1393 ();
 b15zdnd11an1n64x5 FILLER_308_1457 ();
 b15zdnd11an1n64x5 FILLER_308_1521 ();
 b15zdnd11an1n64x5 FILLER_308_1585 ();
 b15zdnd11an1n64x5 FILLER_308_1649 ();
 b15zdnd11an1n64x5 FILLER_308_1713 ();
 b15zdnd11an1n64x5 FILLER_308_1777 ();
 b15zdnd11an1n64x5 FILLER_308_1841 ();
 b15zdnd11an1n64x5 FILLER_308_1905 ();
 b15zdnd11an1n64x5 FILLER_308_1969 ();
 b15zdnd11an1n64x5 FILLER_308_2033 ();
 b15zdnd11an1n32x5 FILLER_308_2097 ();
 b15zdnd11an1n16x5 FILLER_308_2129 ();
 b15zdnd11an1n08x5 FILLER_308_2145 ();
 b15zdnd00an1n01x5 FILLER_308_2153 ();
 b15zdnd11an1n64x5 FILLER_308_2162 ();
 b15zdnd11an1n32x5 FILLER_308_2226 ();
 b15zdnd11an1n16x5 FILLER_308_2258 ();
 b15zdnd00an1n02x5 FILLER_308_2274 ();
 b15zdnd11an1n64x5 FILLER_309_0 ();
 b15zdnd11an1n64x5 FILLER_309_64 ();
 b15zdnd11an1n64x5 FILLER_309_128 ();
 b15zdnd11an1n64x5 FILLER_309_192 ();
 b15zdnd11an1n64x5 FILLER_309_256 ();
 b15zdnd11an1n64x5 FILLER_309_320 ();
 b15zdnd11an1n64x5 FILLER_309_384 ();
 b15zdnd11an1n64x5 FILLER_309_448 ();
 b15zdnd11an1n64x5 FILLER_309_512 ();
 b15zdnd11an1n64x5 FILLER_309_576 ();
 b15zdnd11an1n64x5 FILLER_309_640 ();
 b15zdnd11an1n64x5 FILLER_309_704 ();
 b15zdnd11an1n64x5 FILLER_309_768 ();
 b15zdnd11an1n64x5 FILLER_309_832 ();
 b15zdnd11an1n64x5 FILLER_309_896 ();
 b15zdnd11an1n64x5 FILLER_309_960 ();
 b15zdnd11an1n64x5 FILLER_309_1024 ();
 b15zdnd11an1n64x5 FILLER_309_1088 ();
 b15zdnd11an1n64x5 FILLER_309_1152 ();
 b15zdnd11an1n64x5 FILLER_309_1216 ();
 b15zdnd11an1n64x5 FILLER_309_1280 ();
 b15zdnd11an1n64x5 FILLER_309_1344 ();
 b15zdnd11an1n64x5 FILLER_309_1408 ();
 b15zdnd11an1n64x5 FILLER_309_1472 ();
 b15zdnd11an1n64x5 FILLER_309_1536 ();
 b15zdnd11an1n64x5 FILLER_309_1600 ();
 b15zdnd11an1n64x5 FILLER_309_1664 ();
 b15zdnd11an1n64x5 FILLER_309_1728 ();
 b15zdnd11an1n64x5 FILLER_309_1792 ();
 b15zdnd11an1n64x5 FILLER_309_1856 ();
 b15zdnd11an1n64x5 FILLER_309_1920 ();
 b15zdnd11an1n64x5 FILLER_309_1984 ();
 b15zdnd11an1n64x5 FILLER_309_2048 ();
 b15zdnd11an1n64x5 FILLER_309_2112 ();
 b15zdnd11an1n64x5 FILLER_309_2176 ();
 b15zdnd11an1n32x5 FILLER_309_2240 ();
 b15zdnd11an1n08x5 FILLER_309_2272 ();
 b15zdnd11an1n04x5 FILLER_309_2280 ();
 b15zdnd11an1n64x5 FILLER_310_8 ();
 b15zdnd11an1n64x5 FILLER_310_72 ();
 b15zdnd11an1n64x5 FILLER_310_136 ();
 b15zdnd11an1n64x5 FILLER_310_200 ();
 b15zdnd11an1n64x5 FILLER_310_264 ();
 b15zdnd11an1n64x5 FILLER_310_328 ();
 b15zdnd11an1n64x5 FILLER_310_392 ();
 b15zdnd11an1n64x5 FILLER_310_456 ();
 b15zdnd11an1n64x5 FILLER_310_520 ();
 b15zdnd11an1n64x5 FILLER_310_584 ();
 b15zdnd11an1n64x5 FILLER_310_648 ();
 b15zdnd11an1n04x5 FILLER_310_712 ();
 b15zdnd00an1n02x5 FILLER_310_716 ();
 b15zdnd11an1n64x5 FILLER_310_726 ();
 b15zdnd11an1n64x5 FILLER_310_790 ();
 b15zdnd11an1n64x5 FILLER_310_854 ();
 b15zdnd11an1n64x5 FILLER_310_918 ();
 b15zdnd11an1n64x5 FILLER_310_982 ();
 b15zdnd11an1n64x5 FILLER_310_1046 ();
 b15zdnd11an1n64x5 FILLER_310_1110 ();
 b15zdnd11an1n64x5 FILLER_310_1174 ();
 b15zdnd11an1n64x5 FILLER_310_1238 ();
 b15zdnd11an1n64x5 FILLER_310_1302 ();
 b15zdnd11an1n64x5 FILLER_310_1366 ();
 b15zdnd11an1n64x5 FILLER_310_1430 ();
 b15zdnd11an1n64x5 FILLER_310_1494 ();
 b15zdnd11an1n64x5 FILLER_310_1558 ();
 b15zdnd11an1n64x5 FILLER_310_1622 ();
 b15zdnd11an1n64x5 FILLER_310_1686 ();
 b15zdnd11an1n64x5 FILLER_310_1750 ();
 b15zdnd11an1n64x5 FILLER_310_1814 ();
 b15zdnd11an1n64x5 FILLER_310_1878 ();
 b15zdnd11an1n64x5 FILLER_310_1942 ();
 b15zdnd11an1n64x5 FILLER_310_2006 ();
 b15zdnd11an1n64x5 FILLER_310_2070 ();
 b15zdnd11an1n16x5 FILLER_310_2134 ();
 b15zdnd11an1n04x5 FILLER_310_2150 ();
 b15zdnd11an1n64x5 FILLER_310_2162 ();
 b15zdnd11an1n32x5 FILLER_310_2226 ();
 b15zdnd11an1n16x5 FILLER_310_2258 ();
 b15zdnd00an1n02x5 FILLER_310_2274 ();
 b15zdnd11an1n64x5 FILLER_311_0 ();
 b15zdnd11an1n64x5 FILLER_311_64 ();
 b15zdnd11an1n64x5 FILLER_311_128 ();
 b15zdnd11an1n64x5 FILLER_311_192 ();
 b15zdnd11an1n64x5 FILLER_311_256 ();
 b15zdnd11an1n64x5 FILLER_311_320 ();
 b15zdnd11an1n64x5 FILLER_311_384 ();
 b15zdnd11an1n64x5 FILLER_311_448 ();
 b15zdnd11an1n64x5 FILLER_311_512 ();
 b15zdnd11an1n64x5 FILLER_311_576 ();
 b15zdnd11an1n64x5 FILLER_311_640 ();
 b15zdnd11an1n64x5 FILLER_311_704 ();
 b15zdnd11an1n64x5 FILLER_311_768 ();
 b15zdnd11an1n64x5 FILLER_311_832 ();
 b15zdnd11an1n64x5 FILLER_311_896 ();
 b15zdnd11an1n64x5 FILLER_311_960 ();
 b15zdnd11an1n64x5 FILLER_311_1024 ();
 b15zdnd11an1n64x5 FILLER_311_1088 ();
 b15zdnd11an1n64x5 FILLER_311_1152 ();
 b15zdnd11an1n64x5 FILLER_311_1216 ();
 b15zdnd11an1n64x5 FILLER_311_1280 ();
 b15zdnd11an1n64x5 FILLER_311_1344 ();
 b15zdnd11an1n64x5 FILLER_311_1408 ();
 b15zdnd11an1n64x5 FILLER_311_1472 ();
 b15zdnd11an1n64x5 FILLER_311_1536 ();
 b15zdnd11an1n64x5 FILLER_311_1600 ();
 b15zdnd11an1n64x5 FILLER_311_1664 ();
 b15zdnd11an1n64x5 FILLER_311_1728 ();
 b15zdnd11an1n64x5 FILLER_311_1792 ();
 b15zdnd11an1n64x5 FILLER_311_1856 ();
 b15zdnd11an1n64x5 FILLER_311_1920 ();
 b15zdnd11an1n64x5 FILLER_311_1984 ();
 b15zdnd11an1n64x5 FILLER_311_2048 ();
 b15zdnd11an1n64x5 FILLER_311_2112 ();
 b15zdnd11an1n64x5 FILLER_311_2176 ();
 b15zdnd11an1n32x5 FILLER_311_2240 ();
 b15zdnd11an1n08x5 FILLER_311_2272 ();
 b15zdnd11an1n04x5 FILLER_311_2280 ();
 b15zdnd11an1n64x5 FILLER_312_8 ();
 b15zdnd11an1n64x5 FILLER_312_72 ();
 b15zdnd11an1n64x5 FILLER_312_136 ();
 b15zdnd11an1n64x5 FILLER_312_200 ();
 b15zdnd11an1n64x5 FILLER_312_264 ();
 b15zdnd11an1n64x5 FILLER_312_328 ();
 b15zdnd11an1n64x5 FILLER_312_392 ();
 b15zdnd11an1n64x5 FILLER_312_456 ();
 b15zdnd11an1n64x5 FILLER_312_520 ();
 b15zdnd11an1n64x5 FILLER_312_584 ();
 b15zdnd11an1n64x5 FILLER_312_648 ();
 b15zdnd11an1n04x5 FILLER_312_712 ();
 b15zdnd00an1n02x5 FILLER_312_716 ();
 b15zdnd11an1n64x5 FILLER_312_726 ();
 b15zdnd11an1n64x5 FILLER_312_790 ();
 b15zdnd11an1n64x5 FILLER_312_854 ();
 b15zdnd11an1n64x5 FILLER_312_918 ();
 b15zdnd11an1n64x5 FILLER_312_982 ();
 b15zdnd11an1n64x5 FILLER_312_1046 ();
 b15zdnd11an1n64x5 FILLER_312_1110 ();
 b15zdnd11an1n64x5 FILLER_312_1174 ();
 b15zdnd11an1n64x5 FILLER_312_1238 ();
 b15zdnd11an1n64x5 FILLER_312_1302 ();
 b15zdnd11an1n64x5 FILLER_312_1366 ();
 b15zdnd11an1n64x5 FILLER_312_1430 ();
 b15zdnd11an1n64x5 FILLER_312_1494 ();
 b15zdnd11an1n64x5 FILLER_312_1558 ();
 b15zdnd11an1n64x5 FILLER_312_1622 ();
 b15zdnd11an1n64x5 FILLER_312_1686 ();
 b15zdnd11an1n64x5 FILLER_312_1750 ();
 b15zdnd11an1n64x5 FILLER_312_1814 ();
 b15zdnd11an1n64x5 FILLER_312_1878 ();
 b15zdnd11an1n64x5 FILLER_312_1942 ();
 b15zdnd11an1n64x5 FILLER_312_2006 ();
 b15zdnd11an1n64x5 FILLER_312_2070 ();
 b15zdnd11an1n16x5 FILLER_312_2134 ();
 b15zdnd11an1n04x5 FILLER_312_2150 ();
 b15zdnd11an1n64x5 FILLER_312_2162 ();
 b15zdnd11an1n32x5 FILLER_312_2226 ();
 b15zdnd11an1n16x5 FILLER_312_2258 ();
 b15zdnd00an1n02x5 FILLER_312_2274 ();
 b15zdnd11an1n64x5 FILLER_313_0 ();
 b15zdnd11an1n64x5 FILLER_313_64 ();
 b15zdnd11an1n64x5 FILLER_313_128 ();
 b15zdnd11an1n64x5 FILLER_313_192 ();
 b15zdnd11an1n64x5 FILLER_313_256 ();
 b15zdnd11an1n64x5 FILLER_313_320 ();
 b15zdnd11an1n64x5 FILLER_313_384 ();
 b15zdnd11an1n64x5 FILLER_313_448 ();
 b15zdnd11an1n64x5 FILLER_313_512 ();
 b15zdnd11an1n64x5 FILLER_313_576 ();
 b15zdnd11an1n64x5 FILLER_313_640 ();
 b15zdnd11an1n64x5 FILLER_313_704 ();
 b15zdnd11an1n64x5 FILLER_313_768 ();
 b15zdnd11an1n64x5 FILLER_313_832 ();
 b15zdnd11an1n64x5 FILLER_313_896 ();
 b15zdnd11an1n64x5 FILLER_313_960 ();
 b15zdnd11an1n64x5 FILLER_313_1024 ();
 b15zdnd11an1n64x5 FILLER_313_1088 ();
 b15zdnd11an1n64x5 FILLER_313_1152 ();
 b15zdnd11an1n64x5 FILLER_313_1216 ();
 b15zdnd11an1n64x5 FILLER_313_1280 ();
 b15zdnd11an1n64x5 FILLER_313_1344 ();
 b15zdnd11an1n64x5 FILLER_313_1408 ();
 b15zdnd11an1n64x5 FILLER_313_1472 ();
 b15zdnd11an1n64x5 FILLER_313_1536 ();
 b15zdnd11an1n64x5 FILLER_313_1600 ();
 b15zdnd11an1n64x5 FILLER_313_1664 ();
 b15zdnd11an1n64x5 FILLER_313_1728 ();
 b15zdnd11an1n64x5 FILLER_313_1792 ();
 b15zdnd11an1n64x5 FILLER_313_1856 ();
 b15zdnd11an1n64x5 FILLER_313_1920 ();
 b15zdnd11an1n64x5 FILLER_313_1984 ();
 b15zdnd11an1n64x5 FILLER_313_2048 ();
 b15zdnd11an1n64x5 FILLER_313_2112 ();
 b15zdnd11an1n64x5 FILLER_313_2176 ();
 b15zdnd11an1n32x5 FILLER_313_2240 ();
 b15zdnd11an1n08x5 FILLER_313_2272 ();
 b15zdnd11an1n04x5 FILLER_313_2280 ();
 b15zdnd11an1n64x5 FILLER_314_8 ();
 b15zdnd11an1n64x5 FILLER_314_72 ();
 b15zdnd11an1n64x5 FILLER_314_136 ();
 b15zdnd11an1n64x5 FILLER_314_200 ();
 b15zdnd11an1n64x5 FILLER_314_264 ();
 b15zdnd11an1n64x5 FILLER_314_328 ();
 b15zdnd11an1n64x5 FILLER_314_392 ();
 b15zdnd11an1n64x5 FILLER_314_456 ();
 b15zdnd11an1n64x5 FILLER_314_520 ();
 b15zdnd11an1n64x5 FILLER_314_584 ();
 b15zdnd11an1n64x5 FILLER_314_648 ();
 b15zdnd11an1n04x5 FILLER_314_712 ();
 b15zdnd00an1n02x5 FILLER_314_716 ();
 b15zdnd11an1n64x5 FILLER_314_726 ();
 b15zdnd11an1n64x5 FILLER_314_790 ();
 b15zdnd11an1n64x5 FILLER_314_854 ();
 b15zdnd11an1n64x5 FILLER_314_918 ();
 b15zdnd11an1n64x5 FILLER_314_982 ();
 b15zdnd11an1n64x5 FILLER_314_1046 ();
 b15zdnd11an1n64x5 FILLER_314_1110 ();
 b15zdnd11an1n64x5 FILLER_314_1174 ();
 b15zdnd11an1n64x5 FILLER_314_1238 ();
 b15zdnd11an1n64x5 FILLER_314_1302 ();
 b15zdnd11an1n64x5 FILLER_314_1366 ();
 b15zdnd11an1n64x5 FILLER_314_1430 ();
 b15zdnd11an1n64x5 FILLER_314_1494 ();
 b15zdnd11an1n64x5 FILLER_314_1558 ();
 b15zdnd11an1n64x5 FILLER_314_1622 ();
 b15zdnd11an1n64x5 FILLER_314_1686 ();
 b15zdnd11an1n64x5 FILLER_314_1750 ();
 b15zdnd11an1n64x5 FILLER_314_1814 ();
 b15zdnd11an1n64x5 FILLER_314_1878 ();
 b15zdnd11an1n64x5 FILLER_314_1942 ();
 b15zdnd11an1n64x5 FILLER_314_2006 ();
 b15zdnd11an1n64x5 FILLER_314_2070 ();
 b15zdnd11an1n16x5 FILLER_314_2134 ();
 b15zdnd11an1n04x5 FILLER_314_2150 ();
 b15zdnd11an1n64x5 FILLER_314_2162 ();
 b15zdnd11an1n32x5 FILLER_314_2226 ();
 b15zdnd11an1n16x5 FILLER_314_2258 ();
 b15zdnd00an1n02x5 FILLER_314_2274 ();
 b15zdnd11an1n64x5 FILLER_315_0 ();
 b15zdnd11an1n64x5 FILLER_315_64 ();
 b15zdnd11an1n64x5 FILLER_315_128 ();
 b15zdnd11an1n64x5 FILLER_315_192 ();
 b15zdnd11an1n64x5 FILLER_315_256 ();
 b15zdnd11an1n64x5 FILLER_315_320 ();
 b15zdnd11an1n64x5 FILLER_315_384 ();
 b15zdnd11an1n64x5 FILLER_315_448 ();
 b15zdnd11an1n64x5 FILLER_315_512 ();
 b15zdnd11an1n64x5 FILLER_315_576 ();
 b15zdnd11an1n64x5 FILLER_315_640 ();
 b15zdnd11an1n64x5 FILLER_315_704 ();
 b15zdnd11an1n64x5 FILLER_315_768 ();
 b15zdnd11an1n64x5 FILLER_315_832 ();
 b15zdnd11an1n64x5 FILLER_315_896 ();
 b15zdnd11an1n64x5 FILLER_315_960 ();
 b15zdnd11an1n64x5 FILLER_315_1024 ();
 b15zdnd11an1n64x5 FILLER_315_1088 ();
 b15zdnd11an1n64x5 FILLER_315_1152 ();
 b15zdnd11an1n64x5 FILLER_315_1216 ();
 b15zdnd11an1n64x5 FILLER_315_1280 ();
 b15zdnd11an1n64x5 FILLER_315_1344 ();
 b15zdnd11an1n64x5 FILLER_315_1408 ();
 b15zdnd11an1n64x5 FILLER_315_1472 ();
 b15zdnd11an1n64x5 FILLER_315_1536 ();
 b15zdnd11an1n64x5 FILLER_315_1600 ();
 b15zdnd11an1n64x5 FILLER_315_1664 ();
 b15zdnd11an1n64x5 FILLER_315_1728 ();
 b15zdnd11an1n64x5 FILLER_315_1792 ();
 b15zdnd11an1n64x5 FILLER_315_1856 ();
 b15zdnd11an1n64x5 FILLER_315_1920 ();
 b15zdnd11an1n64x5 FILLER_315_1984 ();
 b15zdnd11an1n64x5 FILLER_315_2048 ();
 b15zdnd11an1n64x5 FILLER_315_2112 ();
 b15zdnd11an1n64x5 FILLER_315_2176 ();
 b15zdnd11an1n32x5 FILLER_315_2240 ();
 b15zdnd11an1n08x5 FILLER_315_2272 ();
 b15zdnd11an1n04x5 FILLER_315_2280 ();
 b15zdnd11an1n64x5 FILLER_316_8 ();
 b15zdnd11an1n64x5 FILLER_316_72 ();
 b15zdnd11an1n64x5 FILLER_316_136 ();
 b15zdnd11an1n64x5 FILLER_316_200 ();
 b15zdnd11an1n64x5 FILLER_316_264 ();
 b15zdnd11an1n64x5 FILLER_316_328 ();
 b15zdnd11an1n64x5 FILLER_316_392 ();
 b15zdnd11an1n64x5 FILLER_316_456 ();
 b15zdnd11an1n64x5 FILLER_316_520 ();
 b15zdnd11an1n64x5 FILLER_316_584 ();
 b15zdnd11an1n64x5 FILLER_316_648 ();
 b15zdnd11an1n04x5 FILLER_316_712 ();
 b15zdnd00an1n02x5 FILLER_316_716 ();
 b15zdnd11an1n64x5 FILLER_316_726 ();
 b15zdnd11an1n64x5 FILLER_316_790 ();
 b15zdnd11an1n16x5 FILLER_316_854 ();
 b15zdnd00an1n02x5 FILLER_316_870 ();
 b15zdnd00an1n01x5 FILLER_316_872 ();
 b15zdnd11an1n64x5 FILLER_316_915 ();
 b15zdnd11an1n64x5 FILLER_316_979 ();
 b15zdnd11an1n64x5 FILLER_316_1043 ();
 b15zdnd11an1n64x5 FILLER_316_1107 ();
 b15zdnd11an1n64x5 FILLER_316_1171 ();
 b15zdnd11an1n64x5 FILLER_316_1235 ();
 b15zdnd11an1n64x5 FILLER_316_1299 ();
 b15zdnd11an1n64x5 FILLER_316_1363 ();
 b15zdnd11an1n64x5 FILLER_316_1427 ();
 b15zdnd11an1n64x5 FILLER_316_1491 ();
 b15zdnd11an1n64x5 FILLER_316_1555 ();
 b15zdnd11an1n64x5 FILLER_316_1619 ();
 b15zdnd11an1n64x5 FILLER_316_1683 ();
 b15zdnd11an1n64x5 FILLER_316_1747 ();
 b15zdnd11an1n64x5 FILLER_316_1811 ();
 b15zdnd11an1n64x5 FILLER_316_1875 ();
 b15zdnd11an1n64x5 FILLER_316_1939 ();
 b15zdnd11an1n64x5 FILLER_316_2003 ();
 b15zdnd11an1n64x5 FILLER_316_2067 ();
 b15zdnd11an1n16x5 FILLER_316_2131 ();
 b15zdnd11an1n04x5 FILLER_316_2147 ();
 b15zdnd00an1n02x5 FILLER_316_2151 ();
 b15zdnd00an1n01x5 FILLER_316_2153 ();
 b15zdnd11an1n64x5 FILLER_316_2162 ();
 b15zdnd11an1n32x5 FILLER_316_2226 ();
 b15zdnd11an1n16x5 FILLER_316_2258 ();
 b15zdnd00an1n02x5 FILLER_316_2274 ();
 b15zdnd11an1n64x5 FILLER_317_0 ();
 b15zdnd11an1n64x5 FILLER_317_64 ();
 b15zdnd11an1n64x5 FILLER_317_128 ();
 b15zdnd11an1n64x5 FILLER_317_192 ();
 b15zdnd11an1n64x5 FILLER_317_256 ();
 b15zdnd11an1n64x5 FILLER_317_320 ();
 b15zdnd11an1n64x5 FILLER_317_384 ();
 b15zdnd11an1n64x5 FILLER_317_448 ();
 b15zdnd11an1n64x5 FILLER_317_512 ();
 b15zdnd11an1n64x5 FILLER_317_576 ();
 b15zdnd11an1n64x5 FILLER_317_640 ();
 b15zdnd11an1n64x5 FILLER_317_704 ();
 b15zdnd11an1n64x5 FILLER_317_768 ();
 b15zdnd11an1n64x5 FILLER_317_832 ();
 b15zdnd11an1n64x5 FILLER_317_896 ();
 b15zdnd11an1n64x5 FILLER_317_960 ();
 b15zdnd11an1n64x5 FILLER_317_1024 ();
 b15zdnd11an1n64x5 FILLER_317_1088 ();
 b15zdnd11an1n64x5 FILLER_317_1152 ();
 b15zdnd11an1n64x5 FILLER_317_1216 ();
 b15zdnd11an1n64x5 FILLER_317_1280 ();
 b15zdnd11an1n64x5 FILLER_317_1344 ();
 b15zdnd11an1n64x5 FILLER_317_1408 ();
 b15zdnd11an1n64x5 FILLER_317_1472 ();
 b15zdnd11an1n64x5 FILLER_317_1536 ();
 b15zdnd11an1n64x5 FILLER_317_1600 ();
 b15zdnd11an1n64x5 FILLER_317_1664 ();
 b15zdnd11an1n64x5 FILLER_317_1728 ();
 b15zdnd11an1n64x5 FILLER_317_1792 ();
 b15zdnd11an1n64x5 FILLER_317_1856 ();
 b15zdnd11an1n64x5 FILLER_317_1920 ();
 b15zdnd11an1n64x5 FILLER_317_1984 ();
 b15zdnd11an1n64x5 FILLER_317_2048 ();
 b15zdnd11an1n64x5 FILLER_317_2112 ();
 b15zdnd11an1n64x5 FILLER_317_2176 ();
 b15zdnd11an1n32x5 FILLER_317_2240 ();
 b15zdnd11an1n08x5 FILLER_317_2272 ();
 b15zdnd11an1n04x5 FILLER_317_2280 ();
 b15zdnd11an1n64x5 FILLER_318_8 ();
 b15zdnd11an1n64x5 FILLER_318_72 ();
 b15zdnd11an1n64x5 FILLER_318_136 ();
 b15zdnd11an1n64x5 FILLER_318_200 ();
 b15zdnd11an1n64x5 FILLER_318_264 ();
 b15zdnd11an1n64x5 FILLER_318_328 ();
 b15zdnd11an1n64x5 FILLER_318_392 ();
 b15zdnd11an1n64x5 FILLER_318_456 ();
 b15zdnd11an1n64x5 FILLER_318_520 ();
 b15zdnd11an1n64x5 FILLER_318_584 ();
 b15zdnd11an1n64x5 FILLER_318_648 ();
 b15zdnd11an1n04x5 FILLER_318_712 ();
 b15zdnd00an1n02x5 FILLER_318_716 ();
 b15zdnd11an1n64x5 FILLER_318_726 ();
 b15zdnd11an1n64x5 FILLER_318_790 ();
 b15zdnd11an1n64x5 FILLER_318_854 ();
 b15zdnd11an1n64x5 FILLER_318_918 ();
 b15zdnd11an1n64x5 FILLER_318_982 ();
 b15zdnd11an1n64x5 FILLER_318_1046 ();
 b15zdnd11an1n64x5 FILLER_318_1110 ();
 b15zdnd11an1n64x5 FILLER_318_1174 ();
 b15zdnd11an1n64x5 FILLER_318_1238 ();
 b15zdnd11an1n64x5 FILLER_318_1302 ();
 b15zdnd11an1n64x5 FILLER_318_1366 ();
 b15zdnd11an1n64x5 FILLER_318_1430 ();
 b15zdnd11an1n64x5 FILLER_318_1494 ();
 b15zdnd11an1n64x5 FILLER_318_1558 ();
 b15zdnd11an1n64x5 FILLER_318_1622 ();
 b15zdnd11an1n64x5 FILLER_318_1686 ();
 b15zdnd11an1n64x5 FILLER_318_1750 ();
 b15zdnd11an1n64x5 FILLER_318_1814 ();
 b15zdnd11an1n64x5 FILLER_318_1878 ();
 b15zdnd11an1n64x5 FILLER_318_1942 ();
 b15zdnd11an1n64x5 FILLER_318_2006 ();
 b15zdnd11an1n64x5 FILLER_318_2070 ();
 b15zdnd11an1n16x5 FILLER_318_2134 ();
 b15zdnd11an1n04x5 FILLER_318_2150 ();
 b15zdnd11an1n64x5 FILLER_318_2162 ();
 b15zdnd11an1n32x5 FILLER_318_2226 ();
 b15zdnd11an1n16x5 FILLER_318_2258 ();
 b15zdnd00an1n02x5 FILLER_318_2274 ();
 b15zdnd11an1n64x5 FILLER_319_0 ();
 b15zdnd11an1n64x5 FILLER_319_64 ();
 b15zdnd11an1n64x5 FILLER_319_128 ();
 b15zdnd11an1n64x5 FILLER_319_192 ();
 b15zdnd11an1n64x5 FILLER_319_256 ();
 b15zdnd11an1n64x5 FILLER_319_320 ();
 b15zdnd11an1n64x5 FILLER_319_384 ();
 b15zdnd11an1n64x5 FILLER_319_448 ();
 b15zdnd11an1n64x5 FILLER_319_512 ();
 b15zdnd11an1n64x5 FILLER_319_576 ();
 b15zdnd11an1n64x5 FILLER_319_640 ();
 b15zdnd11an1n64x5 FILLER_319_704 ();
 b15zdnd11an1n64x5 FILLER_319_768 ();
 b15zdnd11an1n64x5 FILLER_319_832 ();
 b15zdnd11an1n64x5 FILLER_319_896 ();
 b15zdnd11an1n64x5 FILLER_319_960 ();
 b15zdnd11an1n64x5 FILLER_319_1024 ();
 b15zdnd11an1n64x5 FILLER_319_1088 ();
 b15zdnd11an1n64x5 FILLER_319_1152 ();
 b15zdnd11an1n64x5 FILLER_319_1216 ();
 b15zdnd11an1n64x5 FILLER_319_1280 ();
 b15zdnd11an1n64x5 FILLER_319_1344 ();
 b15zdnd11an1n64x5 FILLER_319_1408 ();
 b15zdnd11an1n64x5 FILLER_319_1472 ();
 b15zdnd11an1n64x5 FILLER_319_1536 ();
 b15zdnd11an1n64x5 FILLER_319_1600 ();
 b15zdnd11an1n64x5 FILLER_319_1664 ();
 b15zdnd11an1n64x5 FILLER_319_1728 ();
 b15zdnd11an1n64x5 FILLER_319_1792 ();
 b15zdnd11an1n64x5 FILLER_319_1856 ();
 b15zdnd11an1n64x5 FILLER_319_1920 ();
 b15zdnd11an1n64x5 FILLER_319_1984 ();
 b15zdnd11an1n64x5 FILLER_319_2048 ();
 b15zdnd11an1n64x5 FILLER_319_2112 ();
 b15zdnd11an1n64x5 FILLER_319_2176 ();
 b15zdnd11an1n32x5 FILLER_319_2240 ();
 b15zdnd11an1n08x5 FILLER_319_2272 ();
 b15zdnd11an1n04x5 FILLER_319_2280 ();
 b15zdnd11an1n64x5 FILLER_320_8 ();
 b15zdnd11an1n64x5 FILLER_320_72 ();
 b15zdnd11an1n64x5 FILLER_320_136 ();
 b15zdnd11an1n64x5 FILLER_320_200 ();
 b15zdnd11an1n64x5 FILLER_320_264 ();
 b15zdnd11an1n64x5 FILLER_320_328 ();
 b15zdnd11an1n64x5 FILLER_320_392 ();
 b15zdnd11an1n64x5 FILLER_320_456 ();
 b15zdnd11an1n64x5 FILLER_320_520 ();
 b15zdnd11an1n64x5 FILLER_320_584 ();
 b15zdnd11an1n64x5 FILLER_320_648 ();
 b15zdnd11an1n04x5 FILLER_320_712 ();
 b15zdnd00an1n02x5 FILLER_320_716 ();
 b15zdnd11an1n64x5 FILLER_320_726 ();
 b15zdnd11an1n64x5 FILLER_320_790 ();
 b15zdnd11an1n64x5 FILLER_320_854 ();
 b15zdnd11an1n64x5 FILLER_320_918 ();
 b15zdnd11an1n64x5 FILLER_320_982 ();
 b15zdnd11an1n64x5 FILLER_320_1046 ();
 b15zdnd11an1n64x5 FILLER_320_1110 ();
 b15zdnd11an1n64x5 FILLER_320_1174 ();
 b15zdnd11an1n64x5 FILLER_320_1238 ();
 b15zdnd11an1n64x5 FILLER_320_1302 ();
 b15zdnd11an1n64x5 FILLER_320_1366 ();
 b15zdnd11an1n64x5 FILLER_320_1430 ();
 b15zdnd11an1n64x5 FILLER_320_1494 ();
 b15zdnd11an1n64x5 FILLER_320_1558 ();
 b15zdnd11an1n64x5 FILLER_320_1622 ();
 b15zdnd11an1n64x5 FILLER_320_1686 ();
 b15zdnd11an1n64x5 FILLER_320_1750 ();
 b15zdnd11an1n64x5 FILLER_320_1814 ();
 b15zdnd11an1n64x5 FILLER_320_1878 ();
 b15zdnd11an1n64x5 FILLER_320_1942 ();
 b15zdnd11an1n64x5 FILLER_320_2006 ();
 b15zdnd11an1n64x5 FILLER_320_2070 ();
 b15zdnd11an1n16x5 FILLER_320_2134 ();
 b15zdnd11an1n04x5 FILLER_320_2150 ();
 b15zdnd11an1n64x5 FILLER_320_2162 ();
 b15zdnd11an1n32x5 FILLER_320_2226 ();
 b15zdnd11an1n16x5 FILLER_320_2258 ();
 b15zdnd00an1n02x5 FILLER_320_2274 ();
 b15zdnd11an1n64x5 FILLER_321_0 ();
 b15zdnd11an1n64x5 FILLER_321_64 ();
 b15zdnd11an1n64x5 FILLER_321_128 ();
 b15zdnd11an1n64x5 FILLER_321_192 ();
 b15zdnd11an1n64x5 FILLER_321_256 ();
 b15zdnd11an1n64x5 FILLER_321_320 ();
 b15zdnd11an1n64x5 FILLER_321_384 ();
 b15zdnd11an1n64x5 FILLER_321_448 ();
 b15zdnd11an1n64x5 FILLER_321_512 ();
 b15zdnd11an1n64x5 FILLER_321_576 ();
 b15zdnd11an1n64x5 FILLER_321_640 ();
 b15zdnd11an1n64x5 FILLER_321_704 ();
 b15zdnd11an1n64x5 FILLER_321_768 ();
 b15zdnd11an1n64x5 FILLER_321_832 ();
 b15zdnd11an1n64x5 FILLER_321_896 ();
 b15zdnd11an1n64x5 FILLER_321_960 ();
 b15zdnd11an1n64x5 FILLER_321_1024 ();
 b15zdnd11an1n64x5 FILLER_321_1088 ();
 b15zdnd11an1n64x5 FILLER_321_1152 ();
 b15zdnd11an1n64x5 FILLER_321_1216 ();
 b15zdnd11an1n64x5 FILLER_321_1280 ();
 b15zdnd11an1n64x5 FILLER_321_1344 ();
 b15zdnd11an1n64x5 FILLER_321_1408 ();
 b15zdnd11an1n64x5 FILLER_321_1472 ();
 b15zdnd11an1n64x5 FILLER_321_1536 ();
 b15zdnd11an1n64x5 FILLER_321_1600 ();
 b15zdnd11an1n64x5 FILLER_321_1664 ();
 b15zdnd11an1n64x5 FILLER_321_1728 ();
 b15zdnd11an1n64x5 FILLER_321_1792 ();
 b15zdnd11an1n64x5 FILLER_321_1856 ();
 b15zdnd11an1n64x5 FILLER_321_1920 ();
 b15zdnd11an1n64x5 FILLER_321_1984 ();
 b15zdnd11an1n64x5 FILLER_321_2048 ();
 b15zdnd11an1n64x5 FILLER_321_2112 ();
 b15zdnd11an1n64x5 FILLER_321_2176 ();
 b15zdnd11an1n32x5 FILLER_321_2240 ();
 b15zdnd11an1n08x5 FILLER_321_2272 ();
 b15zdnd11an1n04x5 FILLER_321_2280 ();
 b15zdnd11an1n64x5 FILLER_322_8 ();
 b15zdnd11an1n64x5 FILLER_322_72 ();
 b15zdnd11an1n64x5 FILLER_322_136 ();
 b15zdnd11an1n64x5 FILLER_322_200 ();
 b15zdnd11an1n64x5 FILLER_322_264 ();
 b15zdnd11an1n64x5 FILLER_322_328 ();
 b15zdnd11an1n64x5 FILLER_322_392 ();
 b15zdnd11an1n64x5 FILLER_322_456 ();
 b15zdnd11an1n64x5 FILLER_322_520 ();
 b15zdnd11an1n64x5 FILLER_322_584 ();
 b15zdnd11an1n64x5 FILLER_322_648 ();
 b15zdnd11an1n04x5 FILLER_322_712 ();
 b15zdnd00an1n02x5 FILLER_322_716 ();
 b15zdnd11an1n64x5 FILLER_322_726 ();
 b15zdnd11an1n64x5 FILLER_322_790 ();
 b15zdnd11an1n64x5 FILLER_322_854 ();
 b15zdnd11an1n64x5 FILLER_322_918 ();
 b15zdnd11an1n64x5 FILLER_322_982 ();
 b15zdnd11an1n64x5 FILLER_322_1046 ();
 b15zdnd11an1n64x5 FILLER_322_1110 ();
 b15zdnd11an1n64x5 FILLER_322_1174 ();
 b15zdnd11an1n32x5 FILLER_322_1238 ();
 b15zdnd11an1n16x5 FILLER_322_1270 ();
 b15zdnd11an1n08x5 FILLER_322_1286 ();
 b15zdnd11an1n04x5 FILLER_322_1294 ();
 b15zdnd00an1n01x5 FILLER_322_1298 ();
 b15zdnd11an1n64x5 FILLER_322_1341 ();
 b15zdnd11an1n64x5 FILLER_322_1405 ();
 b15zdnd11an1n64x5 FILLER_322_1469 ();
 b15zdnd11an1n64x5 FILLER_322_1533 ();
 b15zdnd11an1n64x5 FILLER_322_1597 ();
 b15zdnd11an1n64x5 FILLER_322_1661 ();
 b15zdnd11an1n64x5 FILLER_322_1725 ();
 b15zdnd11an1n64x5 FILLER_322_1789 ();
 b15zdnd11an1n64x5 FILLER_322_1853 ();
 b15zdnd11an1n64x5 FILLER_322_1917 ();
 b15zdnd11an1n64x5 FILLER_322_1981 ();
 b15zdnd11an1n64x5 FILLER_322_2045 ();
 b15zdnd11an1n32x5 FILLER_322_2109 ();
 b15zdnd11an1n08x5 FILLER_322_2141 ();
 b15zdnd11an1n04x5 FILLER_322_2149 ();
 b15zdnd00an1n01x5 FILLER_322_2153 ();
 b15zdnd11an1n64x5 FILLER_322_2162 ();
 b15zdnd11an1n32x5 FILLER_322_2226 ();
 b15zdnd11an1n16x5 FILLER_322_2258 ();
 b15zdnd00an1n02x5 FILLER_322_2274 ();
 b15zdnd11an1n64x5 FILLER_323_0 ();
 b15zdnd11an1n64x5 FILLER_323_64 ();
 b15zdnd11an1n64x5 FILLER_323_128 ();
 b15zdnd11an1n64x5 FILLER_323_192 ();
 b15zdnd11an1n64x5 FILLER_323_256 ();
 b15zdnd11an1n64x5 FILLER_323_320 ();
 b15zdnd11an1n64x5 FILLER_323_384 ();
 b15zdnd11an1n64x5 FILLER_323_448 ();
 b15zdnd11an1n64x5 FILLER_323_512 ();
 b15zdnd11an1n64x5 FILLER_323_576 ();
 b15zdnd11an1n64x5 FILLER_323_640 ();
 b15zdnd11an1n64x5 FILLER_323_704 ();
 b15zdnd11an1n64x5 FILLER_323_768 ();
 b15zdnd11an1n64x5 FILLER_323_832 ();
 b15zdnd11an1n64x5 FILLER_323_896 ();
 b15zdnd11an1n64x5 FILLER_323_960 ();
 b15zdnd11an1n64x5 FILLER_323_1024 ();
 b15zdnd11an1n64x5 FILLER_323_1088 ();
 b15zdnd11an1n64x5 FILLER_323_1152 ();
 b15zdnd11an1n32x5 FILLER_323_1216 ();
 b15zdnd11an1n16x5 FILLER_323_1248 ();
 b15zdnd11an1n08x5 FILLER_323_1264 ();
 b15zdnd11an1n04x5 FILLER_323_1272 ();
 b15zdnd00an1n02x5 FILLER_323_1276 ();
 b15zdnd11an1n64x5 FILLER_323_1320 ();
 b15zdnd11an1n64x5 FILLER_323_1384 ();
 b15zdnd11an1n64x5 FILLER_323_1448 ();
 b15zdnd11an1n64x5 FILLER_323_1512 ();
 b15zdnd11an1n64x5 FILLER_323_1576 ();
 b15zdnd11an1n64x5 FILLER_323_1640 ();
 b15zdnd11an1n64x5 FILLER_323_1704 ();
 b15zdnd11an1n64x5 FILLER_323_1768 ();
 b15zdnd11an1n64x5 FILLER_323_1832 ();
 b15zdnd11an1n64x5 FILLER_323_1896 ();
 b15zdnd11an1n64x5 FILLER_323_1960 ();
 b15zdnd11an1n64x5 FILLER_323_2024 ();
 b15zdnd11an1n64x5 FILLER_323_2088 ();
 b15zdnd11an1n64x5 FILLER_323_2152 ();
 b15zdnd11an1n64x5 FILLER_323_2216 ();
 b15zdnd11an1n04x5 FILLER_323_2280 ();
 b15zdnd11an1n64x5 FILLER_324_8 ();
 b15zdnd11an1n64x5 FILLER_324_72 ();
 b15zdnd11an1n64x5 FILLER_324_136 ();
 b15zdnd11an1n64x5 FILLER_324_200 ();
 b15zdnd11an1n64x5 FILLER_324_264 ();
 b15zdnd11an1n64x5 FILLER_324_328 ();
 b15zdnd11an1n64x5 FILLER_324_392 ();
 b15zdnd11an1n64x5 FILLER_324_456 ();
 b15zdnd11an1n64x5 FILLER_324_520 ();
 b15zdnd11an1n64x5 FILLER_324_584 ();
 b15zdnd11an1n64x5 FILLER_324_648 ();
 b15zdnd11an1n04x5 FILLER_324_712 ();
 b15zdnd00an1n02x5 FILLER_324_716 ();
 b15zdnd11an1n64x5 FILLER_324_726 ();
 b15zdnd11an1n64x5 FILLER_324_790 ();
 b15zdnd11an1n64x5 FILLER_324_854 ();
 b15zdnd11an1n64x5 FILLER_324_918 ();
 b15zdnd11an1n64x5 FILLER_324_982 ();
 b15zdnd11an1n64x5 FILLER_324_1046 ();
 b15zdnd11an1n64x5 FILLER_324_1110 ();
 b15zdnd11an1n64x5 FILLER_324_1174 ();
 b15zdnd11an1n64x5 FILLER_324_1238 ();
 b15zdnd11an1n64x5 FILLER_324_1302 ();
 b15zdnd11an1n64x5 FILLER_324_1366 ();
 b15zdnd11an1n64x5 FILLER_324_1430 ();
 b15zdnd11an1n64x5 FILLER_324_1494 ();
 b15zdnd11an1n64x5 FILLER_324_1558 ();
 b15zdnd11an1n64x5 FILLER_324_1622 ();
 b15zdnd11an1n64x5 FILLER_324_1686 ();
 b15zdnd11an1n64x5 FILLER_324_1750 ();
 b15zdnd11an1n64x5 FILLER_324_1814 ();
 b15zdnd11an1n64x5 FILLER_324_1878 ();
 b15zdnd11an1n64x5 FILLER_324_1942 ();
 b15zdnd11an1n64x5 FILLER_324_2006 ();
 b15zdnd11an1n64x5 FILLER_324_2070 ();
 b15zdnd11an1n16x5 FILLER_324_2134 ();
 b15zdnd11an1n04x5 FILLER_324_2150 ();
 b15zdnd11an1n64x5 FILLER_324_2162 ();
 b15zdnd11an1n32x5 FILLER_324_2226 ();
 b15zdnd11an1n16x5 FILLER_324_2258 ();
 b15zdnd00an1n02x5 FILLER_324_2274 ();
 b15zdnd11an1n64x5 FILLER_325_0 ();
 b15zdnd11an1n64x5 FILLER_325_64 ();
 b15zdnd11an1n64x5 FILLER_325_128 ();
 b15zdnd11an1n64x5 FILLER_325_192 ();
 b15zdnd11an1n64x5 FILLER_325_256 ();
 b15zdnd11an1n64x5 FILLER_325_320 ();
 b15zdnd11an1n64x5 FILLER_325_384 ();
 b15zdnd11an1n64x5 FILLER_325_448 ();
 b15zdnd11an1n64x5 FILLER_325_512 ();
 b15zdnd11an1n64x5 FILLER_325_576 ();
 b15zdnd11an1n64x5 FILLER_325_640 ();
 b15zdnd11an1n64x5 FILLER_325_704 ();
 b15zdnd11an1n64x5 FILLER_325_768 ();
 b15zdnd11an1n64x5 FILLER_325_832 ();
 b15zdnd11an1n64x5 FILLER_325_896 ();
 b15zdnd11an1n64x5 FILLER_325_960 ();
 b15zdnd11an1n64x5 FILLER_325_1024 ();
 b15zdnd11an1n64x5 FILLER_325_1088 ();
 b15zdnd11an1n64x5 FILLER_325_1152 ();
 b15zdnd11an1n64x5 FILLER_325_1216 ();
 b15zdnd11an1n64x5 FILLER_325_1280 ();
 b15zdnd11an1n64x5 FILLER_325_1344 ();
 b15zdnd11an1n64x5 FILLER_325_1408 ();
 b15zdnd11an1n64x5 FILLER_325_1472 ();
 b15zdnd11an1n64x5 FILLER_325_1536 ();
 b15zdnd11an1n64x5 FILLER_325_1600 ();
 b15zdnd11an1n64x5 FILLER_325_1664 ();
 b15zdnd11an1n64x5 FILLER_325_1728 ();
 b15zdnd11an1n64x5 FILLER_325_1792 ();
 b15zdnd11an1n64x5 FILLER_325_1856 ();
 b15zdnd11an1n64x5 FILLER_325_1920 ();
 b15zdnd11an1n64x5 FILLER_325_1984 ();
 b15zdnd11an1n64x5 FILLER_325_2048 ();
 b15zdnd11an1n64x5 FILLER_325_2112 ();
 b15zdnd11an1n64x5 FILLER_325_2176 ();
 b15zdnd11an1n32x5 FILLER_325_2240 ();
 b15zdnd11an1n08x5 FILLER_325_2272 ();
 b15zdnd11an1n04x5 FILLER_325_2280 ();
 b15zdnd11an1n64x5 FILLER_326_8 ();
 b15zdnd11an1n64x5 FILLER_326_72 ();
 b15zdnd11an1n64x5 FILLER_326_136 ();
 b15zdnd11an1n64x5 FILLER_326_200 ();
 b15zdnd11an1n64x5 FILLER_326_264 ();
 b15zdnd11an1n64x5 FILLER_326_328 ();
 b15zdnd11an1n64x5 FILLER_326_392 ();
 b15zdnd11an1n64x5 FILLER_326_456 ();
 b15zdnd11an1n64x5 FILLER_326_520 ();
 b15zdnd11an1n64x5 FILLER_326_584 ();
 b15zdnd11an1n64x5 FILLER_326_648 ();
 b15zdnd11an1n04x5 FILLER_326_712 ();
 b15zdnd00an1n02x5 FILLER_326_716 ();
 b15zdnd11an1n64x5 FILLER_326_726 ();
 b15zdnd11an1n64x5 FILLER_326_790 ();
 b15zdnd11an1n64x5 FILLER_326_854 ();
 b15zdnd11an1n64x5 FILLER_326_918 ();
 b15zdnd11an1n64x5 FILLER_326_982 ();
 b15zdnd11an1n64x5 FILLER_326_1046 ();
 b15zdnd11an1n64x5 FILLER_326_1110 ();
 b15zdnd11an1n64x5 FILLER_326_1174 ();
 b15zdnd11an1n64x5 FILLER_326_1238 ();
 b15zdnd11an1n64x5 FILLER_326_1302 ();
 b15zdnd11an1n64x5 FILLER_326_1366 ();
 b15zdnd11an1n64x5 FILLER_326_1430 ();
 b15zdnd11an1n64x5 FILLER_326_1494 ();
 b15zdnd11an1n64x5 FILLER_326_1558 ();
 b15zdnd11an1n64x5 FILLER_326_1622 ();
 b15zdnd11an1n64x5 FILLER_326_1686 ();
 b15zdnd11an1n64x5 FILLER_326_1750 ();
 b15zdnd11an1n64x5 FILLER_326_1814 ();
 b15zdnd11an1n64x5 FILLER_326_1878 ();
 b15zdnd11an1n64x5 FILLER_326_1942 ();
 b15zdnd11an1n64x5 FILLER_326_2006 ();
 b15zdnd11an1n64x5 FILLER_326_2070 ();
 b15zdnd11an1n16x5 FILLER_326_2134 ();
 b15zdnd11an1n04x5 FILLER_326_2150 ();
 b15zdnd11an1n64x5 FILLER_326_2162 ();
 b15zdnd11an1n32x5 FILLER_326_2226 ();
 b15zdnd11an1n16x5 FILLER_326_2258 ();
 b15zdnd00an1n02x5 FILLER_326_2274 ();
 b15zdnd11an1n64x5 FILLER_327_0 ();
 b15zdnd11an1n64x5 FILLER_327_64 ();
 b15zdnd11an1n64x5 FILLER_327_128 ();
 b15zdnd11an1n64x5 FILLER_327_192 ();
 b15zdnd11an1n64x5 FILLER_327_256 ();
 b15zdnd11an1n64x5 FILLER_327_320 ();
 b15zdnd11an1n64x5 FILLER_327_384 ();
 b15zdnd11an1n64x5 FILLER_327_448 ();
 b15zdnd11an1n64x5 FILLER_327_512 ();
 b15zdnd11an1n64x5 FILLER_327_576 ();
 b15zdnd11an1n64x5 FILLER_327_640 ();
 b15zdnd11an1n64x5 FILLER_327_704 ();
 b15zdnd11an1n64x5 FILLER_327_768 ();
 b15zdnd11an1n64x5 FILLER_327_832 ();
 b15zdnd11an1n64x5 FILLER_327_896 ();
 b15zdnd11an1n64x5 FILLER_327_960 ();
 b15zdnd11an1n64x5 FILLER_327_1024 ();
 b15zdnd11an1n64x5 FILLER_327_1088 ();
 b15zdnd11an1n64x5 FILLER_327_1152 ();
 b15zdnd11an1n64x5 FILLER_327_1216 ();
 b15zdnd11an1n64x5 FILLER_327_1280 ();
 b15zdnd11an1n64x5 FILLER_327_1344 ();
 b15zdnd11an1n64x5 FILLER_327_1408 ();
 b15zdnd11an1n64x5 FILLER_327_1472 ();
 b15zdnd11an1n64x5 FILLER_327_1536 ();
 b15zdnd11an1n64x5 FILLER_327_1600 ();
 b15zdnd11an1n64x5 FILLER_327_1664 ();
 b15zdnd11an1n64x5 FILLER_327_1728 ();
 b15zdnd11an1n64x5 FILLER_327_1792 ();
 b15zdnd11an1n64x5 FILLER_327_1856 ();
 b15zdnd11an1n64x5 FILLER_327_1920 ();
 b15zdnd11an1n64x5 FILLER_327_1984 ();
 b15zdnd11an1n64x5 FILLER_327_2048 ();
 b15zdnd11an1n64x5 FILLER_327_2112 ();
 b15zdnd11an1n64x5 FILLER_327_2176 ();
 b15zdnd11an1n32x5 FILLER_327_2240 ();
 b15zdnd11an1n08x5 FILLER_327_2272 ();
 b15zdnd11an1n04x5 FILLER_327_2280 ();
 b15zdnd11an1n64x5 FILLER_328_8 ();
 b15zdnd11an1n64x5 FILLER_328_72 ();
 b15zdnd11an1n64x5 FILLER_328_136 ();
 b15zdnd11an1n64x5 FILLER_328_200 ();
 b15zdnd11an1n64x5 FILLER_328_264 ();
 b15zdnd11an1n64x5 FILLER_328_328 ();
 b15zdnd11an1n64x5 FILLER_328_392 ();
 b15zdnd11an1n64x5 FILLER_328_456 ();
 b15zdnd11an1n64x5 FILLER_328_520 ();
 b15zdnd11an1n64x5 FILLER_328_584 ();
 b15zdnd11an1n64x5 FILLER_328_648 ();
 b15zdnd11an1n04x5 FILLER_328_712 ();
 b15zdnd00an1n02x5 FILLER_328_716 ();
 b15zdnd11an1n64x5 FILLER_328_726 ();
 b15zdnd11an1n64x5 FILLER_328_790 ();
 b15zdnd11an1n64x5 FILLER_328_854 ();
 b15zdnd11an1n64x5 FILLER_328_918 ();
 b15zdnd11an1n64x5 FILLER_328_982 ();
 b15zdnd11an1n64x5 FILLER_328_1046 ();
 b15zdnd11an1n64x5 FILLER_328_1110 ();
 b15zdnd11an1n64x5 FILLER_328_1174 ();
 b15zdnd11an1n64x5 FILLER_328_1238 ();
 b15zdnd11an1n64x5 FILLER_328_1302 ();
 b15zdnd11an1n64x5 FILLER_328_1366 ();
 b15zdnd11an1n64x5 FILLER_328_1430 ();
 b15zdnd11an1n64x5 FILLER_328_1494 ();
 b15zdnd11an1n64x5 FILLER_328_1558 ();
 b15zdnd11an1n64x5 FILLER_328_1622 ();
 b15zdnd11an1n64x5 FILLER_328_1686 ();
 b15zdnd11an1n64x5 FILLER_328_1750 ();
 b15zdnd11an1n64x5 FILLER_328_1814 ();
 b15zdnd11an1n64x5 FILLER_328_1878 ();
 b15zdnd11an1n64x5 FILLER_328_1942 ();
 b15zdnd11an1n64x5 FILLER_328_2006 ();
 b15zdnd11an1n64x5 FILLER_328_2070 ();
 b15zdnd11an1n16x5 FILLER_328_2134 ();
 b15zdnd11an1n04x5 FILLER_328_2150 ();
 b15zdnd11an1n64x5 FILLER_328_2162 ();
 b15zdnd11an1n32x5 FILLER_328_2226 ();
 b15zdnd11an1n16x5 FILLER_328_2258 ();
 b15zdnd00an1n02x5 FILLER_328_2274 ();
 b15zdnd11an1n64x5 FILLER_329_0 ();
 b15zdnd11an1n64x5 FILLER_329_64 ();
 b15zdnd11an1n64x5 FILLER_329_128 ();
 b15zdnd11an1n64x5 FILLER_329_192 ();
 b15zdnd11an1n64x5 FILLER_329_256 ();
 b15zdnd11an1n64x5 FILLER_329_320 ();
 b15zdnd11an1n64x5 FILLER_329_384 ();
 b15zdnd11an1n64x5 FILLER_329_448 ();
 b15zdnd11an1n64x5 FILLER_329_512 ();
 b15zdnd11an1n64x5 FILLER_329_576 ();
 b15zdnd11an1n64x5 FILLER_329_640 ();
 b15zdnd11an1n64x5 FILLER_329_704 ();
 b15zdnd11an1n64x5 FILLER_329_768 ();
 b15zdnd11an1n64x5 FILLER_329_832 ();
 b15zdnd11an1n64x5 FILLER_329_896 ();
 b15zdnd11an1n64x5 FILLER_329_960 ();
 b15zdnd11an1n64x5 FILLER_329_1024 ();
 b15zdnd11an1n64x5 FILLER_329_1088 ();
 b15zdnd11an1n64x5 FILLER_329_1152 ();
 b15zdnd11an1n64x5 FILLER_329_1216 ();
 b15zdnd11an1n64x5 FILLER_329_1280 ();
 b15zdnd11an1n64x5 FILLER_329_1344 ();
 b15zdnd11an1n64x5 FILLER_329_1408 ();
 b15zdnd11an1n64x5 FILLER_329_1472 ();
 b15zdnd11an1n64x5 FILLER_329_1536 ();
 b15zdnd11an1n64x5 FILLER_329_1600 ();
 b15zdnd11an1n64x5 FILLER_329_1664 ();
 b15zdnd11an1n64x5 FILLER_329_1728 ();
 b15zdnd11an1n64x5 FILLER_329_1792 ();
 b15zdnd11an1n64x5 FILLER_329_1856 ();
 b15zdnd11an1n64x5 FILLER_329_1920 ();
 b15zdnd11an1n64x5 FILLER_329_1984 ();
 b15zdnd11an1n64x5 FILLER_329_2048 ();
 b15zdnd11an1n64x5 FILLER_329_2112 ();
 b15zdnd11an1n64x5 FILLER_329_2176 ();
 b15zdnd11an1n32x5 FILLER_329_2240 ();
 b15zdnd11an1n08x5 FILLER_329_2272 ();
 b15zdnd11an1n04x5 FILLER_329_2280 ();
 b15zdnd11an1n64x5 FILLER_330_8 ();
 b15zdnd11an1n64x5 FILLER_330_72 ();
 b15zdnd11an1n64x5 FILLER_330_136 ();
 b15zdnd11an1n64x5 FILLER_330_200 ();
 b15zdnd11an1n64x5 FILLER_330_264 ();
 b15zdnd11an1n64x5 FILLER_330_328 ();
 b15zdnd11an1n64x5 FILLER_330_392 ();
 b15zdnd11an1n64x5 FILLER_330_456 ();
 b15zdnd11an1n64x5 FILLER_330_520 ();
 b15zdnd11an1n64x5 FILLER_330_584 ();
 b15zdnd11an1n64x5 FILLER_330_648 ();
 b15zdnd11an1n04x5 FILLER_330_712 ();
 b15zdnd00an1n02x5 FILLER_330_716 ();
 b15zdnd11an1n64x5 FILLER_330_726 ();
 b15zdnd11an1n64x5 FILLER_330_790 ();
 b15zdnd11an1n64x5 FILLER_330_854 ();
 b15zdnd11an1n64x5 FILLER_330_918 ();
 b15zdnd11an1n64x5 FILLER_330_982 ();
 b15zdnd11an1n64x5 FILLER_330_1046 ();
 b15zdnd11an1n64x5 FILLER_330_1110 ();
 b15zdnd11an1n64x5 FILLER_330_1174 ();
 b15zdnd11an1n64x5 FILLER_330_1238 ();
 b15zdnd11an1n64x5 FILLER_330_1302 ();
 b15zdnd11an1n64x5 FILLER_330_1366 ();
 b15zdnd11an1n64x5 FILLER_330_1430 ();
 b15zdnd11an1n64x5 FILLER_330_1494 ();
 b15zdnd11an1n64x5 FILLER_330_1558 ();
 b15zdnd11an1n64x5 FILLER_330_1622 ();
 b15zdnd11an1n64x5 FILLER_330_1686 ();
 b15zdnd11an1n64x5 FILLER_330_1750 ();
 b15zdnd11an1n64x5 FILLER_330_1814 ();
 b15zdnd11an1n64x5 FILLER_330_1878 ();
 b15zdnd11an1n64x5 FILLER_330_1942 ();
 b15zdnd11an1n64x5 FILLER_330_2006 ();
 b15zdnd11an1n64x5 FILLER_330_2070 ();
 b15zdnd11an1n16x5 FILLER_330_2134 ();
 b15zdnd11an1n04x5 FILLER_330_2150 ();
 b15zdnd11an1n64x5 FILLER_330_2162 ();
 b15zdnd11an1n32x5 FILLER_330_2226 ();
 b15zdnd11an1n16x5 FILLER_330_2258 ();
 b15zdnd00an1n02x5 FILLER_330_2274 ();
 b15zdnd11an1n64x5 FILLER_331_0 ();
 b15zdnd11an1n64x5 FILLER_331_64 ();
 b15zdnd11an1n64x5 FILLER_331_128 ();
 b15zdnd11an1n64x5 FILLER_331_192 ();
 b15zdnd11an1n64x5 FILLER_331_256 ();
 b15zdnd11an1n64x5 FILLER_331_320 ();
 b15zdnd11an1n64x5 FILLER_331_384 ();
 b15zdnd11an1n64x5 FILLER_331_448 ();
 b15zdnd11an1n64x5 FILLER_331_512 ();
 b15zdnd11an1n64x5 FILLER_331_576 ();
 b15zdnd11an1n64x5 FILLER_331_640 ();
 b15zdnd11an1n64x5 FILLER_331_704 ();
 b15zdnd11an1n64x5 FILLER_331_768 ();
 b15zdnd11an1n64x5 FILLER_331_832 ();
 b15zdnd11an1n64x5 FILLER_331_896 ();
 b15zdnd11an1n64x5 FILLER_331_960 ();
 b15zdnd11an1n64x5 FILLER_331_1024 ();
 b15zdnd11an1n64x5 FILLER_331_1088 ();
 b15zdnd11an1n64x5 FILLER_331_1152 ();
 b15zdnd11an1n64x5 FILLER_331_1216 ();
 b15zdnd11an1n64x5 FILLER_331_1280 ();
 b15zdnd11an1n64x5 FILLER_331_1344 ();
 b15zdnd11an1n64x5 FILLER_331_1408 ();
 b15zdnd11an1n64x5 FILLER_331_1472 ();
 b15zdnd11an1n64x5 FILLER_331_1536 ();
 b15zdnd11an1n64x5 FILLER_331_1600 ();
 b15zdnd11an1n64x5 FILLER_331_1664 ();
 b15zdnd11an1n64x5 FILLER_331_1728 ();
 b15zdnd11an1n64x5 FILLER_331_1792 ();
 b15zdnd11an1n64x5 FILLER_331_1856 ();
 b15zdnd11an1n64x5 FILLER_331_1920 ();
 b15zdnd11an1n64x5 FILLER_331_1984 ();
 b15zdnd11an1n64x5 FILLER_331_2048 ();
 b15zdnd11an1n64x5 FILLER_331_2112 ();
 b15zdnd11an1n64x5 FILLER_331_2176 ();
 b15zdnd11an1n32x5 FILLER_331_2240 ();
 b15zdnd11an1n08x5 FILLER_331_2272 ();
 b15zdnd11an1n04x5 FILLER_331_2280 ();
 b15zdnd11an1n64x5 FILLER_332_8 ();
 b15zdnd11an1n64x5 FILLER_332_72 ();
 b15zdnd11an1n64x5 FILLER_332_136 ();
 b15zdnd11an1n64x5 FILLER_332_200 ();
 b15zdnd11an1n64x5 FILLER_332_264 ();
 b15zdnd11an1n64x5 FILLER_332_328 ();
 b15zdnd11an1n64x5 FILLER_332_392 ();
 b15zdnd11an1n64x5 FILLER_332_456 ();
 b15zdnd11an1n64x5 FILLER_332_520 ();
 b15zdnd11an1n64x5 FILLER_332_584 ();
 b15zdnd11an1n64x5 FILLER_332_648 ();
 b15zdnd11an1n04x5 FILLER_332_712 ();
 b15zdnd00an1n02x5 FILLER_332_716 ();
 b15zdnd11an1n64x5 FILLER_332_726 ();
 b15zdnd11an1n64x5 FILLER_332_790 ();
 b15zdnd11an1n64x5 FILLER_332_854 ();
 b15zdnd11an1n64x5 FILLER_332_918 ();
 b15zdnd11an1n64x5 FILLER_332_982 ();
 b15zdnd11an1n64x5 FILLER_332_1046 ();
 b15zdnd11an1n64x5 FILLER_332_1110 ();
 b15zdnd11an1n64x5 FILLER_332_1174 ();
 b15zdnd11an1n64x5 FILLER_332_1238 ();
 b15zdnd11an1n64x5 FILLER_332_1302 ();
 b15zdnd11an1n64x5 FILLER_332_1366 ();
 b15zdnd11an1n64x5 FILLER_332_1430 ();
 b15zdnd11an1n64x5 FILLER_332_1494 ();
 b15zdnd11an1n64x5 FILLER_332_1558 ();
 b15zdnd11an1n64x5 FILLER_332_1622 ();
 b15zdnd11an1n64x5 FILLER_332_1686 ();
 b15zdnd11an1n64x5 FILLER_332_1750 ();
 b15zdnd11an1n64x5 FILLER_332_1814 ();
 b15zdnd11an1n64x5 FILLER_332_1878 ();
 b15zdnd11an1n64x5 FILLER_332_1942 ();
 b15zdnd11an1n64x5 FILLER_332_2006 ();
 b15zdnd11an1n64x5 FILLER_332_2070 ();
 b15zdnd11an1n16x5 FILLER_332_2134 ();
 b15zdnd11an1n04x5 FILLER_332_2150 ();
 b15zdnd11an1n64x5 FILLER_332_2162 ();
 b15zdnd11an1n32x5 FILLER_332_2226 ();
 b15zdnd11an1n16x5 FILLER_332_2258 ();
 b15zdnd00an1n02x5 FILLER_332_2274 ();
 b15zdnd11an1n64x5 FILLER_333_0 ();
 b15zdnd11an1n64x5 FILLER_333_64 ();
 b15zdnd11an1n64x5 FILLER_333_128 ();
 b15zdnd11an1n64x5 FILLER_333_192 ();
 b15zdnd11an1n64x5 FILLER_333_256 ();
 b15zdnd11an1n64x5 FILLER_333_320 ();
 b15zdnd11an1n64x5 FILLER_333_384 ();
 b15zdnd11an1n64x5 FILLER_333_448 ();
 b15zdnd11an1n64x5 FILLER_333_512 ();
 b15zdnd11an1n64x5 FILLER_333_576 ();
 b15zdnd11an1n64x5 FILLER_333_640 ();
 b15zdnd11an1n64x5 FILLER_333_704 ();
 b15zdnd11an1n64x5 FILLER_333_768 ();
 b15zdnd11an1n64x5 FILLER_333_832 ();
 b15zdnd11an1n64x5 FILLER_333_896 ();
 b15zdnd11an1n64x5 FILLER_333_960 ();
 b15zdnd11an1n64x5 FILLER_333_1024 ();
 b15zdnd11an1n64x5 FILLER_333_1088 ();
 b15zdnd11an1n64x5 FILLER_333_1152 ();
 b15zdnd11an1n64x5 FILLER_333_1216 ();
 b15zdnd11an1n64x5 FILLER_333_1280 ();
 b15zdnd11an1n64x5 FILLER_333_1344 ();
 b15zdnd11an1n64x5 FILLER_333_1408 ();
 b15zdnd11an1n64x5 FILLER_333_1472 ();
 b15zdnd11an1n64x5 FILLER_333_1536 ();
 b15zdnd11an1n64x5 FILLER_333_1600 ();
 b15zdnd11an1n64x5 FILLER_333_1664 ();
 b15zdnd11an1n64x5 FILLER_333_1728 ();
 b15zdnd11an1n64x5 FILLER_333_1792 ();
 b15zdnd11an1n64x5 FILLER_333_1856 ();
 b15zdnd11an1n64x5 FILLER_333_1920 ();
 b15zdnd11an1n64x5 FILLER_333_1984 ();
 b15zdnd11an1n64x5 FILLER_333_2048 ();
 b15zdnd11an1n64x5 FILLER_333_2112 ();
 b15zdnd11an1n64x5 FILLER_333_2176 ();
 b15zdnd11an1n32x5 FILLER_333_2240 ();
 b15zdnd11an1n08x5 FILLER_333_2272 ();
 b15zdnd11an1n04x5 FILLER_333_2280 ();
 b15zdnd11an1n64x5 FILLER_334_8 ();
 b15zdnd11an1n64x5 FILLER_334_72 ();
 b15zdnd11an1n64x5 FILLER_334_136 ();
 b15zdnd11an1n64x5 FILLER_334_200 ();
 b15zdnd11an1n64x5 FILLER_334_264 ();
 b15zdnd11an1n64x5 FILLER_334_328 ();
 b15zdnd11an1n64x5 FILLER_334_392 ();
 b15zdnd11an1n64x5 FILLER_334_456 ();
 b15zdnd11an1n64x5 FILLER_334_520 ();
 b15zdnd11an1n64x5 FILLER_334_584 ();
 b15zdnd11an1n64x5 FILLER_334_648 ();
 b15zdnd11an1n04x5 FILLER_334_712 ();
 b15zdnd00an1n02x5 FILLER_334_716 ();
 b15zdnd11an1n64x5 FILLER_334_726 ();
 b15zdnd11an1n64x5 FILLER_334_790 ();
 b15zdnd11an1n64x5 FILLER_334_854 ();
 b15zdnd11an1n64x5 FILLER_334_918 ();
 b15zdnd11an1n64x5 FILLER_334_982 ();
 b15zdnd11an1n64x5 FILLER_334_1046 ();
 b15zdnd11an1n64x5 FILLER_334_1110 ();
 b15zdnd11an1n64x5 FILLER_334_1174 ();
 b15zdnd11an1n64x5 FILLER_334_1238 ();
 b15zdnd11an1n64x5 FILLER_334_1302 ();
 b15zdnd11an1n64x5 FILLER_334_1366 ();
 b15zdnd11an1n64x5 FILLER_334_1430 ();
 b15zdnd11an1n64x5 FILLER_334_1494 ();
 b15zdnd11an1n64x5 FILLER_334_1558 ();
 b15zdnd11an1n64x5 FILLER_334_1622 ();
 b15zdnd11an1n64x5 FILLER_334_1686 ();
 b15zdnd11an1n64x5 FILLER_334_1750 ();
 b15zdnd11an1n64x5 FILLER_334_1814 ();
 b15zdnd11an1n64x5 FILLER_334_1878 ();
 b15zdnd11an1n64x5 FILLER_334_1942 ();
 b15zdnd11an1n64x5 FILLER_334_2006 ();
 b15zdnd11an1n64x5 FILLER_334_2070 ();
 b15zdnd11an1n16x5 FILLER_334_2134 ();
 b15zdnd11an1n04x5 FILLER_334_2150 ();
 b15zdnd11an1n64x5 FILLER_334_2162 ();
 b15zdnd11an1n32x5 FILLER_334_2226 ();
 b15zdnd11an1n16x5 FILLER_334_2258 ();
 b15zdnd00an1n02x5 FILLER_334_2274 ();
 b15zdnd11an1n64x5 FILLER_335_0 ();
 b15zdnd11an1n64x5 FILLER_335_64 ();
 b15zdnd11an1n64x5 FILLER_335_128 ();
 b15zdnd11an1n64x5 FILLER_335_192 ();
 b15zdnd11an1n64x5 FILLER_335_256 ();
 b15zdnd11an1n64x5 FILLER_335_320 ();
 b15zdnd11an1n64x5 FILLER_335_384 ();
 b15zdnd11an1n64x5 FILLER_335_448 ();
 b15zdnd11an1n64x5 FILLER_335_512 ();
 b15zdnd11an1n64x5 FILLER_335_576 ();
 b15zdnd11an1n64x5 FILLER_335_640 ();
 b15zdnd11an1n64x5 FILLER_335_704 ();
 b15zdnd11an1n64x5 FILLER_335_768 ();
 b15zdnd11an1n64x5 FILLER_335_832 ();
 b15zdnd11an1n64x5 FILLER_335_896 ();
 b15zdnd11an1n64x5 FILLER_335_960 ();
 b15zdnd11an1n64x5 FILLER_335_1024 ();
 b15zdnd11an1n64x5 FILLER_335_1088 ();
 b15zdnd11an1n64x5 FILLER_335_1152 ();
 b15zdnd11an1n64x5 FILLER_335_1216 ();
 b15zdnd11an1n64x5 FILLER_335_1280 ();
 b15zdnd11an1n64x5 FILLER_335_1344 ();
 b15zdnd11an1n64x5 FILLER_335_1408 ();
 b15zdnd11an1n64x5 FILLER_335_1472 ();
 b15zdnd11an1n64x5 FILLER_335_1536 ();
 b15zdnd11an1n64x5 FILLER_335_1600 ();
 b15zdnd11an1n64x5 FILLER_335_1664 ();
 b15zdnd11an1n64x5 FILLER_335_1728 ();
 b15zdnd11an1n64x5 FILLER_335_1792 ();
 b15zdnd11an1n64x5 FILLER_335_1856 ();
 b15zdnd11an1n64x5 FILLER_335_1920 ();
 b15zdnd11an1n64x5 FILLER_335_1984 ();
 b15zdnd11an1n64x5 FILLER_335_2048 ();
 b15zdnd11an1n64x5 FILLER_335_2112 ();
 b15zdnd11an1n64x5 FILLER_335_2176 ();
 b15zdnd11an1n32x5 FILLER_335_2240 ();
 b15zdnd11an1n08x5 FILLER_335_2272 ();
 b15zdnd11an1n04x5 FILLER_335_2280 ();
 b15zdnd11an1n64x5 FILLER_336_8 ();
 b15zdnd11an1n64x5 FILLER_336_72 ();
 b15zdnd11an1n64x5 FILLER_336_136 ();
 b15zdnd11an1n64x5 FILLER_336_200 ();
 b15zdnd11an1n64x5 FILLER_336_264 ();
 b15zdnd11an1n64x5 FILLER_336_328 ();
 b15zdnd11an1n64x5 FILLER_336_392 ();
 b15zdnd11an1n64x5 FILLER_336_456 ();
 b15zdnd11an1n64x5 FILLER_336_520 ();
 b15zdnd11an1n64x5 FILLER_336_584 ();
 b15zdnd11an1n64x5 FILLER_336_648 ();
 b15zdnd11an1n04x5 FILLER_336_712 ();
 b15zdnd00an1n02x5 FILLER_336_716 ();
 b15zdnd11an1n64x5 FILLER_336_726 ();
 b15zdnd11an1n64x5 FILLER_336_790 ();
 b15zdnd11an1n64x5 FILLER_336_854 ();
 b15zdnd11an1n64x5 FILLER_336_918 ();
 b15zdnd11an1n64x5 FILLER_336_982 ();
 b15zdnd11an1n64x5 FILLER_336_1046 ();
 b15zdnd11an1n64x5 FILLER_336_1110 ();
 b15zdnd11an1n64x5 FILLER_336_1174 ();
 b15zdnd11an1n64x5 FILLER_336_1238 ();
 b15zdnd11an1n64x5 FILLER_336_1302 ();
 b15zdnd11an1n64x5 FILLER_336_1366 ();
 b15zdnd11an1n64x5 FILLER_336_1430 ();
 b15zdnd11an1n64x5 FILLER_336_1494 ();
 b15zdnd11an1n64x5 FILLER_336_1558 ();
 b15zdnd11an1n64x5 FILLER_336_1622 ();
 b15zdnd11an1n64x5 FILLER_336_1686 ();
 b15zdnd11an1n64x5 FILLER_336_1750 ();
 b15zdnd11an1n64x5 FILLER_336_1814 ();
 b15zdnd11an1n64x5 FILLER_336_1878 ();
 b15zdnd11an1n64x5 FILLER_336_1942 ();
 b15zdnd11an1n64x5 FILLER_336_2006 ();
 b15zdnd11an1n64x5 FILLER_336_2070 ();
 b15zdnd11an1n16x5 FILLER_336_2134 ();
 b15zdnd11an1n04x5 FILLER_336_2150 ();
 b15zdnd11an1n64x5 FILLER_336_2162 ();
 b15zdnd11an1n32x5 FILLER_336_2226 ();
 b15zdnd11an1n16x5 FILLER_336_2258 ();
 b15zdnd00an1n02x5 FILLER_336_2274 ();
 b15zdnd11an1n64x5 FILLER_337_0 ();
 b15zdnd11an1n64x5 FILLER_337_64 ();
 b15zdnd11an1n64x5 FILLER_337_128 ();
 b15zdnd11an1n64x5 FILLER_337_192 ();
 b15zdnd11an1n64x5 FILLER_337_256 ();
 b15zdnd11an1n64x5 FILLER_337_320 ();
 b15zdnd11an1n64x5 FILLER_337_384 ();
 b15zdnd11an1n64x5 FILLER_337_448 ();
 b15zdnd11an1n64x5 FILLER_337_512 ();
 b15zdnd11an1n64x5 FILLER_337_576 ();
 b15zdnd11an1n64x5 FILLER_337_640 ();
 b15zdnd11an1n64x5 FILLER_337_704 ();
 b15zdnd11an1n64x5 FILLER_337_768 ();
 b15zdnd11an1n64x5 FILLER_337_832 ();
 b15zdnd11an1n64x5 FILLER_337_896 ();
 b15zdnd11an1n64x5 FILLER_337_960 ();
 b15zdnd11an1n64x5 FILLER_337_1024 ();
 b15zdnd11an1n64x5 FILLER_337_1088 ();
 b15zdnd11an1n64x5 FILLER_337_1152 ();
 b15zdnd11an1n64x5 FILLER_337_1216 ();
 b15zdnd11an1n64x5 FILLER_337_1280 ();
 b15zdnd11an1n64x5 FILLER_337_1344 ();
 b15zdnd11an1n64x5 FILLER_337_1408 ();
 b15zdnd11an1n64x5 FILLER_337_1472 ();
 b15zdnd11an1n64x5 FILLER_337_1536 ();
 b15zdnd11an1n64x5 FILLER_337_1600 ();
 b15zdnd11an1n64x5 FILLER_337_1664 ();
 b15zdnd11an1n64x5 FILLER_337_1728 ();
 b15zdnd11an1n64x5 FILLER_337_1792 ();
 b15zdnd11an1n64x5 FILLER_337_1856 ();
 b15zdnd11an1n64x5 FILLER_337_1920 ();
 b15zdnd11an1n64x5 FILLER_337_1984 ();
 b15zdnd11an1n64x5 FILLER_337_2048 ();
 b15zdnd11an1n64x5 FILLER_337_2112 ();
 b15zdnd11an1n64x5 FILLER_337_2176 ();
 b15zdnd11an1n32x5 FILLER_337_2240 ();
 b15zdnd11an1n08x5 FILLER_337_2272 ();
 b15zdnd11an1n04x5 FILLER_337_2280 ();
 b15zdnd11an1n64x5 FILLER_338_8 ();
 b15zdnd11an1n64x5 FILLER_338_72 ();
 b15zdnd11an1n64x5 FILLER_338_136 ();
 b15zdnd11an1n64x5 FILLER_338_200 ();
 b15zdnd11an1n64x5 FILLER_338_264 ();
 b15zdnd11an1n64x5 FILLER_338_328 ();
 b15zdnd11an1n64x5 FILLER_338_392 ();
 b15zdnd11an1n64x5 FILLER_338_456 ();
 b15zdnd11an1n64x5 FILLER_338_520 ();
 b15zdnd11an1n64x5 FILLER_338_584 ();
 b15zdnd11an1n64x5 FILLER_338_648 ();
 b15zdnd11an1n04x5 FILLER_338_712 ();
 b15zdnd00an1n02x5 FILLER_338_716 ();
 b15zdnd11an1n64x5 FILLER_338_726 ();
 b15zdnd11an1n64x5 FILLER_338_790 ();
 b15zdnd11an1n64x5 FILLER_338_854 ();
 b15zdnd11an1n64x5 FILLER_338_918 ();
 b15zdnd11an1n64x5 FILLER_338_982 ();
 b15zdnd11an1n64x5 FILLER_338_1046 ();
 b15zdnd11an1n64x5 FILLER_338_1110 ();
 b15zdnd11an1n64x5 FILLER_338_1174 ();
 b15zdnd11an1n64x5 FILLER_338_1238 ();
 b15zdnd11an1n64x5 FILLER_338_1302 ();
 b15zdnd11an1n64x5 FILLER_338_1366 ();
 b15zdnd11an1n64x5 FILLER_338_1430 ();
 b15zdnd11an1n64x5 FILLER_338_1494 ();
 b15zdnd11an1n64x5 FILLER_338_1558 ();
 b15zdnd11an1n64x5 FILLER_338_1622 ();
 b15zdnd11an1n64x5 FILLER_338_1686 ();
 b15zdnd11an1n64x5 FILLER_338_1750 ();
 b15zdnd11an1n64x5 FILLER_338_1814 ();
 b15zdnd11an1n64x5 FILLER_338_1878 ();
 b15zdnd11an1n64x5 FILLER_338_1942 ();
 b15zdnd11an1n64x5 FILLER_338_2006 ();
 b15zdnd11an1n64x5 FILLER_338_2070 ();
 b15zdnd11an1n16x5 FILLER_338_2134 ();
 b15zdnd11an1n04x5 FILLER_338_2150 ();
 b15zdnd11an1n64x5 FILLER_338_2162 ();
 b15zdnd11an1n32x5 FILLER_338_2226 ();
 b15zdnd11an1n16x5 FILLER_338_2258 ();
 b15zdnd00an1n02x5 FILLER_338_2274 ();
 b15zdnd11an1n64x5 FILLER_339_0 ();
 b15zdnd11an1n64x5 FILLER_339_64 ();
 b15zdnd11an1n64x5 FILLER_339_128 ();
 b15zdnd11an1n64x5 FILLER_339_192 ();
 b15zdnd11an1n64x5 FILLER_339_256 ();
 b15zdnd11an1n64x5 FILLER_339_320 ();
 b15zdnd11an1n64x5 FILLER_339_384 ();
 b15zdnd11an1n64x5 FILLER_339_448 ();
 b15zdnd11an1n64x5 FILLER_339_512 ();
 b15zdnd11an1n64x5 FILLER_339_576 ();
 b15zdnd11an1n64x5 FILLER_339_640 ();
 b15zdnd11an1n64x5 FILLER_339_704 ();
 b15zdnd11an1n64x5 FILLER_339_768 ();
 b15zdnd11an1n64x5 FILLER_339_832 ();
 b15zdnd11an1n64x5 FILLER_339_896 ();
 b15zdnd11an1n64x5 FILLER_339_960 ();
 b15zdnd11an1n64x5 FILLER_339_1024 ();
 b15zdnd11an1n64x5 FILLER_339_1088 ();
 b15zdnd11an1n64x5 FILLER_339_1152 ();
 b15zdnd11an1n64x5 FILLER_339_1216 ();
 b15zdnd11an1n64x5 FILLER_339_1280 ();
 b15zdnd11an1n64x5 FILLER_339_1344 ();
 b15zdnd11an1n64x5 FILLER_339_1408 ();
 b15zdnd11an1n64x5 FILLER_339_1472 ();
 b15zdnd11an1n64x5 FILLER_339_1536 ();
 b15zdnd11an1n64x5 FILLER_339_1600 ();
 b15zdnd11an1n64x5 FILLER_339_1664 ();
 b15zdnd11an1n64x5 FILLER_339_1728 ();
 b15zdnd11an1n64x5 FILLER_339_1792 ();
 b15zdnd11an1n64x5 FILLER_339_1856 ();
 b15zdnd11an1n64x5 FILLER_339_1920 ();
 b15zdnd11an1n64x5 FILLER_339_1984 ();
 b15zdnd11an1n64x5 FILLER_339_2048 ();
 b15zdnd11an1n64x5 FILLER_339_2112 ();
 b15zdnd11an1n64x5 FILLER_339_2176 ();
 b15zdnd11an1n32x5 FILLER_339_2240 ();
 b15zdnd11an1n08x5 FILLER_339_2272 ();
 b15zdnd11an1n04x5 FILLER_339_2280 ();
 b15zdnd11an1n64x5 FILLER_340_8 ();
 b15zdnd11an1n64x5 FILLER_340_72 ();
 b15zdnd11an1n64x5 FILLER_340_136 ();
 b15zdnd11an1n64x5 FILLER_340_200 ();
 b15zdnd11an1n64x5 FILLER_340_264 ();
 b15zdnd11an1n64x5 FILLER_340_328 ();
 b15zdnd11an1n64x5 FILLER_340_392 ();
 b15zdnd11an1n64x5 FILLER_340_456 ();
 b15zdnd11an1n64x5 FILLER_340_520 ();
 b15zdnd11an1n64x5 FILLER_340_584 ();
 b15zdnd11an1n64x5 FILLER_340_648 ();
 b15zdnd11an1n04x5 FILLER_340_712 ();
 b15zdnd00an1n02x5 FILLER_340_716 ();
 b15zdnd11an1n64x5 FILLER_340_726 ();
 b15zdnd11an1n64x5 FILLER_340_790 ();
 b15zdnd11an1n64x5 FILLER_340_854 ();
 b15zdnd11an1n64x5 FILLER_340_918 ();
 b15zdnd11an1n64x5 FILLER_340_982 ();
 b15zdnd11an1n64x5 FILLER_340_1046 ();
 b15zdnd11an1n64x5 FILLER_340_1110 ();
 b15zdnd11an1n64x5 FILLER_340_1174 ();
 b15zdnd11an1n64x5 FILLER_340_1238 ();
 b15zdnd11an1n64x5 FILLER_340_1302 ();
 b15zdnd11an1n64x5 FILLER_340_1366 ();
 b15zdnd11an1n64x5 FILLER_340_1430 ();
 b15zdnd11an1n64x5 FILLER_340_1494 ();
 b15zdnd11an1n64x5 FILLER_340_1558 ();
 b15zdnd11an1n64x5 FILLER_340_1622 ();
 b15zdnd11an1n64x5 FILLER_340_1686 ();
 b15zdnd11an1n64x5 FILLER_340_1750 ();
 b15zdnd11an1n64x5 FILLER_340_1814 ();
 b15zdnd11an1n64x5 FILLER_340_1878 ();
 b15zdnd11an1n64x5 FILLER_340_1942 ();
 b15zdnd11an1n64x5 FILLER_340_2006 ();
 b15zdnd11an1n64x5 FILLER_340_2070 ();
 b15zdnd11an1n16x5 FILLER_340_2134 ();
 b15zdnd11an1n04x5 FILLER_340_2150 ();
 b15zdnd11an1n64x5 FILLER_340_2162 ();
 b15zdnd11an1n32x5 FILLER_340_2226 ();
 b15zdnd11an1n16x5 FILLER_340_2258 ();
 b15zdnd00an1n02x5 FILLER_340_2274 ();
 b15zdnd11an1n64x5 FILLER_341_0 ();
 b15zdnd11an1n64x5 FILLER_341_64 ();
 b15zdnd11an1n64x5 FILLER_341_128 ();
 b15zdnd11an1n64x5 FILLER_341_192 ();
 b15zdnd11an1n64x5 FILLER_341_256 ();
 b15zdnd11an1n64x5 FILLER_341_320 ();
 b15zdnd11an1n64x5 FILLER_341_384 ();
 b15zdnd11an1n64x5 FILLER_341_448 ();
 b15zdnd11an1n64x5 FILLER_341_512 ();
 b15zdnd11an1n64x5 FILLER_341_576 ();
 b15zdnd11an1n64x5 FILLER_341_640 ();
 b15zdnd11an1n64x5 FILLER_341_704 ();
 b15zdnd11an1n64x5 FILLER_341_768 ();
 b15zdnd11an1n64x5 FILLER_341_832 ();
 b15zdnd11an1n64x5 FILLER_341_896 ();
 b15zdnd11an1n64x5 FILLER_341_960 ();
 b15zdnd11an1n64x5 FILLER_341_1024 ();
 b15zdnd11an1n64x5 FILLER_341_1088 ();
 b15zdnd11an1n64x5 FILLER_341_1152 ();
 b15zdnd11an1n64x5 FILLER_341_1216 ();
 b15zdnd11an1n64x5 FILLER_341_1280 ();
 b15zdnd11an1n64x5 FILLER_341_1344 ();
 b15zdnd11an1n64x5 FILLER_341_1408 ();
 b15zdnd11an1n64x5 FILLER_341_1472 ();
 b15zdnd11an1n64x5 FILLER_341_1536 ();
 b15zdnd11an1n64x5 FILLER_341_1600 ();
 b15zdnd11an1n64x5 FILLER_341_1664 ();
 b15zdnd11an1n64x5 FILLER_341_1728 ();
 b15zdnd11an1n64x5 FILLER_341_1792 ();
 b15zdnd11an1n64x5 FILLER_341_1856 ();
 b15zdnd11an1n64x5 FILLER_341_1920 ();
 b15zdnd11an1n64x5 FILLER_341_1984 ();
 b15zdnd11an1n64x5 FILLER_341_2048 ();
 b15zdnd11an1n64x5 FILLER_341_2112 ();
 b15zdnd11an1n64x5 FILLER_341_2176 ();
 b15zdnd11an1n32x5 FILLER_341_2240 ();
 b15zdnd11an1n08x5 FILLER_341_2272 ();
 b15zdnd11an1n04x5 FILLER_341_2280 ();
 b15zdnd11an1n64x5 FILLER_342_8 ();
 b15zdnd11an1n64x5 FILLER_342_72 ();
 b15zdnd11an1n64x5 FILLER_342_136 ();
 b15zdnd11an1n64x5 FILLER_342_200 ();
 b15zdnd11an1n64x5 FILLER_342_264 ();
 b15zdnd11an1n64x5 FILLER_342_328 ();
 b15zdnd11an1n64x5 FILLER_342_392 ();
 b15zdnd11an1n64x5 FILLER_342_456 ();
 b15zdnd11an1n64x5 FILLER_342_520 ();
 b15zdnd11an1n64x5 FILLER_342_584 ();
 b15zdnd11an1n64x5 FILLER_342_648 ();
 b15zdnd11an1n04x5 FILLER_342_712 ();
 b15zdnd00an1n02x5 FILLER_342_716 ();
 b15zdnd11an1n64x5 FILLER_342_726 ();
 b15zdnd11an1n64x5 FILLER_342_790 ();
 b15zdnd11an1n64x5 FILLER_342_854 ();
 b15zdnd11an1n64x5 FILLER_342_918 ();
 b15zdnd11an1n64x5 FILLER_342_982 ();
 b15zdnd11an1n64x5 FILLER_342_1046 ();
 b15zdnd11an1n64x5 FILLER_342_1110 ();
 b15zdnd11an1n64x5 FILLER_342_1174 ();
 b15zdnd11an1n64x5 FILLER_342_1238 ();
 b15zdnd11an1n64x5 FILLER_342_1302 ();
 b15zdnd11an1n64x5 FILLER_342_1366 ();
 b15zdnd11an1n64x5 FILLER_342_1430 ();
 b15zdnd11an1n64x5 FILLER_342_1494 ();
 b15zdnd11an1n64x5 FILLER_342_1558 ();
 b15zdnd11an1n64x5 FILLER_342_1622 ();
 b15zdnd11an1n64x5 FILLER_342_1686 ();
 b15zdnd11an1n64x5 FILLER_342_1750 ();
 b15zdnd11an1n64x5 FILLER_342_1814 ();
 b15zdnd11an1n64x5 FILLER_342_1878 ();
 b15zdnd11an1n64x5 FILLER_342_1942 ();
 b15zdnd11an1n64x5 FILLER_342_2006 ();
 b15zdnd11an1n64x5 FILLER_342_2070 ();
 b15zdnd11an1n16x5 FILLER_342_2134 ();
 b15zdnd11an1n04x5 FILLER_342_2150 ();
 b15zdnd11an1n64x5 FILLER_342_2162 ();
 b15zdnd11an1n32x5 FILLER_342_2226 ();
 b15zdnd11an1n16x5 FILLER_342_2258 ();
 b15zdnd00an1n02x5 FILLER_342_2274 ();
 b15zdnd11an1n64x5 FILLER_343_0 ();
 b15zdnd11an1n64x5 FILLER_343_64 ();
 b15zdnd11an1n64x5 FILLER_343_128 ();
 b15zdnd11an1n64x5 FILLER_343_192 ();
 b15zdnd11an1n64x5 FILLER_343_256 ();
 b15zdnd11an1n64x5 FILLER_343_320 ();
 b15zdnd11an1n64x5 FILLER_343_384 ();
 b15zdnd11an1n64x5 FILLER_343_448 ();
 b15zdnd11an1n64x5 FILLER_343_512 ();
 b15zdnd11an1n64x5 FILLER_343_576 ();
 b15zdnd11an1n64x5 FILLER_343_640 ();
 b15zdnd11an1n64x5 FILLER_343_704 ();
 b15zdnd11an1n64x5 FILLER_343_768 ();
 b15zdnd11an1n64x5 FILLER_343_832 ();
 b15zdnd11an1n64x5 FILLER_343_896 ();
 b15zdnd11an1n64x5 FILLER_343_960 ();
 b15zdnd11an1n64x5 FILLER_343_1024 ();
 b15zdnd11an1n64x5 FILLER_343_1088 ();
 b15zdnd11an1n64x5 FILLER_343_1152 ();
 b15zdnd11an1n64x5 FILLER_343_1216 ();
 b15zdnd11an1n64x5 FILLER_343_1280 ();
 b15zdnd11an1n64x5 FILLER_343_1344 ();
 b15zdnd11an1n64x5 FILLER_343_1408 ();
 b15zdnd11an1n64x5 FILLER_343_1472 ();
 b15zdnd11an1n64x5 FILLER_343_1536 ();
 b15zdnd11an1n64x5 FILLER_343_1600 ();
 b15zdnd11an1n64x5 FILLER_343_1664 ();
 b15zdnd11an1n64x5 FILLER_343_1728 ();
 b15zdnd11an1n64x5 FILLER_343_1792 ();
 b15zdnd11an1n64x5 FILLER_343_1856 ();
 b15zdnd11an1n64x5 FILLER_343_1920 ();
 b15zdnd11an1n64x5 FILLER_343_1984 ();
 b15zdnd11an1n64x5 FILLER_343_2048 ();
 b15zdnd11an1n64x5 FILLER_343_2112 ();
 b15zdnd11an1n64x5 FILLER_343_2176 ();
 b15zdnd11an1n32x5 FILLER_343_2240 ();
 b15zdnd11an1n08x5 FILLER_343_2272 ();
 b15zdnd11an1n04x5 FILLER_343_2280 ();
 b15zdnd11an1n64x5 FILLER_344_8 ();
 b15zdnd11an1n64x5 FILLER_344_72 ();
 b15zdnd11an1n64x5 FILLER_344_136 ();
 b15zdnd11an1n64x5 FILLER_344_200 ();
 b15zdnd11an1n64x5 FILLER_344_264 ();
 b15zdnd11an1n64x5 FILLER_344_328 ();
 b15zdnd11an1n64x5 FILLER_344_392 ();
 b15zdnd11an1n64x5 FILLER_344_456 ();
 b15zdnd11an1n64x5 FILLER_344_520 ();
 b15zdnd11an1n64x5 FILLER_344_584 ();
 b15zdnd11an1n64x5 FILLER_344_648 ();
 b15zdnd11an1n04x5 FILLER_344_712 ();
 b15zdnd00an1n02x5 FILLER_344_716 ();
 b15zdnd11an1n64x5 FILLER_344_726 ();
 b15zdnd11an1n64x5 FILLER_344_790 ();
 b15zdnd11an1n64x5 FILLER_344_854 ();
 b15zdnd11an1n64x5 FILLER_344_918 ();
 b15zdnd11an1n64x5 FILLER_344_982 ();
 b15zdnd11an1n64x5 FILLER_344_1046 ();
 b15zdnd11an1n64x5 FILLER_344_1110 ();
 b15zdnd11an1n64x5 FILLER_344_1174 ();
 b15zdnd11an1n64x5 FILLER_344_1238 ();
 b15zdnd11an1n64x5 FILLER_344_1302 ();
 b15zdnd11an1n64x5 FILLER_344_1366 ();
 b15zdnd11an1n64x5 FILLER_344_1430 ();
 b15zdnd11an1n64x5 FILLER_344_1494 ();
 b15zdnd11an1n64x5 FILLER_344_1558 ();
 b15zdnd11an1n64x5 FILLER_344_1622 ();
 b15zdnd11an1n64x5 FILLER_344_1686 ();
 b15zdnd11an1n64x5 FILLER_344_1750 ();
 b15zdnd11an1n64x5 FILLER_344_1814 ();
 b15zdnd11an1n64x5 FILLER_344_1878 ();
 b15zdnd11an1n64x5 FILLER_344_1942 ();
 b15zdnd11an1n64x5 FILLER_344_2006 ();
 b15zdnd11an1n64x5 FILLER_344_2070 ();
 b15zdnd11an1n16x5 FILLER_344_2134 ();
 b15zdnd11an1n04x5 FILLER_344_2150 ();
 b15zdnd11an1n64x5 FILLER_344_2162 ();
 b15zdnd11an1n32x5 FILLER_344_2226 ();
 b15zdnd11an1n16x5 FILLER_344_2258 ();
 b15zdnd00an1n02x5 FILLER_344_2274 ();
 b15zdnd11an1n64x5 FILLER_345_0 ();
 b15zdnd11an1n64x5 FILLER_345_64 ();
 b15zdnd11an1n64x5 FILLER_345_128 ();
 b15zdnd11an1n64x5 FILLER_345_192 ();
 b15zdnd11an1n64x5 FILLER_345_256 ();
 b15zdnd11an1n64x5 FILLER_345_320 ();
 b15zdnd11an1n64x5 FILLER_345_384 ();
 b15zdnd11an1n64x5 FILLER_345_448 ();
 b15zdnd11an1n64x5 FILLER_345_512 ();
 b15zdnd11an1n64x5 FILLER_345_576 ();
 b15zdnd11an1n64x5 FILLER_345_640 ();
 b15zdnd11an1n64x5 FILLER_345_704 ();
 b15zdnd11an1n64x5 FILLER_345_768 ();
 b15zdnd11an1n64x5 FILLER_345_832 ();
 b15zdnd11an1n64x5 FILLER_345_896 ();
 b15zdnd11an1n64x5 FILLER_345_960 ();
 b15zdnd11an1n64x5 FILLER_345_1024 ();
 b15zdnd11an1n64x5 FILLER_345_1088 ();
 b15zdnd11an1n64x5 FILLER_345_1152 ();
 b15zdnd11an1n64x5 FILLER_345_1216 ();
 b15zdnd11an1n64x5 FILLER_345_1280 ();
 b15zdnd11an1n64x5 FILLER_345_1344 ();
 b15zdnd11an1n64x5 FILLER_345_1408 ();
 b15zdnd11an1n64x5 FILLER_345_1472 ();
 b15zdnd11an1n64x5 FILLER_345_1536 ();
 b15zdnd11an1n64x5 FILLER_345_1600 ();
 b15zdnd11an1n64x5 FILLER_345_1664 ();
 b15zdnd11an1n64x5 FILLER_345_1728 ();
 b15zdnd11an1n64x5 FILLER_345_1792 ();
 b15zdnd11an1n64x5 FILLER_345_1856 ();
 b15zdnd11an1n64x5 FILLER_345_1920 ();
 b15zdnd11an1n64x5 FILLER_345_1984 ();
 b15zdnd11an1n64x5 FILLER_345_2048 ();
 b15zdnd11an1n64x5 FILLER_345_2112 ();
 b15zdnd11an1n64x5 FILLER_345_2176 ();
 b15zdnd11an1n32x5 FILLER_345_2240 ();
 b15zdnd11an1n08x5 FILLER_345_2272 ();
 b15zdnd11an1n04x5 FILLER_345_2280 ();
 b15zdnd11an1n64x5 FILLER_346_8 ();
 b15zdnd11an1n64x5 FILLER_346_72 ();
 b15zdnd11an1n64x5 FILLER_346_136 ();
 b15zdnd11an1n64x5 FILLER_346_200 ();
 b15zdnd11an1n64x5 FILLER_346_264 ();
 b15zdnd11an1n64x5 FILLER_346_328 ();
 b15zdnd11an1n64x5 FILLER_346_392 ();
 b15zdnd11an1n64x5 FILLER_346_456 ();
 b15zdnd11an1n64x5 FILLER_346_520 ();
 b15zdnd11an1n64x5 FILLER_346_584 ();
 b15zdnd11an1n64x5 FILLER_346_648 ();
 b15zdnd11an1n04x5 FILLER_346_712 ();
 b15zdnd00an1n02x5 FILLER_346_716 ();
 b15zdnd11an1n64x5 FILLER_346_726 ();
 b15zdnd11an1n64x5 FILLER_346_790 ();
 b15zdnd11an1n64x5 FILLER_346_854 ();
 b15zdnd11an1n64x5 FILLER_346_918 ();
 b15zdnd11an1n64x5 FILLER_346_982 ();
 b15zdnd11an1n64x5 FILLER_346_1046 ();
 b15zdnd11an1n64x5 FILLER_346_1110 ();
 b15zdnd11an1n64x5 FILLER_346_1174 ();
 b15zdnd11an1n64x5 FILLER_346_1238 ();
 b15zdnd11an1n64x5 FILLER_346_1302 ();
 b15zdnd11an1n64x5 FILLER_346_1366 ();
 b15zdnd11an1n64x5 FILLER_346_1430 ();
 b15zdnd11an1n64x5 FILLER_346_1494 ();
 b15zdnd11an1n64x5 FILLER_346_1558 ();
 b15zdnd11an1n64x5 FILLER_346_1622 ();
 b15zdnd11an1n64x5 FILLER_346_1686 ();
 b15zdnd11an1n64x5 FILLER_346_1750 ();
 b15zdnd11an1n64x5 FILLER_346_1814 ();
 b15zdnd11an1n64x5 FILLER_346_1878 ();
 b15zdnd11an1n64x5 FILLER_346_1942 ();
 b15zdnd11an1n64x5 FILLER_346_2006 ();
 b15zdnd11an1n64x5 FILLER_346_2070 ();
 b15zdnd11an1n16x5 FILLER_346_2134 ();
 b15zdnd11an1n04x5 FILLER_346_2150 ();
 b15zdnd11an1n64x5 FILLER_346_2162 ();
 b15zdnd11an1n32x5 FILLER_346_2226 ();
 b15zdnd11an1n16x5 FILLER_346_2258 ();
 b15zdnd00an1n02x5 FILLER_346_2274 ();
 b15zdnd11an1n64x5 FILLER_347_0 ();
 b15zdnd11an1n64x5 FILLER_347_64 ();
 b15zdnd11an1n64x5 FILLER_347_128 ();
 b15zdnd11an1n64x5 FILLER_347_192 ();
 b15zdnd11an1n64x5 FILLER_347_256 ();
 b15zdnd11an1n64x5 FILLER_347_320 ();
 b15zdnd11an1n64x5 FILLER_347_384 ();
 b15zdnd11an1n64x5 FILLER_347_448 ();
 b15zdnd11an1n64x5 FILLER_347_512 ();
 b15zdnd11an1n64x5 FILLER_347_576 ();
 b15zdnd11an1n64x5 FILLER_347_640 ();
 b15zdnd11an1n64x5 FILLER_347_704 ();
 b15zdnd11an1n64x5 FILLER_347_768 ();
 b15zdnd11an1n64x5 FILLER_347_832 ();
 b15zdnd11an1n64x5 FILLER_347_896 ();
 b15zdnd11an1n64x5 FILLER_347_960 ();
 b15zdnd11an1n64x5 FILLER_347_1024 ();
 b15zdnd11an1n64x5 FILLER_347_1088 ();
 b15zdnd11an1n64x5 FILLER_347_1152 ();
 b15zdnd11an1n64x5 FILLER_347_1216 ();
 b15zdnd11an1n64x5 FILLER_347_1280 ();
 b15zdnd11an1n64x5 FILLER_347_1344 ();
 b15zdnd11an1n64x5 FILLER_347_1408 ();
 b15zdnd11an1n64x5 FILLER_347_1472 ();
 b15zdnd11an1n64x5 FILLER_347_1536 ();
 b15zdnd11an1n64x5 FILLER_347_1600 ();
 b15zdnd11an1n64x5 FILLER_347_1664 ();
 b15zdnd11an1n64x5 FILLER_347_1728 ();
 b15zdnd11an1n64x5 FILLER_347_1792 ();
 b15zdnd11an1n64x5 FILLER_347_1856 ();
 b15zdnd11an1n64x5 FILLER_347_1920 ();
 b15zdnd11an1n64x5 FILLER_347_1984 ();
 b15zdnd11an1n64x5 FILLER_347_2048 ();
 b15zdnd11an1n64x5 FILLER_347_2112 ();
 b15zdnd11an1n64x5 FILLER_347_2176 ();
 b15zdnd11an1n32x5 FILLER_347_2240 ();
 b15zdnd11an1n08x5 FILLER_347_2272 ();
 b15zdnd11an1n04x5 FILLER_347_2280 ();
 b15zdnd11an1n64x5 FILLER_348_8 ();
 b15zdnd11an1n64x5 FILLER_348_72 ();
 b15zdnd11an1n64x5 FILLER_348_136 ();
 b15zdnd11an1n64x5 FILLER_348_200 ();
 b15zdnd11an1n64x5 FILLER_348_264 ();
 b15zdnd11an1n64x5 FILLER_348_328 ();
 b15zdnd11an1n64x5 FILLER_348_392 ();
 b15zdnd11an1n64x5 FILLER_348_456 ();
 b15zdnd11an1n64x5 FILLER_348_520 ();
 b15zdnd11an1n64x5 FILLER_348_584 ();
 b15zdnd11an1n64x5 FILLER_348_648 ();
 b15zdnd11an1n04x5 FILLER_348_712 ();
 b15zdnd00an1n02x5 FILLER_348_716 ();
 b15zdnd11an1n64x5 FILLER_348_726 ();
 b15zdnd11an1n64x5 FILLER_348_790 ();
 b15zdnd11an1n64x5 FILLER_348_854 ();
 b15zdnd11an1n64x5 FILLER_348_918 ();
 b15zdnd11an1n64x5 FILLER_348_982 ();
 b15zdnd11an1n64x5 FILLER_348_1046 ();
 b15zdnd11an1n64x5 FILLER_348_1110 ();
 b15zdnd11an1n64x5 FILLER_348_1174 ();
 b15zdnd11an1n64x5 FILLER_348_1238 ();
 b15zdnd11an1n64x5 FILLER_348_1302 ();
 b15zdnd11an1n64x5 FILLER_348_1366 ();
 b15zdnd11an1n64x5 FILLER_348_1430 ();
 b15zdnd11an1n64x5 FILLER_348_1494 ();
 b15zdnd11an1n64x5 FILLER_348_1558 ();
 b15zdnd11an1n64x5 FILLER_348_1622 ();
 b15zdnd11an1n64x5 FILLER_348_1686 ();
 b15zdnd11an1n64x5 FILLER_348_1750 ();
 b15zdnd11an1n64x5 FILLER_348_1814 ();
 b15zdnd11an1n64x5 FILLER_348_1878 ();
 b15zdnd11an1n64x5 FILLER_348_1942 ();
 b15zdnd11an1n64x5 FILLER_348_2006 ();
 b15zdnd11an1n64x5 FILLER_348_2070 ();
 b15zdnd11an1n16x5 FILLER_348_2134 ();
 b15zdnd11an1n04x5 FILLER_348_2150 ();
 b15zdnd11an1n64x5 FILLER_348_2162 ();
 b15zdnd11an1n32x5 FILLER_348_2226 ();
 b15zdnd11an1n16x5 FILLER_348_2258 ();
 b15zdnd00an1n02x5 FILLER_348_2274 ();
 b15zdnd11an1n64x5 FILLER_349_0 ();
 b15zdnd11an1n64x5 FILLER_349_64 ();
 b15zdnd11an1n64x5 FILLER_349_128 ();
 b15zdnd11an1n64x5 FILLER_349_192 ();
 b15zdnd11an1n64x5 FILLER_349_256 ();
 b15zdnd11an1n64x5 FILLER_349_320 ();
 b15zdnd11an1n64x5 FILLER_349_384 ();
 b15zdnd11an1n64x5 FILLER_349_448 ();
 b15zdnd11an1n64x5 FILLER_349_512 ();
 b15zdnd11an1n64x5 FILLER_349_576 ();
 b15zdnd11an1n64x5 FILLER_349_640 ();
 b15zdnd11an1n64x5 FILLER_349_704 ();
 b15zdnd11an1n64x5 FILLER_349_768 ();
 b15zdnd11an1n64x5 FILLER_349_832 ();
 b15zdnd11an1n64x5 FILLER_349_896 ();
 b15zdnd11an1n64x5 FILLER_349_960 ();
 b15zdnd11an1n64x5 FILLER_349_1024 ();
 b15zdnd11an1n64x5 FILLER_349_1088 ();
 b15zdnd11an1n64x5 FILLER_349_1152 ();
 b15zdnd11an1n64x5 FILLER_349_1216 ();
 b15zdnd11an1n64x5 FILLER_349_1280 ();
 b15zdnd11an1n64x5 FILLER_349_1344 ();
 b15zdnd11an1n64x5 FILLER_349_1408 ();
 b15zdnd11an1n64x5 FILLER_349_1472 ();
 b15zdnd11an1n64x5 FILLER_349_1536 ();
 b15zdnd11an1n64x5 FILLER_349_1600 ();
 b15zdnd11an1n64x5 FILLER_349_1664 ();
 b15zdnd11an1n64x5 FILLER_349_1728 ();
 b15zdnd11an1n64x5 FILLER_349_1792 ();
 b15zdnd11an1n64x5 FILLER_349_1856 ();
 b15zdnd11an1n64x5 FILLER_349_1920 ();
 b15zdnd11an1n64x5 FILLER_349_1984 ();
 b15zdnd11an1n64x5 FILLER_349_2048 ();
 b15zdnd11an1n64x5 FILLER_349_2112 ();
 b15zdnd11an1n64x5 FILLER_349_2176 ();
 b15zdnd11an1n32x5 FILLER_349_2240 ();
 b15zdnd11an1n08x5 FILLER_349_2272 ();
 b15zdnd11an1n04x5 FILLER_349_2280 ();
 b15zdnd11an1n64x5 FILLER_350_8 ();
 b15zdnd11an1n64x5 FILLER_350_72 ();
 b15zdnd11an1n64x5 FILLER_350_136 ();
 b15zdnd11an1n64x5 FILLER_350_200 ();
 b15zdnd11an1n64x5 FILLER_350_264 ();
 b15zdnd11an1n64x5 FILLER_350_328 ();
 b15zdnd11an1n64x5 FILLER_350_392 ();
 b15zdnd11an1n64x5 FILLER_350_456 ();
 b15zdnd11an1n64x5 FILLER_350_520 ();
 b15zdnd11an1n64x5 FILLER_350_584 ();
 b15zdnd11an1n64x5 FILLER_350_648 ();
 b15zdnd11an1n04x5 FILLER_350_712 ();
 b15zdnd00an1n02x5 FILLER_350_716 ();
 b15zdnd11an1n64x5 FILLER_350_726 ();
 b15zdnd11an1n64x5 FILLER_350_790 ();
 b15zdnd11an1n64x5 FILLER_350_854 ();
 b15zdnd11an1n64x5 FILLER_350_918 ();
 b15zdnd11an1n64x5 FILLER_350_982 ();
 b15zdnd11an1n64x5 FILLER_350_1046 ();
 b15zdnd11an1n64x5 FILLER_350_1110 ();
 b15zdnd11an1n64x5 FILLER_350_1174 ();
 b15zdnd11an1n64x5 FILLER_350_1238 ();
 b15zdnd11an1n64x5 FILLER_350_1302 ();
 b15zdnd11an1n64x5 FILLER_350_1366 ();
 b15zdnd11an1n64x5 FILLER_350_1430 ();
 b15zdnd11an1n64x5 FILLER_350_1494 ();
 b15zdnd11an1n64x5 FILLER_350_1558 ();
 b15zdnd11an1n64x5 FILLER_350_1622 ();
 b15zdnd11an1n64x5 FILLER_350_1686 ();
 b15zdnd11an1n64x5 FILLER_350_1750 ();
 b15zdnd11an1n64x5 FILLER_350_1814 ();
 b15zdnd11an1n64x5 FILLER_350_1878 ();
 b15zdnd11an1n64x5 FILLER_350_1942 ();
 b15zdnd11an1n64x5 FILLER_350_2006 ();
 b15zdnd11an1n64x5 FILLER_350_2070 ();
 b15zdnd11an1n16x5 FILLER_350_2134 ();
 b15zdnd11an1n04x5 FILLER_350_2150 ();
 b15zdnd11an1n64x5 FILLER_350_2162 ();
 b15zdnd11an1n32x5 FILLER_350_2226 ();
 b15zdnd11an1n16x5 FILLER_350_2258 ();
 b15zdnd00an1n02x5 FILLER_350_2274 ();
 b15zdnd11an1n64x5 FILLER_351_0 ();
 b15zdnd11an1n64x5 FILLER_351_64 ();
 b15zdnd11an1n64x5 FILLER_351_128 ();
 b15zdnd11an1n64x5 FILLER_351_192 ();
 b15zdnd11an1n64x5 FILLER_351_256 ();
 b15zdnd11an1n64x5 FILLER_351_320 ();
 b15zdnd11an1n64x5 FILLER_351_384 ();
 b15zdnd11an1n64x5 FILLER_351_448 ();
 b15zdnd11an1n64x5 FILLER_351_512 ();
 b15zdnd11an1n64x5 FILLER_351_576 ();
 b15zdnd11an1n64x5 FILLER_351_640 ();
 b15zdnd11an1n64x5 FILLER_351_704 ();
 b15zdnd11an1n64x5 FILLER_351_768 ();
 b15zdnd11an1n64x5 FILLER_351_832 ();
 b15zdnd11an1n64x5 FILLER_351_896 ();
 b15zdnd11an1n64x5 FILLER_351_960 ();
 b15zdnd11an1n64x5 FILLER_351_1024 ();
 b15zdnd11an1n64x5 FILLER_351_1088 ();
 b15zdnd11an1n64x5 FILLER_351_1152 ();
 b15zdnd11an1n64x5 FILLER_351_1216 ();
 b15zdnd11an1n64x5 FILLER_351_1280 ();
 b15zdnd11an1n64x5 FILLER_351_1344 ();
 b15zdnd11an1n64x5 FILLER_351_1408 ();
 b15zdnd11an1n64x5 FILLER_351_1472 ();
 b15zdnd11an1n64x5 FILLER_351_1536 ();
 b15zdnd11an1n64x5 FILLER_351_1600 ();
 b15zdnd11an1n64x5 FILLER_351_1664 ();
 b15zdnd11an1n64x5 FILLER_351_1728 ();
 b15zdnd11an1n64x5 FILLER_351_1792 ();
 b15zdnd11an1n64x5 FILLER_351_1856 ();
 b15zdnd11an1n64x5 FILLER_351_1920 ();
 b15zdnd11an1n64x5 FILLER_351_1984 ();
 b15zdnd11an1n64x5 FILLER_351_2048 ();
 b15zdnd11an1n64x5 FILLER_351_2112 ();
 b15zdnd11an1n64x5 FILLER_351_2176 ();
 b15zdnd11an1n32x5 FILLER_351_2240 ();
 b15zdnd11an1n08x5 FILLER_351_2272 ();
 b15zdnd11an1n04x5 FILLER_351_2280 ();
 b15zdnd11an1n64x5 FILLER_352_8 ();
 b15zdnd11an1n64x5 FILLER_352_72 ();
 b15zdnd11an1n64x5 FILLER_352_136 ();
 b15zdnd11an1n64x5 FILLER_352_200 ();
 b15zdnd11an1n64x5 FILLER_352_264 ();
 b15zdnd11an1n64x5 FILLER_352_328 ();
 b15zdnd11an1n64x5 FILLER_352_392 ();
 b15zdnd11an1n64x5 FILLER_352_456 ();
 b15zdnd11an1n64x5 FILLER_352_520 ();
 b15zdnd11an1n64x5 FILLER_352_584 ();
 b15zdnd11an1n64x5 FILLER_352_648 ();
 b15zdnd11an1n04x5 FILLER_352_712 ();
 b15zdnd00an1n02x5 FILLER_352_716 ();
 b15zdnd11an1n64x5 FILLER_352_726 ();
 b15zdnd11an1n64x5 FILLER_352_790 ();
 b15zdnd11an1n64x5 FILLER_352_854 ();
 b15zdnd11an1n64x5 FILLER_352_918 ();
 b15zdnd11an1n64x5 FILLER_352_982 ();
 b15zdnd11an1n64x5 FILLER_352_1046 ();
 b15zdnd11an1n64x5 FILLER_352_1110 ();
 b15zdnd11an1n64x5 FILLER_352_1174 ();
 b15zdnd11an1n64x5 FILLER_352_1238 ();
 b15zdnd11an1n64x5 FILLER_352_1302 ();
 b15zdnd11an1n64x5 FILLER_352_1366 ();
 b15zdnd11an1n64x5 FILLER_352_1430 ();
 b15zdnd11an1n64x5 FILLER_352_1494 ();
 b15zdnd11an1n64x5 FILLER_352_1558 ();
 b15zdnd11an1n64x5 FILLER_352_1622 ();
 b15zdnd11an1n64x5 FILLER_352_1686 ();
 b15zdnd11an1n64x5 FILLER_352_1750 ();
 b15zdnd11an1n64x5 FILLER_352_1814 ();
 b15zdnd11an1n64x5 FILLER_352_1878 ();
 b15zdnd11an1n64x5 FILLER_352_1942 ();
 b15zdnd11an1n64x5 FILLER_352_2006 ();
 b15zdnd11an1n64x5 FILLER_352_2070 ();
 b15zdnd11an1n16x5 FILLER_352_2134 ();
 b15zdnd11an1n04x5 FILLER_352_2150 ();
 b15zdnd11an1n64x5 FILLER_352_2162 ();
 b15zdnd11an1n32x5 FILLER_352_2226 ();
 b15zdnd11an1n16x5 FILLER_352_2258 ();
 b15zdnd00an1n02x5 FILLER_352_2274 ();
 b15zdnd11an1n64x5 FILLER_353_0 ();
 b15zdnd11an1n64x5 FILLER_353_64 ();
 b15zdnd11an1n64x5 FILLER_353_128 ();
 b15zdnd11an1n64x5 FILLER_353_192 ();
 b15zdnd11an1n64x5 FILLER_353_256 ();
 b15zdnd11an1n64x5 FILLER_353_320 ();
 b15zdnd11an1n64x5 FILLER_353_384 ();
 b15zdnd11an1n64x5 FILLER_353_448 ();
 b15zdnd11an1n64x5 FILLER_353_512 ();
 b15zdnd11an1n64x5 FILLER_353_576 ();
 b15zdnd11an1n64x5 FILLER_353_640 ();
 b15zdnd11an1n64x5 FILLER_353_704 ();
 b15zdnd11an1n64x5 FILLER_353_768 ();
 b15zdnd11an1n64x5 FILLER_353_832 ();
 b15zdnd11an1n64x5 FILLER_353_896 ();
 b15zdnd11an1n64x5 FILLER_353_960 ();
 b15zdnd11an1n64x5 FILLER_353_1024 ();
 b15zdnd11an1n64x5 FILLER_353_1088 ();
 b15zdnd11an1n64x5 FILLER_353_1152 ();
 b15zdnd11an1n64x5 FILLER_353_1216 ();
 b15zdnd11an1n64x5 FILLER_353_1280 ();
 b15zdnd11an1n64x5 FILLER_353_1344 ();
 b15zdnd11an1n64x5 FILLER_353_1408 ();
 b15zdnd11an1n64x5 FILLER_353_1472 ();
 b15zdnd11an1n64x5 FILLER_353_1536 ();
 b15zdnd11an1n64x5 FILLER_353_1600 ();
 b15zdnd11an1n64x5 FILLER_353_1664 ();
 b15zdnd11an1n64x5 FILLER_353_1728 ();
 b15zdnd11an1n64x5 FILLER_353_1792 ();
 b15zdnd11an1n64x5 FILLER_353_1856 ();
 b15zdnd11an1n64x5 FILLER_353_1920 ();
 b15zdnd11an1n64x5 FILLER_353_1984 ();
 b15zdnd11an1n64x5 FILLER_353_2048 ();
 b15zdnd11an1n64x5 FILLER_353_2112 ();
 b15zdnd11an1n64x5 FILLER_353_2176 ();
 b15zdnd11an1n32x5 FILLER_353_2240 ();
 b15zdnd11an1n08x5 FILLER_353_2272 ();
 b15zdnd11an1n04x5 FILLER_353_2280 ();
 b15zdnd11an1n64x5 FILLER_354_8 ();
 b15zdnd11an1n64x5 FILLER_354_72 ();
 b15zdnd11an1n64x5 FILLER_354_136 ();
 b15zdnd11an1n64x5 FILLER_354_200 ();
 b15zdnd11an1n64x5 FILLER_354_264 ();
 b15zdnd11an1n64x5 FILLER_354_328 ();
 b15zdnd11an1n64x5 FILLER_354_392 ();
 b15zdnd11an1n64x5 FILLER_354_456 ();
 b15zdnd11an1n64x5 FILLER_354_520 ();
 b15zdnd11an1n64x5 FILLER_354_584 ();
 b15zdnd11an1n64x5 FILLER_354_648 ();
 b15zdnd11an1n04x5 FILLER_354_712 ();
 b15zdnd00an1n02x5 FILLER_354_716 ();
 b15zdnd11an1n64x5 FILLER_354_726 ();
 b15zdnd11an1n64x5 FILLER_354_790 ();
 b15zdnd11an1n64x5 FILLER_354_854 ();
 b15zdnd11an1n64x5 FILLER_354_918 ();
 b15zdnd11an1n64x5 FILLER_354_982 ();
 b15zdnd11an1n64x5 FILLER_354_1046 ();
 b15zdnd11an1n64x5 FILLER_354_1110 ();
 b15zdnd11an1n64x5 FILLER_354_1174 ();
 b15zdnd11an1n64x5 FILLER_354_1238 ();
 b15zdnd11an1n64x5 FILLER_354_1302 ();
 b15zdnd11an1n64x5 FILLER_354_1366 ();
 b15zdnd11an1n64x5 FILLER_354_1430 ();
 b15zdnd11an1n64x5 FILLER_354_1494 ();
 b15zdnd11an1n64x5 FILLER_354_1558 ();
 b15zdnd11an1n64x5 FILLER_354_1622 ();
 b15zdnd11an1n64x5 FILLER_354_1686 ();
 b15zdnd11an1n64x5 FILLER_354_1750 ();
 b15zdnd11an1n64x5 FILLER_354_1814 ();
 b15zdnd11an1n64x5 FILLER_354_1878 ();
 b15zdnd11an1n64x5 FILLER_354_1942 ();
 b15zdnd11an1n64x5 FILLER_354_2006 ();
 b15zdnd11an1n64x5 FILLER_354_2070 ();
 b15zdnd11an1n16x5 FILLER_354_2134 ();
 b15zdnd11an1n04x5 FILLER_354_2150 ();
 b15zdnd11an1n64x5 FILLER_354_2162 ();
 b15zdnd11an1n32x5 FILLER_354_2226 ();
 b15zdnd11an1n16x5 FILLER_354_2258 ();
 b15zdnd00an1n02x5 FILLER_354_2274 ();
 b15zdnd11an1n64x5 FILLER_355_0 ();
 b15zdnd11an1n64x5 FILLER_355_64 ();
 b15zdnd11an1n64x5 FILLER_355_128 ();
 b15zdnd11an1n64x5 FILLER_355_192 ();
 b15zdnd11an1n64x5 FILLER_355_256 ();
 b15zdnd11an1n64x5 FILLER_355_320 ();
 b15zdnd11an1n64x5 FILLER_355_384 ();
 b15zdnd11an1n64x5 FILLER_355_448 ();
 b15zdnd11an1n64x5 FILLER_355_512 ();
 b15zdnd11an1n64x5 FILLER_355_576 ();
 b15zdnd11an1n64x5 FILLER_355_640 ();
 b15zdnd11an1n64x5 FILLER_355_704 ();
 b15zdnd11an1n64x5 FILLER_355_768 ();
 b15zdnd11an1n64x5 FILLER_355_832 ();
 b15zdnd11an1n64x5 FILLER_355_896 ();
 b15zdnd11an1n64x5 FILLER_355_960 ();
 b15zdnd11an1n64x5 FILLER_355_1024 ();
 b15zdnd11an1n64x5 FILLER_355_1088 ();
 b15zdnd11an1n64x5 FILLER_355_1152 ();
 b15zdnd11an1n64x5 FILLER_355_1216 ();
 b15zdnd11an1n64x5 FILLER_355_1280 ();
 b15zdnd11an1n64x5 FILLER_355_1344 ();
 b15zdnd11an1n64x5 FILLER_355_1408 ();
 b15zdnd11an1n64x5 FILLER_355_1472 ();
 b15zdnd11an1n64x5 FILLER_355_1536 ();
 b15zdnd11an1n64x5 FILLER_355_1600 ();
 b15zdnd11an1n64x5 FILLER_355_1664 ();
 b15zdnd11an1n64x5 FILLER_355_1728 ();
 b15zdnd11an1n64x5 FILLER_355_1792 ();
 b15zdnd11an1n64x5 FILLER_355_1856 ();
 b15zdnd11an1n64x5 FILLER_355_1920 ();
 b15zdnd11an1n64x5 FILLER_355_1984 ();
 b15zdnd11an1n64x5 FILLER_355_2048 ();
 b15zdnd11an1n64x5 FILLER_355_2112 ();
 b15zdnd11an1n64x5 FILLER_355_2176 ();
 b15zdnd11an1n32x5 FILLER_355_2240 ();
 b15zdnd11an1n08x5 FILLER_355_2272 ();
 b15zdnd11an1n04x5 FILLER_355_2280 ();
 b15zdnd11an1n64x5 FILLER_356_8 ();
 b15zdnd11an1n64x5 FILLER_356_72 ();
 b15zdnd11an1n64x5 FILLER_356_136 ();
 b15zdnd11an1n64x5 FILLER_356_200 ();
 b15zdnd11an1n64x5 FILLER_356_264 ();
 b15zdnd11an1n64x5 FILLER_356_328 ();
 b15zdnd11an1n64x5 FILLER_356_392 ();
 b15zdnd11an1n64x5 FILLER_356_456 ();
 b15zdnd11an1n64x5 FILLER_356_520 ();
 b15zdnd11an1n64x5 FILLER_356_584 ();
 b15zdnd11an1n64x5 FILLER_356_648 ();
 b15zdnd11an1n04x5 FILLER_356_712 ();
 b15zdnd00an1n02x5 FILLER_356_716 ();
 b15zdnd11an1n64x5 FILLER_356_726 ();
 b15zdnd11an1n64x5 FILLER_356_790 ();
 b15zdnd11an1n64x5 FILLER_356_854 ();
 b15zdnd11an1n64x5 FILLER_356_918 ();
 b15zdnd11an1n64x5 FILLER_356_982 ();
 b15zdnd11an1n64x5 FILLER_356_1046 ();
 b15zdnd11an1n64x5 FILLER_356_1110 ();
 b15zdnd11an1n64x5 FILLER_356_1174 ();
 b15zdnd11an1n64x5 FILLER_356_1238 ();
 b15zdnd11an1n64x5 FILLER_356_1302 ();
 b15zdnd11an1n64x5 FILLER_356_1366 ();
 b15zdnd11an1n64x5 FILLER_356_1430 ();
 b15zdnd11an1n64x5 FILLER_356_1494 ();
 b15zdnd11an1n64x5 FILLER_356_1558 ();
 b15zdnd11an1n64x5 FILLER_356_1622 ();
 b15zdnd11an1n64x5 FILLER_356_1686 ();
 b15zdnd11an1n64x5 FILLER_356_1750 ();
 b15zdnd11an1n64x5 FILLER_356_1814 ();
 b15zdnd11an1n64x5 FILLER_356_1878 ();
 b15zdnd11an1n64x5 FILLER_356_1942 ();
 b15zdnd11an1n64x5 FILLER_356_2006 ();
 b15zdnd11an1n64x5 FILLER_356_2070 ();
 b15zdnd11an1n16x5 FILLER_356_2134 ();
 b15zdnd11an1n04x5 FILLER_356_2150 ();
 b15zdnd11an1n64x5 FILLER_356_2162 ();
 b15zdnd11an1n32x5 FILLER_356_2226 ();
 b15zdnd11an1n16x5 FILLER_356_2258 ();
 b15zdnd00an1n02x5 FILLER_356_2274 ();
 b15zdnd11an1n64x5 FILLER_357_0 ();
 b15zdnd11an1n64x5 FILLER_357_64 ();
 b15zdnd11an1n64x5 FILLER_357_128 ();
 b15zdnd11an1n64x5 FILLER_357_192 ();
 b15zdnd11an1n64x5 FILLER_357_256 ();
 b15zdnd11an1n64x5 FILLER_357_320 ();
 b15zdnd11an1n64x5 FILLER_357_384 ();
 b15zdnd11an1n64x5 FILLER_357_448 ();
 b15zdnd11an1n64x5 FILLER_357_512 ();
 b15zdnd11an1n64x5 FILLER_357_576 ();
 b15zdnd11an1n64x5 FILLER_357_640 ();
 b15zdnd11an1n64x5 FILLER_357_704 ();
 b15zdnd11an1n64x5 FILLER_357_768 ();
 b15zdnd11an1n64x5 FILLER_357_832 ();
 b15zdnd11an1n64x5 FILLER_357_896 ();
 b15zdnd11an1n64x5 FILLER_357_960 ();
 b15zdnd11an1n64x5 FILLER_357_1024 ();
 b15zdnd11an1n64x5 FILLER_357_1088 ();
 b15zdnd11an1n64x5 FILLER_357_1152 ();
 b15zdnd11an1n64x5 FILLER_357_1216 ();
 b15zdnd11an1n64x5 FILLER_357_1280 ();
 b15zdnd11an1n64x5 FILLER_357_1344 ();
 b15zdnd11an1n64x5 FILLER_357_1408 ();
 b15zdnd11an1n64x5 FILLER_357_1472 ();
 b15zdnd11an1n64x5 FILLER_357_1536 ();
 b15zdnd11an1n64x5 FILLER_357_1600 ();
 b15zdnd11an1n64x5 FILLER_357_1664 ();
 b15zdnd11an1n64x5 FILLER_357_1728 ();
 b15zdnd11an1n64x5 FILLER_357_1792 ();
 b15zdnd11an1n64x5 FILLER_357_1856 ();
 b15zdnd11an1n64x5 FILLER_357_1920 ();
 b15zdnd11an1n64x5 FILLER_357_1984 ();
 b15zdnd11an1n64x5 FILLER_357_2048 ();
 b15zdnd11an1n64x5 FILLER_357_2112 ();
 b15zdnd11an1n64x5 FILLER_357_2176 ();
 b15zdnd11an1n32x5 FILLER_357_2240 ();
 b15zdnd11an1n08x5 FILLER_357_2272 ();
 b15zdnd11an1n04x5 FILLER_357_2280 ();
 b15zdnd11an1n64x5 FILLER_358_8 ();
 b15zdnd11an1n64x5 FILLER_358_72 ();
 b15zdnd11an1n64x5 FILLER_358_136 ();
 b15zdnd11an1n64x5 FILLER_358_200 ();
 b15zdnd11an1n64x5 FILLER_358_264 ();
 b15zdnd11an1n64x5 FILLER_358_328 ();
 b15zdnd11an1n64x5 FILLER_358_392 ();
 b15zdnd11an1n64x5 FILLER_358_456 ();
 b15zdnd11an1n64x5 FILLER_358_520 ();
 b15zdnd11an1n64x5 FILLER_358_584 ();
 b15zdnd11an1n64x5 FILLER_358_648 ();
 b15zdnd11an1n04x5 FILLER_358_712 ();
 b15zdnd00an1n02x5 FILLER_358_716 ();
 b15zdnd11an1n64x5 FILLER_358_726 ();
 b15zdnd11an1n64x5 FILLER_358_790 ();
 b15zdnd11an1n64x5 FILLER_358_854 ();
 b15zdnd11an1n64x5 FILLER_358_918 ();
 b15zdnd11an1n64x5 FILLER_358_982 ();
 b15zdnd11an1n64x5 FILLER_358_1046 ();
 b15zdnd11an1n64x5 FILLER_358_1110 ();
 b15zdnd11an1n64x5 FILLER_358_1174 ();
 b15zdnd11an1n64x5 FILLER_358_1238 ();
 b15zdnd11an1n64x5 FILLER_358_1302 ();
 b15zdnd11an1n64x5 FILLER_358_1366 ();
 b15zdnd11an1n64x5 FILLER_358_1430 ();
 b15zdnd11an1n64x5 FILLER_358_1494 ();
 b15zdnd11an1n64x5 FILLER_358_1558 ();
 b15zdnd11an1n64x5 FILLER_358_1622 ();
 b15zdnd11an1n64x5 FILLER_358_1686 ();
 b15zdnd11an1n64x5 FILLER_358_1750 ();
 b15zdnd11an1n64x5 FILLER_358_1814 ();
 b15zdnd11an1n64x5 FILLER_358_1878 ();
 b15zdnd11an1n64x5 FILLER_358_1942 ();
 b15zdnd11an1n64x5 FILLER_358_2006 ();
 b15zdnd11an1n64x5 FILLER_358_2070 ();
 b15zdnd11an1n16x5 FILLER_358_2134 ();
 b15zdnd11an1n04x5 FILLER_358_2150 ();
 b15zdnd11an1n64x5 FILLER_358_2162 ();
 b15zdnd11an1n32x5 FILLER_358_2226 ();
 b15zdnd11an1n16x5 FILLER_358_2258 ();
 b15zdnd00an1n02x5 FILLER_358_2274 ();
 b15zdnd11an1n64x5 FILLER_359_0 ();
 b15zdnd11an1n64x5 FILLER_359_64 ();
 b15zdnd11an1n64x5 FILLER_359_128 ();
 b15zdnd11an1n64x5 FILLER_359_192 ();
 b15zdnd11an1n64x5 FILLER_359_256 ();
 b15zdnd11an1n64x5 FILLER_359_320 ();
 b15zdnd11an1n64x5 FILLER_359_384 ();
 b15zdnd11an1n64x5 FILLER_359_448 ();
 b15zdnd11an1n64x5 FILLER_359_512 ();
 b15zdnd11an1n64x5 FILLER_359_576 ();
 b15zdnd11an1n64x5 FILLER_359_640 ();
 b15zdnd11an1n64x5 FILLER_359_704 ();
 b15zdnd11an1n64x5 FILLER_359_768 ();
 b15zdnd11an1n64x5 FILLER_359_832 ();
 b15zdnd11an1n64x5 FILLER_359_896 ();
 b15zdnd11an1n64x5 FILLER_359_960 ();
 b15zdnd11an1n64x5 FILLER_359_1024 ();
 b15zdnd11an1n64x5 FILLER_359_1088 ();
 b15zdnd11an1n64x5 FILLER_359_1152 ();
 b15zdnd11an1n64x5 FILLER_359_1216 ();
 b15zdnd11an1n64x5 FILLER_359_1280 ();
 b15zdnd11an1n64x5 FILLER_359_1344 ();
 b15zdnd11an1n64x5 FILLER_359_1408 ();
 b15zdnd11an1n64x5 FILLER_359_1472 ();
 b15zdnd11an1n64x5 FILLER_359_1536 ();
 b15zdnd11an1n64x5 FILLER_359_1600 ();
 b15zdnd11an1n64x5 FILLER_359_1664 ();
 b15zdnd11an1n64x5 FILLER_359_1728 ();
 b15zdnd11an1n64x5 FILLER_359_1792 ();
 b15zdnd11an1n64x5 FILLER_359_1856 ();
 b15zdnd11an1n64x5 FILLER_359_1920 ();
 b15zdnd11an1n64x5 FILLER_359_1984 ();
 b15zdnd11an1n64x5 FILLER_359_2048 ();
 b15zdnd11an1n64x5 FILLER_359_2112 ();
 b15zdnd11an1n64x5 FILLER_359_2176 ();
 b15zdnd11an1n32x5 FILLER_359_2240 ();
 b15zdnd11an1n08x5 FILLER_359_2272 ();
 b15zdnd11an1n04x5 FILLER_359_2280 ();
 b15zdnd11an1n64x5 FILLER_360_8 ();
 b15zdnd11an1n64x5 FILLER_360_72 ();
 b15zdnd11an1n64x5 FILLER_360_136 ();
 b15zdnd11an1n64x5 FILLER_360_200 ();
 b15zdnd11an1n64x5 FILLER_360_264 ();
 b15zdnd11an1n64x5 FILLER_360_328 ();
 b15zdnd11an1n64x5 FILLER_360_392 ();
 b15zdnd11an1n64x5 FILLER_360_456 ();
 b15zdnd11an1n64x5 FILLER_360_520 ();
 b15zdnd11an1n64x5 FILLER_360_584 ();
 b15zdnd11an1n64x5 FILLER_360_648 ();
 b15zdnd11an1n04x5 FILLER_360_712 ();
 b15zdnd00an1n02x5 FILLER_360_716 ();
 b15zdnd11an1n64x5 FILLER_360_726 ();
 b15zdnd11an1n64x5 FILLER_360_790 ();
 b15zdnd11an1n64x5 FILLER_360_854 ();
 b15zdnd11an1n64x5 FILLER_360_918 ();
 b15zdnd11an1n64x5 FILLER_360_982 ();
 b15zdnd11an1n64x5 FILLER_360_1046 ();
 b15zdnd11an1n64x5 FILLER_360_1110 ();
 b15zdnd11an1n64x5 FILLER_360_1174 ();
 b15zdnd11an1n64x5 FILLER_360_1238 ();
 b15zdnd11an1n64x5 FILLER_360_1302 ();
 b15zdnd11an1n64x5 FILLER_360_1366 ();
 b15zdnd11an1n64x5 FILLER_360_1430 ();
 b15zdnd11an1n64x5 FILLER_360_1494 ();
 b15zdnd11an1n64x5 FILLER_360_1558 ();
 b15zdnd11an1n64x5 FILLER_360_1622 ();
 b15zdnd11an1n64x5 FILLER_360_1686 ();
 b15zdnd11an1n64x5 FILLER_360_1750 ();
 b15zdnd11an1n64x5 FILLER_360_1814 ();
 b15zdnd11an1n64x5 FILLER_360_1878 ();
 b15zdnd11an1n64x5 FILLER_360_1942 ();
 b15zdnd11an1n64x5 FILLER_360_2006 ();
 b15zdnd11an1n64x5 FILLER_360_2070 ();
 b15zdnd11an1n16x5 FILLER_360_2134 ();
 b15zdnd11an1n04x5 FILLER_360_2150 ();
 b15zdnd11an1n64x5 FILLER_360_2162 ();
 b15zdnd11an1n32x5 FILLER_360_2226 ();
 b15zdnd11an1n16x5 FILLER_360_2258 ();
 b15zdnd00an1n02x5 FILLER_360_2274 ();
 b15zdnd11an1n64x5 FILLER_361_0 ();
 b15zdnd11an1n64x5 FILLER_361_64 ();
 b15zdnd11an1n64x5 FILLER_361_128 ();
 b15zdnd11an1n64x5 FILLER_361_192 ();
 b15zdnd11an1n64x5 FILLER_361_256 ();
 b15zdnd11an1n64x5 FILLER_361_320 ();
 b15zdnd11an1n64x5 FILLER_361_384 ();
 b15zdnd11an1n64x5 FILLER_361_448 ();
 b15zdnd11an1n64x5 FILLER_361_512 ();
 b15zdnd11an1n64x5 FILLER_361_576 ();
 b15zdnd11an1n64x5 FILLER_361_640 ();
 b15zdnd11an1n64x5 FILLER_361_704 ();
 b15zdnd11an1n64x5 FILLER_361_768 ();
 b15zdnd11an1n64x5 FILLER_361_832 ();
 b15zdnd11an1n64x5 FILLER_361_896 ();
 b15zdnd11an1n64x5 FILLER_361_960 ();
 b15zdnd11an1n64x5 FILLER_361_1024 ();
 b15zdnd11an1n64x5 FILLER_361_1088 ();
 b15zdnd11an1n64x5 FILLER_361_1152 ();
 b15zdnd11an1n64x5 FILLER_361_1216 ();
 b15zdnd11an1n64x5 FILLER_361_1280 ();
 b15zdnd11an1n64x5 FILLER_361_1344 ();
 b15zdnd11an1n64x5 FILLER_361_1408 ();
 b15zdnd11an1n64x5 FILLER_361_1472 ();
 b15zdnd11an1n64x5 FILLER_361_1536 ();
 b15zdnd11an1n64x5 FILLER_361_1600 ();
 b15zdnd11an1n64x5 FILLER_361_1664 ();
 b15zdnd11an1n64x5 FILLER_361_1728 ();
 b15zdnd11an1n64x5 FILLER_361_1792 ();
 b15zdnd11an1n64x5 FILLER_361_1856 ();
 b15zdnd11an1n64x5 FILLER_361_1920 ();
 b15zdnd11an1n64x5 FILLER_361_1984 ();
 b15zdnd11an1n64x5 FILLER_361_2048 ();
 b15zdnd11an1n64x5 FILLER_361_2112 ();
 b15zdnd11an1n64x5 FILLER_361_2176 ();
 b15zdnd11an1n32x5 FILLER_361_2240 ();
 b15zdnd11an1n08x5 FILLER_361_2272 ();
 b15zdnd11an1n04x5 FILLER_361_2280 ();
 b15zdnd11an1n64x5 FILLER_362_8 ();
 b15zdnd11an1n64x5 FILLER_362_72 ();
 b15zdnd11an1n64x5 FILLER_362_136 ();
 b15zdnd11an1n64x5 FILLER_362_200 ();
 b15zdnd11an1n64x5 FILLER_362_264 ();
 b15zdnd11an1n64x5 FILLER_362_328 ();
 b15zdnd11an1n64x5 FILLER_362_392 ();
 b15zdnd11an1n64x5 FILLER_362_456 ();
 b15zdnd11an1n64x5 FILLER_362_520 ();
 b15zdnd11an1n64x5 FILLER_362_584 ();
 b15zdnd11an1n64x5 FILLER_362_648 ();
 b15zdnd11an1n04x5 FILLER_362_712 ();
 b15zdnd00an1n02x5 FILLER_362_716 ();
 b15zdnd11an1n64x5 FILLER_362_726 ();
 b15zdnd11an1n64x5 FILLER_362_790 ();
 b15zdnd11an1n64x5 FILLER_362_854 ();
 b15zdnd11an1n64x5 FILLER_362_918 ();
 b15zdnd11an1n64x5 FILLER_362_982 ();
 b15zdnd11an1n64x5 FILLER_362_1046 ();
 b15zdnd11an1n64x5 FILLER_362_1110 ();
 b15zdnd11an1n64x5 FILLER_362_1174 ();
 b15zdnd11an1n64x5 FILLER_362_1238 ();
 b15zdnd11an1n64x5 FILLER_362_1302 ();
 b15zdnd11an1n64x5 FILLER_362_1366 ();
 b15zdnd11an1n64x5 FILLER_362_1430 ();
 b15zdnd11an1n64x5 FILLER_362_1494 ();
 b15zdnd11an1n64x5 FILLER_362_1558 ();
 b15zdnd11an1n64x5 FILLER_362_1622 ();
 b15zdnd11an1n64x5 FILLER_362_1686 ();
 b15zdnd11an1n64x5 FILLER_362_1750 ();
 b15zdnd11an1n64x5 FILLER_362_1814 ();
 b15zdnd11an1n64x5 FILLER_362_1878 ();
 b15zdnd11an1n64x5 FILLER_362_1942 ();
 b15zdnd11an1n64x5 FILLER_362_2006 ();
 b15zdnd11an1n64x5 FILLER_362_2070 ();
 b15zdnd11an1n16x5 FILLER_362_2134 ();
 b15zdnd11an1n04x5 FILLER_362_2150 ();
 b15zdnd11an1n64x5 FILLER_362_2162 ();
 b15zdnd11an1n32x5 FILLER_362_2226 ();
 b15zdnd11an1n16x5 FILLER_362_2258 ();
 b15zdnd00an1n02x5 FILLER_362_2274 ();
 b15zdnd11an1n64x5 FILLER_363_0 ();
 b15zdnd11an1n64x5 FILLER_363_64 ();
 b15zdnd11an1n64x5 FILLER_363_128 ();
 b15zdnd11an1n64x5 FILLER_363_192 ();
 b15zdnd11an1n64x5 FILLER_363_256 ();
 b15zdnd11an1n64x5 FILLER_363_320 ();
 b15zdnd11an1n64x5 FILLER_363_384 ();
 b15zdnd11an1n64x5 FILLER_363_448 ();
 b15zdnd11an1n64x5 FILLER_363_512 ();
 b15zdnd11an1n64x5 FILLER_363_576 ();
 b15zdnd11an1n64x5 FILLER_363_640 ();
 b15zdnd11an1n64x5 FILLER_363_704 ();
 b15zdnd11an1n64x5 FILLER_363_768 ();
 b15zdnd11an1n64x5 FILLER_363_832 ();
 b15zdnd11an1n64x5 FILLER_363_896 ();
 b15zdnd11an1n64x5 FILLER_363_960 ();
 b15zdnd11an1n64x5 FILLER_363_1024 ();
 b15zdnd11an1n64x5 FILLER_363_1088 ();
 b15zdnd11an1n64x5 FILLER_363_1152 ();
 b15zdnd11an1n64x5 FILLER_363_1216 ();
 b15zdnd11an1n64x5 FILLER_363_1280 ();
 b15zdnd11an1n64x5 FILLER_363_1344 ();
 b15zdnd11an1n64x5 FILLER_363_1408 ();
 b15zdnd11an1n64x5 FILLER_363_1472 ();
 b15zdnd11an1n64x5 FILLER_363_1536 ();
 b15zdnd11an1n64x5 FILLER_363_1600 ();
 b15zdnd11an1n64x5 FILLER_363_1664 ();
 b15zdnd11an1n64x5 FILLER_363_1728 ();
 b15zdnd11an1n64x5 FILLER_363_1792 ();
 b15zdnd11an1n64x5 FILLER_363_1856 ();
 b15zdnd11an1n64x5 FILLER_363_1920 ();
 b15zdnd11an1n64x5 FILLER_363_1984 ();
 b15zdnd11an1n64x5 FILLER_363_2048 ();
 b15zdnd11an1n64x5 FILLER_363_2112 ();
 b15zdnd11an1n64x5 FILLER_363_2176 ();
 b15zdnd11an1n32x5 FILLER_363_2240 ();
 b15zdnd11an1n08x5 FILLER_363_2272 ();
 b15zdnd11an1n04x5 FILLER_363_2280 ();
 b15zdnd11an1n64x5 FILLER_364_8 ();
 b15zdnd11an1n64x5 FILLER_364_72 ();
 b15zdnd11an1n64x5 FILLER_364_136 ();
 b15zdnd11an1n64x5 FILLER_364_200 ();
 b15zdnd11an1n64x5 FILLER_364_264 ();
 b15zdnd11an1n64x5 FILLER_364_328 ();
 b15zdnd11an1n64x5 FILLER_364_392 ();
 b15zdnd11an1n64x5 FILLER_364_456 ();
 b15zdnd11an1n64x5 FILLER_364_520 ();
 b15zdnd11an1n64x5 FILLER_364_584 ();
 b15zdnd11an1n64x5 FILLER_364_648 ();
 b15zdnd11an1n04x5 FILLER_364_712 ();
 b15zdnd00an1n02x5 FILLER_364_716 ();
 b15zdnd11an1n64x5 FILLER_364_726 ();
 b15zdnd11an1n64x5 FILLER_364_790 ();
 b15zdnd11an1n64x5 FILLER_364_854 ();
 b15zdnd11an1n64x5 FILLER_364_918 ();
 b15zdnd11an1n64x5 FILLER_364_982 ();
 b15zdnd11an1n64x5 FILLER_364_1046 ();
 b15zdnd11an1n64x5 FILLER_364_1110 ();
 b15zdnd11an1n64x5 FILLER_364_1174 ();
 b15zdnd11an1n64x5 FILLER_364_1238 ();
 b15zdnd11an1n64x5 FILLER_364_1302 ();
 b15zdnd11an1n64x5 FILLER_364_1366 ();
 b15zdnd11an1n64x5 FILLER_364_1430 ();
 b15zdnd11an1n64x5 FILLER_364_1494 ();
 b15zdnd11an1n64x5 FILLER_364_1558 ();
 b15zdnd11an1n64x5 FILLER_364_1622 ();
 b15zdnd11an1n64x5 FILLER_364_1686 ();
 b15zdnd11an1n64x5 FILLER_364_1750 ();
 b15zdnd11an1n64x5 FILLER_364_1814 ();
 b15zdnd11an1n64x5 FILLER_364_1878 ();
 b15zdnd11an1n64x5 FILLER_364_1942 ();
 b15zdnd11an1n64x5 FILLER_364_2006 ();
 b15zdnd11an1n64x5 FILLER_364_2070 ();
 b15zdnd11an1n16x5 FILLER_364_2134 ();
 b15zdnd11an1n04x5 FILLER_364_2150 ();
 b15zdnd11an1n64x5 FILLER_364_2162 ();
 b15zdnd11an1n32x5 FILLER_364_2226 ();
 b15zdnd11an1n16x5 FILLER_364_2258 ();
 b15zdnd00an1n02x5 FILLER_364_2274 ();
 b15zdnd11an1n64x5 FILLER_365_0 ();
 b15zdnd11an1n64x5 FILLER_365_64 ();
 b15zdnd11an1n64x5 FILLER_365_128 ();
 b15zdnd11an1n64x5 FILLER_365_192 ();
 b15zdnd11an1n64x5 FILLER_365_256 ();
 b15zdnd11an1n64x5 FILLER_365_320 ();
 b15zdnd11an1n64x5 FILLER_365_384 ();
 b15zdnd11an1n64x5 FILLER_365_448 ();
 b15zdnd11an1n64x5 FILLER_365_512 ();
 b15zdnd11an1n64x5 FILLER_365_576 ();
 b15zdnd11an1n64x5 FILLER_365_640 ();
 b15zdnd11an1n64x5 FILLER_365_704 ();
 b15zdnd11an1n64x5 FILLER_365_768 ();
 b15zdnd11an1n64x5 FILLER_365_832 ();
 b15zdnd11an1n64x5 FILLER_365_896 ();
 b15zdnd11an1n64x5 FILLER_365_960 ();
 b15zdnd11an1n64x5 FILLER_365_1024 ();
 b15zdnd11an1n64x5 FILLER_365_1088 ();
 b15zdnd11an1n64x5 FILLER_365_1152 ();
 b15zdnd11an1n64x5 FILLER_365_1216 ();
 b15zdnd11an1n64x5 FILLER_365_1280 ();
 b15zdnd11an1n64x5 FILLER_365_1344 ();
 b15zdnd11an1n64x5 FILLER_365_1408 ();
 b15zdnd11an1n64x5 FILLER_365_1472 ();
 b15zdnd11an1n64x5 FILLER_365_1536 ();
 b15zdnd11an1n64x5 FILLER_365_1600 ();
 b15zdnd11an1n64x5 FILLER_365_1664 ();
 b15zdnd11an1n64x5 FILLER_365_1728 ();
 b15zdnd11an1n64x5 FILLER_365_1792 ();
 b15zdnd11an1n64x5 FILLER_365_1856 ();
 b15zdnd11an1n64x5 FILLER_365_1920 ();
 b15zdnd11an1n64x5 FILLER_365_1984 ();
 b15zdnd11an1n64x5 FILLER_365_2048 ();
 b15zdnd11an1n64x5 FILLER_365_2112 ();
 b15zdnd11an1n64x5 FILLER_365_2176 ();
 b15zdnd11an1n32x5 FILLER_365_2240 ();
 b15zdnd11an1n08x5 FILLER_365_2272 ();
 b15zdnd11an1n04x5 FILLER_365_2280 ();
 b15zdnd11an1n64x5 FILLER_366_8 ();
 b15zdnd11an1n64x5 FILLER_366_72 ();
 b15zdnd11an1n64x5 FILLER_366_136 ();
 b15zdnd11an1n64x5 FILLER_366_200 ();
 b15zdnd11an1n64x5 FILLER_366_264 ();
 b15zdnd11an1n64x5 FILLER_366_328 ();
 b15zdnd11an1n64x5 FILLER_366_392 ();
 b15zdnd11an1n64x5 FILLER_366_456 ();
 b15zdnd11an1n64x5 FILLER_366_520 ();
 b15zdnd11an1n64x5 FILLER_366_584 ();
 b15zdnd11an1n64x5 FILLER_366_648 ();
 b15zdnd11an1n04x5 FILLER_366_712 ();
 b15zdnd00an1n02x5 FILLER_366_716 ();
 b15zdnd11an1n64x5 FILLER_366_726 ();
 b15zdnd11an1n64x5 FILLER_366_790 ();
 b15zdnd11an1n64x5 FILLER_366_854 ();
 b15zdnd11an1n64x5 FILLER_366_918 ();
 b15zdnd11an1n64x5 FILLER_366_982 ();
 b15zdnd11an1n64x5 FILLER_366_1046 ();
 b15zdnd11an1n64x5 FILLER_366_1110 ();
 b15zdnd11an1n64x5 FILLER_366_1174 ();
 b15zdnd11an1n64x5 FILLER_366_1238 ();
 b15zdnd11an1n64x5 FILLER_366_1302 ();
 b15zdnd11an1n64x5 FILLER_366_1366 ();
 b15zdnd11an1n64x5 FILLER_366_1430 ();
 b15zdnd11an1n64x5 FILLER_366_1494 ();
 b15zdnd11an1n64x5 FILLER_366_1558 ();
 b15zdnd11an1n64x5 FILLER_366_1622 ();
 b15zdnd11an1n64x5 FILLER_366_1686 ();
 b15zdnd11an1n64x5 FILLER_366_1750 ();
 b15zdnd11an1n64x5 FILLER_366_1814 ();
 b15zdnd11an1n64x5 FILLER_366_1878 ();
 b15zdnd11an1n64x5 FILLER_366_1942 ();
 b15zdnd11an1n64x5 FILLER_366_2006 ();
 b15zdnd11an1n64x5 FILLER_366_2070 ();
 b15zdnd11an1n16x5 FILLER_366_2134 ();
 b15zdnd11an1n04x5 FILLER_366_2150 ();
 b15zdnd11an1n64x5 FILLER_366_2162 ();
 b15zdnd11an1n32x5 FILLER_366_2226 ();
 b15zdnd11an1n16x5 FILLER_366_2258 ();
 b15zdnd00an1n02x5 FILLER_366_2274 ();
 b15zdnd11an1n64x5 FILLER_367_0 ();
 b15zdnd11an1n64x5 FILLER_367_64 ();
 b15zdnd11an1n64x5 FILLER_367_128 ();
 b15zdnd11an1n64x5 FILLER_367_192 ();
 b15zdnd11an1n64x5 FILLER_367_256 ();
 b15zdnd11an1n64x5 FILLER_367_320 ();
 b15zdnd11an1n64x5 FILLER_367_384 ();
 b15zdnd11an1n64x5 FILLER_367_448 ();
 b15zdnd11an1n64x5 FILLER_367_512 ();
 b15zdnd11an1n64x5 FILLER_367_576 ();
 b15zdnd11an1n64x5 FILLER_367_640 ();
 b15zdnd11an1n64x5 FILLER_367_704 ();
 b15zdnd11an1n64x5 FILLER_367_768 ();
 b15zdnd11an1n64x5 FILLER_367_832 ();
 b15zdnd11an1n64x5 FILLER_367_896 ();
 b15zdnd11an1n64x5 FILLER_367_960 ();
 b15zdnd11an1n64x5 FILLER_367_1024 ();
 b15zdnd11an1n64x5 FILLER_367_1088 ();
 b15zdnd11an1n64x5 FILLER_367_1152 ();
 b15zdnd11an1n64x5 FILLER_367_1216 ();
 b15zdnd11an1n64x5 FILLER_367_1280 ();
 b15zdnd11an1n64x5 FILLER_367_1344 ();
 b15zdnd11an1n64x5 FILLER_367_1408 ();
 b15zdnd11an1n64x5 FILLER_367_1472 ();
 b15zdnd11an1n64x5 FILLER_367_1536 ();
 b15zdnd11an1n64x5 FILLER_367_1600 ();
 b15zdnd11an1n64x5 FILLER_367_1664 ();
 b15zdnd11an1n64x5 FILLER_367_1728 ();
 b15zdnd11an1n64x5 FILLER_367_1792 ();
 b15zdnd11an1n64x5 FILLER_367_1856 ();
 b15zdnd11an1n64x5 FILLER_367_1920 ();
 b15zdnd11an1n64x5 FILLER_367_1984 ();
 b15zdnd11an1n64x5 FILLER_367_2048 ();
 b15zdnd11an1n64x5 FILLER_367_2112 ();
 b15zdnd11an1n64x5 FILLER_367_2176 ();
 b15zdnd11an1n32x5 FILLER_367_2240 ();
 b15zdnd11an1n08x5 FILLER_367_2272 ();
 b15zdnd11an1n04x5 FILLER_367_2280 ();
 b15zdnd11an1n64x5 FILLER_368_8 ();
 b15zdnd11an1n64x5 FILLER_368_72 ();
 b15zdnd11an1n64x5 FILLER_368_136 ();
 b15zdnd11an1n64x5 FILLER_368_200 ();
 b15zdnd11an1n64x5 FILLER_368_264 ();
 b15zdnd11an1n64x5 FILLER_368_328 ();
 b15zdnd11an1n64x5 FILLER_368_392 ();
 b15zdnd11an1n64x5 FILLER_368_456 ();
 b15zdnd11an1n64x5 FILLER_368_520 ();
 b15zdnd11an1n64x5 FILLER_368_584 ();
 b15zdnd11an1n64x5 FILLER_368_648 ();
 b15zdnd11an1n04x5 FILLER_368_712 ();
 b15zdnd00an1n02x5 FILLER_368_716 ();
 b15zdnd11an1n64x5 FILLER_368_726 ();
 b15zdnd11an1n64x5 FILLER_368_790 ();
 b15zdnd11an1n64x5 FILLER_368_854 ();
 b15zdnd11an1n64x5 FILLER_368_918 ();
 b15zdnd11an1n64x5 FILLER_368_982 ();
 b15zdnd11an1n64x5 FILLER_368_1046 ();
 b15zdnd11an1n64x5 FILLER_368_1110 ();
 b15zdnd11an1n64x5 FILLER_368_1174 ();
 b15zdnd11an1n64x5 FILLER_368_1238 ();
 b15zdnd11an1n64x5 FILLER_368_1302 ();
 b15zdnd11an1n64x5 FILLER_368_1366 ();
 b15zdnd11an1n64x5 FILLER_368_1430 ();
 b15zdnd11an1n64x5 FILLER_368_1494 ();
 b15zdnd11an1n64x5 FILLER_368_1558 ();
 b15zdnd11an1n64x5 FILLER_368_1622 ();
 b15zdnd11an1n64x5 FILLER_368_1686 ();
 b15zdnd11an1n64x5 FILLER_368_1750 ();
 b15zdnd11an1n64x5 FILLER_368_1814 ();
 b15zdnd11an1n64x5 FILLER_368_1878 ();
 b15zdnd11an1n64x5 FILLER_368_1942 ();
 b15zdnd11an1n64x5 FILLER_368_2006 ();
 b15zdnd11an1n64x5 FILLER_368_2070 ();
 b15zdnd11an1n16x5 FILLER_368_2134 ();
 b15zdnd11an1n04x5 FILLER_368_2150 ();
 b15zdnd11an1n64x5 FILLER_368_2162 ();
 b15zdnd11an1n32x5 FILLER_368_2226 ();
 b15zdnd11an1n16x5 FILLER_368_2258 ();
 b15zdnd00an1n02x5 FILLER_368_2274 ();
 b15zdnd11an1n64x5 FILLER_369_0 ();
 b15zdnd11an1n64x5 FILLER_369_64 ();
 b15zdnd11an1n64x5 FILLER_369_128 ();
 b15zdnd11an1n64x5 FILLER_369_192 ();
 b15zdnd11an1n64x5 FILLER_369_256 ();
 b15zdnd11an1n64x5 FILLER_369_320 ();
 b15zdnd11an1n64x5 FILLER_369_384 ();
 b15zdnd11an1n64x5 FILLER_369_448 ();
 b15zdnd11an1n64x5 FILLER_369_512 ();
 b15zdnd11an1n64x5 FILLER_369_576 ();
 b15zdnd11an1n64x5 FILLER_369_640 ();
 b15zdnd11an1n64x5 FILLER_369_704 ();
 b15zdnd11an1n64x5 FILLER_369_768 ();
 b15zdnd11an1n64x5 FILLER_369_832 ();
 b15zdnd11an1n64x5 FILLER_369_896 ();
 b15zdnd11an1n64x5 FILLER_369_960 ();
 b15zdnd11an1n64x5 FILLER_369_1024 ();
 b15zdnd11an1n64x5 FILLER_369_1088 ();
 b15zdnd11an1n64x5 FILLER_369_1152 ();
 b15zdnd11an1n64x5 FILLER_369_1216 ();
 b15zdnd11an1n64x5 FILLER_369_1280 ();
 b15zdnd11an1n64x5 FILLER_369_1344 ();
 b15zdnd11an1n64x5 FILLER_369_1408 ();
 b15zdnd11an1n64x5 FILLER_369_1472 ();
 b15zdnd11an1n64x5 FILLER_369_1536 ();
 b15zdnd11an1n64x5 FILLER_369_1600 ();
 b15zdnd11an1n64x5 FILLER_369_1664 ();
 b15zdnd11an1n64x5 FILLER_369_1728 ();
 b15zdnd11an1n64x5 FILLER_369_1792 ();
 b15zdnd11an1n64x5 FILLER_369_1856 ();
 b15zdnd11an1n64x5 FILLER_369_1920 ();
 b15zdnd11an1n64x5 FILLER_369_1984 ();
 b15zdnd11an1n64x5 FILLER_369_2048 ();
 b15zdnd11an1n64x5 FILLER_369_2112 ();
 b15zdnd11an1n64x5 FILLER_369_2176 ();
 b15zdnd11an1n32x5 FILLER_369_2240 ();
 b15zdnd11an1n08x5 FILLER_369_2272 ();
 b15zdnd11an1n04x5 FILLER_369_2280 ();
 b15zdnd11an1n64x5 FILLER_370_8 ();
 b15zdnd11an1n64x5 FILLER_370_72 ();
 b15zdnd11an1n64x5 FILLER_370_136 ();
 b15zdnd11an1n64x5 FILLER_370_200 ();
 b15zdnd11an1n64x5 FILLER_370_264 ();
 b15zdnd11an1n64x5 FILLER_370_328 ();
 b15zdnd11an1n64x5 FILLER_370_392 ();
 b15zdnd11an1n64x5 FILLER_370_456 ();
 b15zdnd11an1n64x5 FILLER_370_520 ();
 b15zdnd11an1n64x5 FILLER_370_584 ();
 b15zdnd11an1n64x5 FILLER_370_648 ();
 b15zdnd11an1n04x5 FILLER_370_712 ();
 b15zdnd00an1n02x5 FILLER_370_716 ();
 b15zdnd11an1n64x5 FILLER_370_726 ();
 b15zdnd11an1n64x5 FILLER_370_790 ();
 b15zdnd11an1n64x5 FILLER_370_854 ();
 b15zdnd11an1n64x5 FILLER_370_918 ();
 b15zdnd11an1n64x5 FILLER_370_982 ();
 b15zdnd11an1n64x5 FILLER_370_1046 ();
 b15zdnd11an1n64x5 FILLER_370_1110 ();
 b15zdnd11an1n64x5 FILLER_370_1174 ();
 b15zdnd11an1n64x5 FILLER_370_1238 ();
 b15zdnd11an1n64x5 FILLER_370_1302 ();
 b15zdnd11an1n64x5 FILLER_370_1366 ();
 b15zdnd11an1n64x5 FILLER_370_1430 ();
 b15zdnd11an1n64x5 FILLER_370_1494 ();
 b15zdnd11an1n64x5 FILLER_370_1558 ();
 b15zdnd11an1n64x5 FILLER_370_1622 ();
 b15zdnd11an1n64x5 FILLER_370_1686 ();
 b15zdnd11an1n64x5 FILLER_370_1750 ();
 b15zdnd11an1n64x5 FILLER_370_1814 ();
 b15zdnd11an1n64x5 FILLER_370_1878 ();
 b15zdnd11an1n64x5 FILLER_370_1942 ();
 b15zdnd11an1n64x5 FILLER_370_2006 ();
 b15zdnd11an1n64x5 FILLER_370_2070 ();
 b15zdnd11an1n16x5 FILLER_370_2134 ();
 b15zdnd11an1n04x5 FILLER_370_2150 ();
 b15zdnd11an1n64x5 FILLER_370_2162 ();
 b15zdnd11an1n32x5 FILLER_370_2226 ();
 b15zdnd11an1n16x5 FILLER_370_2258 ();
 b15zdnd00an1n02x5 FILLER_370_2274 ();
 b15zdnd11an1n64x5 FILLER_371_0 ();
 b15zdnd11an1n64x5 FILLER_371_64 ();
 b15zdnd11an1n64x5 FILLER_371_128 ();
 b15zdnd11an1n64x5 FILLER_371_192 ();
 b15zdnd11an1n64x5 FILLER_371_256 ();
 b15zdnd11an1n64x5 FILLER_371_320 ();
 b15zdnd11an1n64x5 FILLER_371_384 ();
 b15zdnd11an1n64x5 FILLER_371_448 ();
 b15zdnd11an1n64x5 FILLER_371_512 ();
 b15zdnd11an1n64x5 FILLER_371_576 ();
 b15zdnd11an1n64x5 FILLER_371_640 ();
 b15zdnd11an1n64x5 FILLER_371_704 ();
 b15zdnd11an1n64x5 FILLER_371_768 ();
 b15zdnd11an1n64x5 FILLER_371_832 ();
 b15zdnd11an1n64x5 FILLER_371_896 ();
 b15zdnd11an1n64x5 FILLER_371_960 ();
 b15zdnd11an1n64x5 FILLER_371_1024 ();
 b15zdnd11an1n64x5 FILLER_371_1088 ();
 b15zdnd11an1n64x5 FILLER_371_1152 ();
 b15zdnd11an1n64x5 FILLER_371_1216 ();
 b15zdnd11an1n64x5 FILLER_371_1280 ();
 b15zdnd11an1n64x5 FILLER_371_1344 ();
 b15zdnd11an1n64x5 FILLER_371_1408 ();
 b15zdnd11an1n64x5 FILLER_371_1472 ();
 b15zdnd11an1n64x5 FILLER_371_1536 ();
 b15zdnd11an1n64x5 FILLER_371_1600 ();
 b15zdnd11an1n64x5 FILLER_371_1664 ();
 b15zdnd11an1n64x5 FILLER_371_1728 ();
 b15zdnd11an1n64x5 FILLER_371_1792 ();
 b15zdnd11an1n64x5 FILLER_371_1856 ();
 b15zdnd11an1n64x5 FILLER_371_1920 ();
 b15zdnd11an1n64x5 FILLER_371_1984 ();
 b15zdnd11an1n64x5 FILLER_371_2048 ();
 b15zdnd11an1n64x5 FILLER_371_2112 ();
 b15zdnd11an1n64x5 FILLER_371_2176 ();
 b15zdnd11an1n32x5 FILLER_371_2240 ();
 b15zdnd11an1n08x5 FILLER_371_2272 ();
 b15zdnd11an1n04x5 FILLER_371_2280 ();
 b15zdnd11an1n64x5 FILLER_372_8 ();
 b15zdnd11an1n64x5 FILLER_372_72 ();
 b15zdnd11an1n64x5 FILLER_372_136 ();
 b15zdnd11an1n64x5 FILLER_372_200 ();
 b15zdnd11an1n64x5 FILLER_372_264 ();
 b15zdnd11an1n64x5 FILLER_372_328 ();
 b15zdnd11an1n64x5 FILLER_372_392 ();
 b15zdnd11an1n64x5 FILLER_372_456 ();
 b15zdnd11an1n64x5 FILLER_372_520 ();
 b15zdnd11an1n64x5 FILLER_372_584 ();
 b15zdnd11an1n64x5 FILLER_372_648 ();
 b15zdnd11an1n04x5 FILLER_372_712 ();
 b15zdnd00an1n02x5 FILLER_372_716 ();
 b15zdnd11an1n64x5 FILLER_372_726 ();
 b15zdnd11an1n64x5 FILLER_372_790 ();
 b15zdnd11an1n64x5 FILLER_372_854 ();
 b15zdnd11an1n64x5 FILLER_372_918 ();
 b15zdnd11an1n64x5 FILLER_372_982 ();
 b15zdnd11an1n64x5 FILLER_372_1046 ();
 b15zdnd11an1n64x5 FILLER_372_1110 ();
 b15zdnd11an1n64x5 FILLER_372_1174 ();
 b15zdnd11an1n64x5 FILLER_372_1238 ();
 b15zdnd11an1n64x5 FILLER_372_1302 ();
 b15zdnd11an1n64x5 FILLER_372_1366 ();
 b15zdnd11an1n64x5 FILLER_372_1430 ();
 b15zdnd11an1n64x5 FILLER_372_1494 ();
 b15zdnd11an1n64x5 FILLER_372_1558 ();
 b15zdnd11an1n64x5 FILLER_372_1622 ();
 b15zdnd11an1n64x5 FILLER_372_1686 ();
 b15zdnd11an1n64x5 FILLER_372_1750 ();
 b15zdnd11an1n64x5 FILLER_372_1814 ();
 b15zdnd11an1n64x5 FILLER_372_1878 ();
 b15zdnd11an1n64x5 FILLER_372_1942 ();
 b15zdnd11an1n64x5 FILLER_372_2006 ();
 b15zdnd11an1n64x5 FILLER_372_2070 ();
 b15zdnd11an1n16x5 FILLER_372_2134 ();
 b15zdnd11an1n04x5 FILLER_372_2150 ();
 b15zdnd11an1n64x5 FILLER_372_2162 ();
 b15zdnd11an1n32x5 FILLER_372_2226 ();
 b15zdnd11an1n16x5 FILLER_372_2258 ();
 b15zdnd00an1n02x5 FILLER_372_2274 ();
 b15zdnd11an1n64x5 FILLER_373_0 ();
 b15zdnd11an1n64x5 FILLER_373_64 ();
 b15zdnd11an1n64x5 FILLER_373_128 ();
 b15zdnd11an1n64x5 FILLER_373_192 ();
 b15zdnd11an1n64x5 FILLER_373_256 ();
 b15zdnd11an1n64x5 FILLER_373_320 ();
 b15zdnd11an1n64x5 FILLER_373_384 ();
 b15zdnd11an1n64x5 FILLER_373_448 ();
 b15zdnd11an1n64x5 FILLER_373_512 ();
 b15zdnd11an1n64x5 FILLER_373_576 ();
 b15zdnd11an1n64x5 FILLER_373_640 ();
 b15zdnd11an1n64x5 FILLER_373_704 ();
 b15zdnd11an1n64x5 FILLER_373_768 ();
 b15zdnd11an1n64x5 FILLER_373_832 ();
 b15zdnd11an1n64x5 FILLER_373_896 ();
 b15zdnd11an1n64x5 FILLER_373_960 ();
 b15zdnd11an1n64x5 FILLER_373_1024 ();
 b15zdnd11an1n64x5 FILLER_373_1088 ();
 b15zdnd11an1n64x5 FILLER_373_1152 ();
 b15zdnd11an1n64x5 FILLER_373_1216 ();
 b15zdnd11an1n64x5 FILLER_373_1280 ();
 b15zdnd11an1n64x5 FILLER_373_1344 ();
 b15zdnd11an1n64x5 FILLER_373_1408 ();
 b15zdnd11an1n64x5 FILLER_373_1472 ();
 b15zdnd11an1n64x5 FILLER_373_1536 ();
 b15zdnd11an1n64x5 FILLER_373_1600 ();
 b15zdnd11an1n64x5 FILLER_373_1664 ();
 b15zdnd11an1n64x5 FILLER_373_1728 ();
 b15zdnd11an1n64x5 FILLER_373_1792 ();
 b15zdnd11an1n64x5 FILLER_373_1856 ();
 b15zdnd11an1n64x5 FILLER_373_1920 ();
 b15zdnd11an1n64x5 FILLER_373_1984 ();
 b15zdnd11an1n64x5 FILLER_373_2048 ();
 b15zdnd11an1n64x5 FILLER_373_2112 ();
 b15zdnd11an1n64x5 FILLER_373_2176 ();
 b15zdnd11an1n32x5 FILLER_373_2240 ();
 b15zdnd11an1n08x5 FILLER_373_2272 ();
 b15zdnd11an1n04x5 FILLER_373_2280 ();
 b15zdnd11an1n64x5 FILLER_374_8 ();
 b15zdnd11an1n64x5 FILLER_374_72 ();
 b15zdnd11an1n64x5 FILLER_374_136 ();
 b15zdnd11an1n64x5 FILLER_374_200 ();
 b15zdnd11an1n64x5 FILLER_374_264 ();
 b15zdnd11an1n64x5 FILLER_374_328 ();
 b15zdnd11an1n64x5 FILLER_374_392 ();
 b15zdnd11an1n64x5 FILLER_374_456 ();
 b15zdnd11an1n64x5 FILLER_374_520 ();
 b15zdnd11an1n64x5 FILLER_374_584 ();
 b15zdnd11an1n64x5 FILLER_374_648 ();
 b15zdnd11an1n04x5 FILLER_374_712 ();
 b15zdnd00an1n02x5 FILLER_374_716 ();
 b15zdnd11an1n64x5 FILLER_374_726 ();
 b15zdnd11an1n64x5 FILLER_374_790 ();
 b15zdnd11an1n64x5 FILLER_374_854 ();
 b15zdnd11an1n64x5 FILLER_374_918 ();
 b15zdnd11an1n64x5 FILLER_374_982 ();
 b15zdnd11an1n64x5 FILLER_374_1046 ();
 b15zdnd11an1n64x5 FILLER_374_1110 ();
 b15zdnd11an1n64x5 FILLER_374_1174 ();
 b15zdnd11an1n64x5 FILLER_374_1238 ();
 b15zdnd11an1n64x5 FILLER_374_1302 ();
 b15zdnd11an1n64x5 FILLER_374_1366 ();
 b15zdnd11an1n64x5 FILLER_374_1430 ();
 b15zdnd11an1n64x5 FILLER_374_1494 ();
 b15zdnd11an1n64x5 FILLER_374_1558 ();
 b15zdnd11an1n64x5 FILLER_374_1622 ();
 b15zdnd11an1n64x5 FILLER_374_1686 ();
 b15zdnd11an1n64x5 FILLER_374_1750 ();
 b15zdnd11an1n64x5 FILLER_374_1814 ();
 b15zdnd11an1n64x5 FILLER_374_1878 ();
 b15zdnd11an1n64x5 FILLER_374_1942 ();
 b15zdnd11an1n64x5 FILLER_374_2006 ();
 b15zdnd11an1n64x5 FILLER_374_2070 ();
 b15zdnd11an1n16x5 FILLER_374_2134 ();
 b15zdnd11an1n04x5 FILLER_374_2150 ();
 b15zdnd11an1n64x5 FILLER_374_2162 ();
 b15zdnd11an1n32x5 FILLER_374_2226 ();
 b15zdnd11an1n16x5 FILLER_374_2258 ();
 b15zdnd00an1n02x5 FILLER_374_2274 ();
 b15zdnd11an1n64x5 FILLER_375_0 ();
 b15zdnd11an1n64x5 FILLER_375_64 ();
 b15zdnd11an1n64x5 FILLER_375_128 ();
 b15zdnd11an1n64x5 FILLER_375_192 ();
 b15zdnd11an1n64x5 FILLER_375_256 ();
 b15zdnd11an1n64x5 FILLER_375_320 ();
 b15zdnd11an1n64x5 FILLER_375_384 ();
 b15zdnd11an1n64x5 FILLER_375_448 ();
 b15zdnd11an1n64x5 FILLER_375_512 ();
 b15zdnd11an1n64x5 FILLER_375_576 ();
 b15zdnd11an1n64x5 FILLER_375_640 ();
 b15zdnd11an1n64x5 FILLER_375_704 ();
 b15zdnd11an1n64x5 FILLER_375_768 ();
 b15zdnd11an1n64x5 FILLER_375_832 ();
 b15zdnd11an1n64x5 FILLER_375_896 ();
 b15zdnd11an1n64x5 FILLER_375_960 ();
 b15zdnd11an1n64x5 FILLER_375_1024 ();
 b15zdnd11an1n64x5 FILLER_375_1088 ();
 b15zdnd11an1n64x5 FILLER_375_1152 ();
 b15zdnd11an1n64x5 FILLER_375_1216 ();
 b15zdnd11an1n64x5 FILLER_375_1280 ();
 b15zdnd11an1n64x5 FILLER_375_1344 ();
 b15zdnd11an1n64x5 FILLER_375_1408 ();
 b15zdnd11an1n64x5 FILLER_375_1472 ();
 b15zdnd11an1n64x5 FILLER_375_1536 ();
 b15zdnd11an1n64x5 FILLER_375_1600 ();
 b15zdnd11an1n64x5 FILLER_375_1664 ();
 b15zdnd11an1n64x5 FILLER_375_1728 ();
 b15zdnd11an1n64x5 FILLER_375_1792 ();
 b15zdnd11an1n64x5 FILLER_375_1856 ();
 b15zdnd11an1n64x5 FILLER_375_1920 ();
 b15zdnd11an1n64x5 FILLER_375_1984 ();
 b15zdnd11an1n64x5 FILLER_375_2048 ();
 b15zdnd11an1n64x5 FILLER_375_2112 ();
 b15zdnd11an1n64x5 FILLER_375_2176 ();
 b15zdnd11an1n32x5 FILLER_375_2240 ();
 b15zdnd11an1n08x5 FILLER_375_2272 ();
 b15zdnd11an1n04x5 FILLER_375_2280 ();
 b15zdnd11an1n64x5 FILLER_376_8 ();
 b15zdnd11an1n64x5 FILLER_376_72 ();
 b15zdnd11an1n64x5 FILLER_376_136 ();
 b15zdnd11an1n64x5 FILLER_376_200 ();
 b15zdnd11an1n64x5 FILLER_376_264 ();
 b15zdnd11an1n64x5 FILLER_376_328 ();
 b15zdnd11an1n64x5 FILLER_376_392 ();
 b15zdnd11an1n64x5 FILLER_376_456 ();
 b15zdnd11an1n64x5 FILLER_376_520 ();
 b15zdnd11an1n64x5 FILLER_376_584 ();
 b15zdnd11an1n64x5 FILLER_376_648 ();
 b15zdnd11an1n04x5 FILLER_376_712 ();
 b15zdnd00an1n02x5 FILLER_376_716 ();
 b15zdnd11an1n64x5 FILLER_376_726 ();
 b15zdnd11an1n64x5 FILLER_376_790 ();
 b15zdnd11an1n64x5 FILLER_376_854 ();
 b15zdnd11an1n64x5 FILLER_376_918 ();
 b15zdnd11an1n64x5 FILLER_376_982 ();
 b15zdnd11an1n64x5 FILLER_376_1046 ();
 b15zdnd11an1n64x5 FILLER_376_1110 ();
 b15zdnd11an1n64x5 FILLER_376_1174 ();
 b15zdnd11an1n64x5 FILLER_376_1238 ();
 b15zdnd11an1n64x5 FILLER_376_1302 ();
 b15zdnd11an1n64x5 FILLER_376_1366 ();
 b15zdnd11an1n64x5 FILLER_376_1430 ();
 b15zdnd11an1n64x5 FILLER_376_1494 ();
 b15zdnd11an1n64x5 FILLER_376_1558 ();
 b15zdnd11an1n64x5 FILLER_376_1622 ();
 b15zdnd11an1n64x5 FILLER_376_1686 ();
 b15zdnd11an1n64x5 FILLER_376_1750 ();
 b15zdnd11an1n64x5 FILLER_376_1814 ();
 b15zdnd11an1n64x5 FILLER_376_1878 ();
 b15zdnd11an1n64x5 FILLER_376_1942 ();
 b15zdnd11an1n64x5 FILLER_376_2006 ();
 b15zdnd11an1n64x5 FILLER_376_2070 ();
 b15zdnd11an1n16x5 FILLER_376_2134 ();
 b15zdnd11an1n04x5 FILLER_376_2150 ();
 b15zdnd11an1n64x5 FILLER_376_2162 ();
 b15zdnd11an1n32x5 FILLER_376_2226 ();
 b15zdnd11an1n16x5 FILLER_376_2258 ();
 b15zdnd00an1n02x5 FILLER_376_2274 ();
 b15zdnd11an1n64x5 FILLER_377_0 ();
 b15zdnd11an1n64x5 FILLER_377_64 ();
 b15zdnd11an1n64x5 FILLER_377_128 ();
 b15zdnd11an1n64x5 FILLER_377_192 ();
 b15zdnd11an1n64x5 FILLER_377_256 ();
 b15zdnd11an1n64x5 FILLER_377_320 ();
 b15zdnd11an1n64x5 FILLER_377_384 ();
 b15zdnd11an1n64x5 FILLER_377_448 ();
 b15zdnd11an1n64x5 FILLER_377_512 ();
 b15zdnd11an1n64x5 FILLER_377_576 ();
 b15zdnd11an1n64x5 FILLER_377_640 ();
 b15zdnd11an1n64x5 FILLER_377_704 ();
 b15zdnd11an1n64x5 FILLER_377_768 ();
 b15zdnd11an1n64x5 FILLER_377_832 ();
 b15zdnd11an1n64x5 FILLER_377_896 ();
 b15zdnd11an1n64x5 FILLER_377_960 ();
 b15zdnd11an1n64x5 FILLER_377_1024 ();
 b15zdnd11an1n64x5 FILLER_377_1088 ();
 b15zdnd11an1n64x5 FILLER_377_1152 ();
 b15zdnd11an1n64x5 FILLER_377_1216 ();
 b15zdnd11an1n64x5 FILLER_377_1280 ();
 b15zdnd11an1n64x5 FILLER_377_1344 ();
 b15zdnd11an1n64x5 FILLER_377_1408 ();
 b15zdnd11an1n64x5 FILLER_377_1472 ();
 b15zdnd11an1n64x5 FILLER_377_1536 ();
 b15zdnd11an1n64x5 FILLER_377_1600 ();
 b15zdnd11an1n64x5 FILLER_377_1664 ();
 b15zdnd11an1n64x5 FILLER_377_1728 ();
 b15zdnd11an1n64x5 FILLER_377_1792 ();
 b15zdnd11an1n64x5 FILLER_377_1856 ();
 b15zdnd11an1n64x5 FILLER_377_1920 ();
 b15zdnd11an1n64x5 FILLER_377_1984 ();
 b15zdnd11an1n64x5 FILLER_377_2048 ();
 b15zdnd11an1n64x5 FILLER_377_2112 ();
 b15zdnd11an1n64x5 FILLER_377_2176 ();
 b15zdnd11an1n32x5 FILLER_377_2240 ();
 b15zdnd11an1n08x5 FILLER_377_2272 ();
 b15zdnd11an1n04x5 FILLER_377_2280 ();
 b15zdnd11an1n64x5 FILLER_378_8 ();
 b15zdnd11an1n64x5 FILLER_378_72 ();
 b15zdnd11an1n64x5 FILLER_378_136 ();
 b15zdnd11an1n64x5 FILLER_378_200 ();
 b15zdnd11an1n64x5 FILLER_378_264 ();
 b15zdnd11an1n64x5 FILLER_378_328 ();
 b15zdnd11an1n64x5 FILLER_378_392 ();
 b15zdnd11an1n64x5 FILLER_378_456 ();
 b15zdnd11an1n64x5 FILLER_378_520 ();
 b15zdnd11an1n64x5 FILLER_378_584 ();
 b15zdnd11an1n64x5 FILLER_378_648 ();
 b15zdnd11an1n04x5 FILLER_378_712 ();
 b15zdnd00an1n02x5 FILLER_378_716 ();
 b15zdnd11an1n64x5 FILLER_378_726 ();
 b15zdnd11an1n64x5 FILLER_378_790 ();
 b15zdnd11an1n64x5 FILLER_378_854 ();
 b15zdnd11an1n64x5 FILLER_378_918 ();
 b15zdnd11an1n64x5 FILLER_378_982 ();
 b15zdnd11an1n64x5 FILLER_378_1046 ();
 b15zdnd11an1n64x5 FILLER_378_1110 ();
 b15zdnd11an1n64x5 FILLER_378_1174 ();
 b15zdnd11an1n64x5 FILLER_378_1238 ();
 b15zdnd11an1n64x5 FILLER_378_1302 ();
 b15zdnd11an1n64x5 FILLER_378_1366 ();
 b15zdnd11an1n64x5 FILLER_378_1430 ();
 b15zdnd11an1n64x5 FILLER_378_1494 ();
 b15zdnd11an1n64x5 FILLER_378_1558 ();
 b15zdnd11an1n64x5 FILLER_378_1622 ();
 b15zdnd11an1n64x5 FILLER_378_1686 ();
 b15zdnd11an1n64x5 FILLER_378_1750 ();
 b15zdnd11an1n64x5 FILLER_378_1814 ();
 b15zdnd11an1n64x5 FILLER_378_1878 ();
 b15zdnd11an1n64x5 FILLER_378_1942 ();
 b15zdnd11an1n64x5 FILLER_378_2006 ();
 b15zdnd11an1n64x5 FILLER_378_2070 ();
 b15zdnd11an1n16x5 FILLER_378_2134 ();
 b15zdnd11an1n04x5 FILLER_378_2150 ();
 b15zdnd11an1n64x5 FILLER_378_2162 ();
 b15zdnd11an1n32x5 FILLER_378_2226 ();
 b15zdnd11an1n16x5 FILLER_378_2258 ();
 b15zdnd00an1n02x5 FILLER_378_2274 ();
 b15zdnd11an1n64x5 FILLER_379_0 ();
 b15zdnd11an1n64x5 FILLER_379_64 ();
 b15zdnd11an1n64x5 FILLER_379_128 ();
 b15zdnd11an1n64x5 FILLER_379_192 ();
 b15zdnd11an1n64x5 FILLER_379_256 ();
 b15zdnd11an1n64x5 FILLER_379_320 ();
 b15zdnd11an1n64x5 FILLER_379_384 ();
 b15zdnd11an1n64x5 FILLER_379_448 ();
 b15zdnd11an1n64x5 FILLER_379_512 ();
 b15zdnd11an1n64x5 FILLER_379_576 ();
 b15zdnd11an1n64x5 FILLER_379_640 ();
 b15zdnd11an1n64x5 FILLER_379_704 ();
 b15zdnd11an1n64x5 FILLER_379_768 ();
 b15zdnd11an1n64x5 FILLER_379_832 ();
 b15zdnd11an1n64x5 FILLER_379_896 ();
 b15zdnd11an1n64x5 FILLER_379_960 ();
 b15zdnd11an1n64x5 FILLER_379_1024 ();
 b15zdnd11an1n64x5 FILLER_379_1088 ();
 b15zdnd11an1n64x5 FILLER_379_1152 ();
 b15zdnd11an1n64x5 FILLER_379_1216 ();
 b15zdnd11an1n64x5 FILLER_379_1280 ();
 b15zdnd11an1n64x5 FILLER_379_1344 ();
 b15zdnd11an1n64x5 FILLER_379_1408 ();
 b15zdnd11an1n64x5 FILLER_379_1472 ();
 b15zdnd11an1n64x5 FILLER_379_1536 ();
 b15zdnd11an1n64x5 FILLER_379_1600 ();
 b15zdnd11an1n64x5 FILLER_379_1664 ();
 b15zdnd11an1n64x5 FILLER_379_1728 ();
 b15zdnd11an1n64x5 FILLER_379_1792 ();
 b15zdnd11an1n64x5 FILLER_379_1856 ();
 b15zdnd11an1n64x5 FILLER_379_1920 ();
 b15zdnd11an1n64x5 FILLER_379_1984 ();
 b15zdnd11an1n64x5 FILLER_379_2048 ();
 b15zdnd11an1n64x5 FILLER_379_2112 ();
 b15zdnd11an1n64x5 FILLER_379_2176 ();
 b15zdnd11an1n32x5 FILLER_379_2240 ();
 b15zdnd11an1n08x5 FILLER_379_2272 ();
 b15zdnd11an1n04x5 FILLER_379_2280 ();
 b15zdnd11an1n64x5 FILLER_380_8 ();
 b15zdnd11an1n64x5 FILLER_380_72 ();
 b15zdnd11an1n64x5 FILLER_380_136 ();
 b15zdnd11an1n64x5 FILLER_380_200 ();
 b15zdnd11an1n64x5 FILLER_380_264 ();
 b15zdnd11an1n64x5 FILLER_380_328 ();
 b15zdnd11an1n64x5 FILLER_380_392 ();
 b15zdnd11an1n64x5 FILLER_380_456 ();
 b15zdnd11an1n64x5 FILLER_380_520 ();
 b15zdnd11an1n64x5 FILLER_380_584 ();
 b15zdnd11an1n64x5 FILLER_380_648 ();
 b15zdnd11an1n04x5 FILLER_380_712 ();
 b15zdnd00an1n02x5 FILLER_380_716 ();
 b15zdnd11an1n64x5 FILLER_380_726 ();
 b15zdnd11an1n64x5 FILLER_380_790 ();
 b15zdnd11an1n64x5 FILLER_380_854 ();
 b15zdnd11an1n64x5 FILLER_380_918 ();
 b15zdnd11an1n64x5 FILLER_380_982 ();
 b15zdnd11an1n64x5 FILLER_380_1046 ();
 b15zdnd11an1n64x5 FILLER_380_1110 ();
 b15zdnd11an1n64x5 FILLER_380_1174 ();
 b15zdnd11an1n64x5 FILLER_380_1238 ();
 b15zdnd11an1n64x5 FILLER_380_1302 ();
 b15zdnd11an1n64x5 FILLER_380_1366 ();
 b15zdnd11an1n64x5 FILLER_380_1430 ();
 b15zdnd11an1n64x5 FILLER_380_1494 ();
 b15zdnd11an1n64x5 FILLER_380_1558 ();
 b15zdnd11an1n64x5 FILLER_380_1622 ();
 b15zdnd11an1n64x5 FILLER_380_1686 ();
 b15zdnd11an1n64x5 FILLER_380_1750 ();
 b15zdnd11an1n64x5 FILLER_380_1814 ();
 b15zdnd11an1n64x5 FILLER_380_1878 ();
 b15zdnd11an1n64x5 FILLER_380_1942 ();
 b15zdnd11an1n64x5 FILLER_380_2006 ();
 b15zdnd11an1n64x5 FILLER_380_2070 ();
 b15zdnd11an1n16x5 FILLER_380_2134 ();
 b15zdnd11an1n04x5 FILLER_380_2150 ();
 b15zdnd11an1n64x5 FILLER_380_2162 ();
 b15zdnd11an1n32x5 FILLER_380_2226 ();
 b15zdnd11an1n16x5 FILLER_380_2258 ();
 b15zdnd00an1n02x5 FILLER_380_2274 ();
 b15zdnd11an1n64x5 FILLER_381_0 ();
 b15zdnd11an1n64x5 FILLER_381_64 ();
 b15zdnd11an1n64x5 FILLER_381_128 ();
 b15zdnd11an1n64x5 FILLER_381_192 ();
 b15zdnd11an1n64x5 FILLER_381_256 ();
 b15zdnd11an1n64x5 FILLER_381_320 ();
 b15zdnd11an1n64x5 FILLER_381_384 ();
 b15zdnd11an1n64x5 FILLER_381_448 ();
 b15zdnd11an1n64x5 FILLER_381_512 ();
 b15zdnd11an1n64x5 FILLER_381_576 ();
 b15zdnd11an1n64x5 FILLER_381_640 ();
 b15zdnd11an1n64x5 FILLER_381_704 ();
 b15zdnd11an1n64x5 FILLER_381_768 ();
 b15zdnd11an1n64x5 FILLER_381_832 ();
 b15zdnd11an1n64x5 FILLER_381_896 ();
 b15zdnd11an1n64x5 FILLER_381_960 ();
 b15zdnd11an1n64x5 FILLER_381_1024 ();
 b15zdnd11an1n64x5 FILLER_381_1088 ();
 b15zdnd11an1n64x5 FILLER_381_1152 ();
 b15zdnd11an1n64x5 FILLER_381_1216 ();
 b15zdnd11an1n64x5 FILLER_381_1280 ();
 b15zdnd11an1n64x5 FILLER_381_1344 ();
 b15zdnd11an1n64x5 FILLER_381_1408 ();
 b15zdnd11an1n64x5 FILLER_381_1472 ();
 b15zdnd11an1n64x5 FILLER_381_1536 ();
 b15zdnd11an1n64x5 FILLER_381_1600 ();
 b15zdnd11an1n64x5 FILLER_381_1664 ();
 b15zdnd11an1n64x5 FILLER_381_1728 ();
 b15zdnd11an1n64x5 FILLER_381_1792 ();
 b15zdnd11an1n64x5 FILLER_381_1856 ();
 b15zdnd11an1n64x5 FILLER_381_1920 ();
 b15zdnd11an1n64x5 FILLER_381_1984 ();
 b15zdnd11an1n64x5 FILLER_381_2048 ();
 b15zdnd11an1n64x5 FILLER_381_2112 ();
 b15zdnd11an1n64x5 FILLER_381_2176 ();
 b15zdnd11an1n32x5 FILLER_381_2240 ();
 b15zdnd11an1n08x5 FILLER_381_2272 ();
 b15zdnd11an1n04x5 FILLER_381_2280 ();
 b15zdnd11an1n64x5 FILLER_382_8 ();
 b15zdnd11an1n64x5 FILLER_382_72 ();
 b15zdnd11an1n64x5 FILLER_382_136 ();
 b15zdnd11an1n64x5 FILLER_382_200 ();
 b15zdnd11an1n64x5 FILLER_382_264 ();
 b15zdnd11an1n64x5 FILLER_382_328 ();
 b15zdnd11an1n64x5 FILLER_382_392 ();
 b15zdnd11an1n64x5 FILLER_382_456 ();
 b15zdnd11an1n64x5 FILLER_382_520 ();
 b15zdnd11an1n64x5 FILLER_382_584 ();
 b15zdnd11an1n64x5 FILLER_382_648 ();
 b15zdnd11an1n04x5 FILLER_382_712 ();
 b15zdnd00an1n02x5 FILLER_382_716 ();
 b15zdnd11an1n64x5 FILLER_382_726 ();
 b15zdnd11an1n64x5 FILLER_382_790 ();
 b15zdnd11an1n64x5 FILLER_382_854 ();
 b15zdnd11an1n64x5 FILLER_382_918 ();
 b15zdnd11an1n64x5 FILLER_382_982 ();
 b15zdnd11an1n64x5 FILLER_382_1046 ();
 b15zdnd11an1n64x5 FILLER_382_1110 ();
 b15zdnd11an1n64x5 FILLER_382_1174 ();
 b15zdnd11an1n64x5 FILLER_382_1238 ();
 b15zdnd11an1n64x5 FILLER_382_1302 ();
 b15zdnd11an1n64x5 FILLER_382_1366 ();
 b15zdnd11an1n64x5 FILLER_382_1430 ();
 b15zdnd11an1n64x5 FILLER_382_1494 ();
 b15zdnd11an1n64x5 FILLER_382_1558 ();
 b15zdnd11an1n64x5 FILLER_382_1622 ();
 b15zdnd11an1n64x5 FILLER_382_1686 ();
 b15zdnd11an1n64x5 FILLER_382_1750 ();
 b15zdnd11an1n64x5 FILLER_382_1814 ();
 b15zdnd11an1n64x5 FILLER_382_1878 ();
 b15zdnd11an1n64x5 FILLER_382_1942 ();
 b15zdnd11an1n64x5 FILLER_382_2006 ();
 b15zdnd11an1n64x5 FILLER_382_2070 ();
 b15zdnd11an1n16x5 FILLER_382_2134 ();
 b15zdnd11an1n04x5 FILLER_382_2150 ();
 b15zdnd11an1n64x5 FILLER_382_2162 ();
 b15zdnd11an1n32x5 FILLER_382_2226 ();
 b15zdnd11an1n16x5 FILLER_382_2258 ();
 b15zdnd00an1n02x5 FILLER_382_2274 ();
 b15zdnd11an1n64x5 FILLER_383_0 ();
 b15zdnd11an1n64x5 FILLER_383_64 ();
 b15zdnd11an1n64x5 FILLER_383_128 ();
 b15zdnd11an1n64x5 FILLER_383_192 ();
 b15zdnd11an1n64x5 FILLER_383_256 ();
 b15zdnd11an1n64x5 FILLER_383_320 ();
 b15zdnd11an1n64x5 FILLER_383_384 ();
 b15zdnd11an1n64x5 FILLER_383_448 ();
 b15zdnd11an1n64x5 FILLER_383_512 ();
 b15zdnd11an1n64x5 FILLER_383_576 ();
 b15zdnd11an1n64x5 FILLER_383_640 ();
 b15zdnd11an1n64x5 FILLER_383_704 ();
 b15zdnd11an1n64x5 FILLER_383_768 ();
 b15zdnd11an1n64x5 FILLER_383_832 ();
 b15zdnd11an1n64x5 FILLER_383_896 ();
 b15zdnd11an1n64x5 FILLER_383_960 ();
 b15zdnd11an1n64x5 FILLER_383_1024 ();
 b15zdnd11an1n64x5 FILLER_383_1088 ();
 b15zdnd11an1n64x5 FILLER_383_1152 ();
 b15zdnd11an1n64x5 FILLER_383_1216 ();
 b15zdnd11an1n64x5 FILLER_383_1280 ();
 b15zdnd11an1n64x5 FILLER_383_1344 ();
 b15zdnd11an1n64x5 FILLER_383_1408 ();
 b15zdnd11an1n64x5 FILLER_383_1472 ();
 b15zdnd11an1n64x5 FILLER_383_1536 ();
 b15zdnd11an1n64x5 FILLER_383_1600 ();
 b15zdnd11an1n64x5 FILLER_383_1664 ();
 b15zdnd11an1n64x5 FILLER_383_1728 ();
 b15zdnd11an1n64x5 FILLER_383_1792 ();
 b15zdnd11an1n64x5 FILLER_383_1856 ();
 b15zdnd11an1n64x5 FILLER_383_1920 ();
 b15zdnd11an1n64x5 FILLER_383_1984 ();
 b15zdnd11an1n64x5 FILLER_383_2048 ();
 b15zdnd11an1n64x5 FILLER_383_2112 ();
 b15zdnd11an1n64x5 FILLER_383_2176 ();
 b15zdnd11an1n32x5 FILLER_383_2240 ();
 b15zdnd11an1n08x5 FILLER_383_2272 ();
 b15zdnd11an1n04x5 FILLER_383_2280 ();
 b15zdnd11an1n64x5 FILLER_384_8 ();
 b15zdnd11an1n64x5 FILLER_384_72 ();
 b15zdnd11an1n64x5 FILLER_384_136 ();
 b15zdnd11an1n64x5 FILLER_384_200 ();
 b15zdnd11an1n64x5 FILLER_384_264 ();
 b15zdnd11an1n64x5 FILLER_384_328 ();
 b15zdnd11an1n64x5 FILLER_384_392 ();
 b15zdnd11an1n64x5 FILLER_384_456 ();
 b15zdnd11an1n64x5 FILLER_384_520 ();
 b15zdnd11an1n64x5 FILLER_384_584 ();
 b15zdnd11an1n64x5 FILLER_384_648 ();
 b15zdnd11an1n04x5 FILLER_384_712 ();
 b15zdnd00an1n02x5 FILLER_384_716 ();
 b15zdnd11an1n64x5 FILLER_384_726 ();
 b15zdnd11an1n64x5 FILLER_384_790 ();
 b15zdnd11an1n64x5 FILLER_384_854 ();
 b15zdnd11an1n64x5 FILLER_384_918 ();
 b15zdnd11an1n64x5 FILLER_384_982 ();
 b15zdnd11an1n64x5 FILLER_384_1046 ();
 b15zdnd11an1n64x5 FILLER_384_1110 ();
 b15zdnd11an1n64x5 FILLER_384_1174 ();
 b15zdnd11an1n64x5 FILLER_384_1238 ();
 b15zdnd11an1n64x5 FILLER_384_1302 ();
 b15zdnd11an1n64x5 FILLER_384_1366 ();
 b15zdnd11an1n64x5 FILLER_384_1430 ();
 b15zdnd11an1n64x5 FILLER_384_1494 ();
 b15zdnd11an1n64x5 FILLER_384_1558 ();
 b15zdnd11an1n64x5 FILLER_384_1622 ();
 b15zdnd11an1n64x5 FILLER_384_1686 ();
 b15zdnd11an1n64x5 FILLER_384_1750 ();
 b15zdnd11an1n64x5 FILLER_384_1814 ();
 b15zdnd11an1n64x5 FILLER_384_1878 ();
 b15zdnd11an1n64x5 FILLER_384_1942 ();
 b15zdnd11an1n64x5 FILLER_384_2006 ();
 b15zdnd11an1n64x5 FILLER_384_2070 ();
 b15zdnd11an1n16x5 FILLER_384_2134 ();
 b15zdnd11an1n04x5 FILLER_384_2150 ();
 b15zdnd11an1n64x5 FILLER_384_2162 ();
 b15zdnd11an1n32x5 FILLER_384_2226 ();
 b15zdnd11an1n16x5 FILLER_384_2258 ();
 b15zdnd00an1n02x5 FILLER_384_2274 ();
 b15zdnd11an1n64x5 FILLER_385_0 ();
 b15zdnd11an1n64x5 FILLER_385_64 ();
 b15zdnd11an1n64x5 FILLER_385_128 ();
 b15zdnd11an1n64x5 FILLER_385_192 ();
 b15zdnd11an1n64x5 FILLER_385_256 ();
 b15zdnd11an1n64x5 FILLER_385_320 ();
 b15zdnd11an1n64x5 FILLER_385_384 ();
 b15zdnd11an1n64x5 FILLER_385_448 ();
 b15zdnd11an1n64x5 FILLER_385_512 ();
 b15zdnd11an1n64x5 FILLER_385_576 ();
 b15zdnd11an1n64x5 FILLER_385_640 ();
 b15zdnd11an1n64x5 FILLER_385_704 ();
 b15zdnd11an1n64x5 FILLER_385_768 ();
 b15zdnd11an1n64x5 FILLER_385_832 ();
 b15zdnd11an1n64x5 FILLER_385_896 ();
 b15zdnd11an1n64x5 FILLER_385_960 ();
 b15zdnd11an1n64x5 FILLER_385_1024 ();
 b15zdnd11an1n64x5 FILLER_385_1088 ();
 b15zdnd11an1n64x5 FILLER_385_1152 ();
 b15zdnd11an1n64x5 FILLER_385_1216 ();
 b15zdnd11an1n64x5 FILLER_385_1280 ();
 b15zdnd11an1n64x5 FILLER_385_1344 ();
 b15zdnd11an1n64x5 FILLER_385_1408 ();
 b15zdnd11an1n64x5 FILLER_385_1472 ();
 b15zdnd11an1n64x5 FILLER_385_1536 ();
 b15zdnd11an1n64x5 FILLER_385_1600 ();
 b15zdnd11an1n64x5 FILLER_385_1664 ();
 b15zdnd11an1n64x5 FILLER_385_1728 ();
 b15zdnd11an1n64x5 FILLER_385_1792 ();
 b15zdnd11an1n64x5 FILLER_385_1856 ();
 b15zdnd11an1n64x5 FILLER_385_1920 ();
 b15zdnd11an1n64x5 FILLER_385_1984 ();
 b15zdnd11an1n64x5 FILLER_385_2048 ();
 b15zdnd11an1n64x5 FILLER_385_2112 ();
 b15zdnd11an1n64x5 FILLER_385_2176 ();
 b15zdnd11an1n32x5 FILLER_385_2240 ();
 b15zdnd11an1n08x5 FILLER_385_2272 ();
 b15zdnd11an1n04x5 FILLER_385_2280 ();
 b15zdnd11an1n64x5 FILLER_386_8 ();
 b15zdnd11an1n64x5 FILLER_386_72 ();
 b15zdnd11an1n64x5 FILLER_386_136 ();
 b15zdnd11an1n64x5 FILLER_386_200 ();
 b15zdnd11an1n64x5 FILLER_386_264 ();
 b15zdnd11an1n64x5 FILLER_386_328 ();
 b15zdnd11an1n64x5 FILLER_386_392 ();
 b15zdnd11an1n64x5 FILLER_386_456 ();
 b15zdnd11an1n64x5 FILLER_386_520 ();
 b15zdnd11an1n64x5 FILLER_386_584 ();
 b15zdnd11an1n64x5 FILLER_386_648 ();
 b15zdnd11an1n04x5 FILLER_386_712 ();
 b15zdnd00an1n02x5 FILLER_386_716 ();
 b15zdnd11an1n64x5 FILLER_386_726 ();
 b15zdnd11an1n64x5 FILLER_386_790 ();
 b15zdnd11an1n64x5 FILLER_386_854 ();
 b15zdnd11an1n64x5 FILLER_386_918 ();
 b15zdnd11an1n64x5 FILLER_386_982 ();
 b15zdnd11an1n64x5 FILLER_386_1046 ();
 b15zdnd11an1n64x5 FILLER_386_1110 ();
 b15zdnd11an1n64x5 FILLER_386_1174 ();
 b15zdnd11an1n64x5 FILLER_386_1238 ();
 b15zdnd11an1n64x5 FILLER_386_1302 ();
 b15zdnd11an1n64x5 FILLER_386_1366 ();
 b15zdnd11an1n64x5 FILLER_386_1430 ();
 b15zdnd11an1n64x5 FILLER_386_1494 ();
 b15zdnd11an1n64x5 FILLER_386_1558 ();
 b15zdnd11an1n64x5 FILLER_386_1622 ();
 b15zdnd11an1n64x5 FILLER_386_1686 ();
 b15zdnd11an1n64x5 FILLER_386_1750 ();
 b15zdnd11an1n64x5 FILLER_386_1814 ();
 b15zdnd11an1n64x5 FILLER_386_1878 ();
 b15zdnd11an1n64x5 FILLER_386_1942 ();
 b15zdnd11an1n64x5 FILLER_386_2006 ();
 b15zdnd11an1n64x5 FILLER_386_2070 ();
 b15zdnd11an1n16x5 FILLER_386_2134 ();
 b15zdnd11an1n04x5 FILLER_386_2150 ();
 b15zdnd11an1n64x5 FILLER_386_2162 ();
 b15zdnd11an1n32x5 FILLER_386_2226 ();
 b15zdnd11an1n16x5 FILLER_386_2258 ();
 b15zdnd00an1n02x5 FILLER_386_2274 ();
 b15zdnd11an1n64x5 FILLER_387_0 ();
 b15zdnd11an1n64x5 FILLER_387_64 ();
 b15zdnd11an1n64x5 FILLER_387_128 ();
 b15zdnd11an1n64x5 FILLER_387_192 ();
 b15zdnd11an1n64x5 FILLER_387_256 ();
 b15zdnd11an1n64x5 FILLER_387_320 ();
 b15zdnd11an1n64x5 FILLER_387_384 ();
 b15zdnd11an1n64x5 FILLER_387_448 ();
 b15zdnd11an1n64x5 FILLER_387_512 ();
 b15zdnd11an1n64x5 FILLER_387_576 ();
 b15zdnd11an1n64x5 FILLER_387_640 ();
 b15zdnd11an1n64x5 FILLER_387_704 ();
 b15zdnd11an1n64x5 FILLER_387_768 ();
 b15zdnd11an1n64x5 FILLER_387_832 ();
 b15zdnd11an1n64x5 FILLER_387_896 ();
 b15zdnd11an1n04x5 FILLER_387_960 ();
 b15zdnd00an1n01x5 FILLER_387_964 ();
 b15zdnd11an1n64x5 FILLER_387_969 ();
 b15zdnd11an1n64x5 FILLER_387_1033 ();
 b15zdnd11an1n64x5 FILLER_387_1097 ();
 b15zdnd11an1n64x5 FILLER_387_1161 ();
 b15zdnd11an1n64x5 FILLER_387_1225 ();
 b15zdnd11an1n64x5 FILLER_387_1289 ();
 b15zdnd11an1n64x5 FILLER_387_1353 ();
 b15zdnd11an1n64x5 FILLER_387_1417 ();
 b15zdnd11an1n64x5 FILLER_387_1481 ();
 b15zdnd11an1n64x5 FILLER_387_1545 ();
 b15zdnd11an1n64x5 FILLER_387_1609 ();
 b15zdnd11an1n64x5 FILLER_387_1673 ();
 b15zdnd11an1n64x5 FILLER_387_1737 ();
 b15zdnd11an1n64x5 FILLER_387_1801 ();
 b15zdnd11an1n64x5 FILLER_387_1865 ();
 b15zdnd11an1n64x5 FILLER_387_1929 ();
 b15zdnd11an1n64x5 FILLER_387_1993 ();
 b15zdnd11an1n64x5 FILLER_387_2057 ();
 b15zdnd11an1n64x5 FILLER_387_2121 ();
 b15zdnd11an1n64x5 FILLER_387_2185 ();
 b15zdnd11an1n32x5 FILLER_387_2249 ();
 b15zdnd00an1n02x5 FILLER_387_2281 ();
 b15zdnd00an1n01x5 FILLER_387_2283 ();
 b15zdnd11an1n64x5 FILLER_388_8 ();
 b15zdnd11an1n64x5 FILLER_388_72 ();
 b15zdnd11an1n64x5 FILLER_388_136 ();
 b15zdnd11an1n64x5 FILLER_388_200 ();
 b15zdnd11an1n64x5 FILLER_388_264 ();
 b15zdnd11an1n64x5 FILLER_388_328 ();
 b15zdnd11an1n64x5 FILLER_388_392 ();
 b15zdnd11an1n64x5 FILLER_388_456 ();
 b15zdnd11an1n64x5 FILLER_388_520 ();
 b15zdnd11an1n64x5 FILLER_388_584 ();
 b15zdnd11an1n64x5 FILLER_388_648 ();
 b15zdnd11an1n04x5 FILLER_388_712 ();
 b15zdnd00an1n02x5 FILLER_388_716 ();
 b15zdnd11an1n64x5 FILLER_388_726 ();
 b15zdnd11an1n32x5 FILLER_388_790 ();
 b15zdnd11an1n16x5 FILLER_388_822 ();
 b15zdnd11an1n08x5 FILLER_388_838 ();
 b15zdnd00an1n02x5 FILLER_388_846 ();
 b15zdnd11an1n08x5 FILLER_388_852 ();
 b15zdnd11an1n64x5 FILLER_388_902 ();
 b15zdnd00an1n02x5 FILLER_388_966 ();
 b15zdnd00an1n01x5 FILLER_388_968 ();
 b15zdnd11an1n64x5 FILLER_388_973 ();
 b15zdnd11an1n64x5 FILLER_388_1037 ();
 b15zdnd11an1n64x5 FILLER_388_1101 ();
 b15zdnd11an1n64x5 FILLER_388_1165 ();
 b15zdnd11an1n64x5 FILLER_388_1229 ();
 b15zdnd11an1n32x5 FILLER_388_1293 ();
 b15zdnd00an1n02x5 FILLER_388_1325 ();
 b15zdnd00an1n01x5 FILLER_388_1327 ();
 b15zdnd11an1n64x5 FILLER_388_1332 ();
 b15zdnd11an1n64x5 FILLER_388_1396 ();
 b15zdnd11an1n64x5 FILLER_388_1460 ();
 b15zdnd11an1n64x5 FILLER_388_1524 ();
 b15zdnd11an1n64x5 FILLER_388_1588 ();
 b15zdnd11an1n64x5 FILLER_388_1652 ();
 b15zdnd11an1n64x5 FILLER_388_1716 ();
 b15zdnd11an1n64x5 FILLER_388_1780 ();
 b15zdnd11an1n64x5 FILLER_388_1844 ();
 b15zdnd11an1n64x5 FILLER_388_1908 ();
 b15zdnd11an1n64x5 FILLER_388_1972 ();
 b15zdnd11an1n64x5 FILLER_388_2036 ();
 b15zdnd11an1n32x5 FILLER_388_2100 ();
 b15zdnd11an1n16x5 FILLER_388_2132 ();
 b15zdnd11an1n04x5 FILLER_388_2148 ();
 b15zdnd00an1n02x5 FILLER_388_2152 ();
 b15zdnd11an1n64x5 FILLER_388_2162 ();
 b15zdnd11an1n32x5 FILLER_388_2226 ();
 b15zdnd11an1n16x5 FILLER_388_2258 ();
 b15zdnd00an1n02x5 FILLER_388_2274 ();
 b15zdnd11an1n64x5 FILLER_389_0 ();
 b15zdnd11an1n64x5 FILLER_389_64 ();
 b15zdnd11an1n64x5 FILLER_389_128 ();
 b15zdnd11an1n64x5 FILLER_389_192 ();
 b15zdnd11an1n64x5 FILLER_389_256 ();
 b15zdnd11an1n64x5 FILLER_389_320 ();
 b15zdnd11an1n64x5 FILLER_389_384 ();
 b15zdnd11an1n64x5 FILLER_389_448 ();
 b15zdnd11an1n64x5 FILLER_389_512 ();
 b15zdnd11an1n64x5 FILLER_389_576 ();
 b15zdnd11an1n64x5 FILLER_389_640 ();
 b15zdnd11an1n64x5 FILLER_389_704 ();
 b15zdnd11an1n16x5 FILLER_389_768 ();
 b15zdnd11an1n04x5 FILLER_389_784 ();
 b15zdnd00an1n02x5 FILLER_389_788 ();
 b15zdnd11an1n32x5 FILLER_389_794 ();
 b15zdnd11an1n16x5 FILLER_389_826 ();
 b15zdnd11an1n04x5 FILLER_389_842 ();
 b15zdnd00an1n02x5 FILLER_389_846 ();
 b15zdnd00an1n01x5 FILLER_389_848 ();
 b15zdnd11an1n04x5 FILLER_389_853 ();
 b15zdnd11an1n04x5 FILLER_389_861 ();
 b15zdnd11an1n32x5 FILLER_389_907 ();
 b15zdnd11an1n16x5 FILLER_389_939 ();
 b15zdnd11an1n04x5 FILLER_389_955 ();
 b15zdnd00an1n02x5 FILLER_389_959 ();
 b15zdnd11an1n04x5 FILLER_389_965 ();
 b15zdnd00an1n01x5 FILLER_389_969 ();
 b15zdnd11an1n64x5 FILLER_389_1012 ();
 b15zdnd11an1n64x5 FILLER_389_1076 ();
 b15zdnd11an1n64x5 FILLER_389_1140 ();
 b15zdnd11an1n64x5 FILLER_389_1204 ();
 b15zdnd11an1n32x5 FILLER_389_1268 ();
 b15zdnd00an1n02x5 FILLER_389_1300 ();
 b15zdnd11an1n04x5 FILLER_389_1306 ();
 b15zdnd11an1n64x5 FILLER_389_1352 ();
 b15zdnd11an1n64x5 FILLER_389_1416 ();
 b15zdnd11an1n64x5 FILLER_389_1480 ();
 b15zdnd11an1n64x5 FILLER_389_1544 ();
 b15zdnd11an1n64x5 FILLER_389_1608 ();
 b15zdnd11an1n64x5 FILLER_389_1672 ();
 b15zdnd11an1n64x5 FILLER_389_1736 ();
 b15zdnd11an1n64x5 FILLER_389_1800 ();
 b15zdnd11an1n64x5 FILLER_389_1864 ();
 b15zdnd11an1n64x5 FILLER_389_1928 ();
 b15zdnd11an1n64x5 FILLER_389_1992 ();
 b15zdnd11an1n64x5 FILLER_389_2056 ();
 b15zdnd11an1n64x5 FILLER_389_2120 ();
 b15zdnd11an1n64x5 FILLER_389_2184 ();
 b15zdnd11an1n32x5 FILLER_389_2248 ();
 b15zdnd11an1n04x5 FILLER_389_2280 ();
endmodule
