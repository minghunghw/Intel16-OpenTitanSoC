VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
	 DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.0005 ;

MACRO ringpll
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN ringpll 0 0 ;
  SIZE 201.96 BY 413.28 ;
  SYMMETRY X Y ;
  PIN fz_vcotrim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 222.908 0.292 222.952 ;
    END
  END fz_vcotrim[3]
  PIN fz_vcotrim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 223.088 0.292 223.132 ;
    END
  END fz_vcotrim[1]
  PIN fz_vcotrim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 222.278 0.292 222.322 ;
    END
  END fz_vcotrim[4]
  PIN fz_vcotrim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 221.828 0.292 221.872 ;
    END
  END fz_vcotrim[5]
  PIN fz_vcotrim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 221.648 0.292 221.692 ;
    END
  END fz_vcotrim[6]
  PIN fz_vcotrim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 221.198 0.292 221.242 ;
    END
  END fz_vcotrim[7]
  PIN fz_vcotrim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 221.018 0.292 221.062 ;
    END
  END fz_vcotrim[8]
  PIN fz_vcotrim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 220.568 0.292 220.612 ;
    END
  END fz_vcotrim[9]
  PIN fz_vcotrim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 219.938 0.292 219.982 ;
    END
  END fz_vcotrim[10]
  PIN fz_vcosel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 224.168 0.292 224.212 ;
    END
  END fz_vcosel
  PIN fz_tight_loopb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 223.718 0.292 223.762 ;
    END
  END fz_tight_loopb
  PIN fz_startup[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 225.608 0.292 225.652 ;
    END
  END fz_startup[0]
  PIN fz_startup[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 226.058 0.292 226.102 ;
    END
  END fz_startup[1]
  PIN fz_startup[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 225.428 0.292 225.472 ;
    END
  END fz_startup[3]
  PIN fz_startup[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 224.348 0.292 224.392 ;
    END
  END fz_startup[4]
  PIN fz_startup[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 224.798 0.292 224.842 ;
    END
  END fz_startup[5]
  PIN fz_startup[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 224.978 0.292 225.022 ;
    END
  END fz_startup[2]
  PIN fz_spare[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 226.868 0.292 226.912 ;
    END
  END fz_spare[1]
  PIN fz_spare[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 227.318 0.292 227.362 ;
    END
  END fz_spare[2]
  PIN fz_spare[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 226.238 0.292 226.282 ;
    END
  END fz_spare[3]
  PIN fz_spare[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 226.688 0.292 226.732 ;
    END
  END fz_spare[4]
  PIN fz_spare[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 227.498 0.292 227.542 ;
    END
  END fz_spare[0]
  PIN fz_skadj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 228.758 0.292 228.802 ;
    END
  END fz_skadj[0]
  PIN fz_skadj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 229.208 0.292 229.252 ;
    END
  END fz_skadj[1]
  PIN fz_skadj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 228.128 0.292 228.172 ;
    END
  END fz_skadj[2]
  PIN fz_skadj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 227.948 0.292 227.992 ;
    END
  END fz_skadj[4]
  PIN fz_pfddly[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 229.838 0.292 229.882 ;
    END
  END fz_pfddly[0]
  PIN fz_pfddly[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 229.388 0.292 229.432 ;
    END
  END fz_pfddly[1]
  PIN fz_pfd_pw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 230.648 0.292 230.692 ;
    END
  END fz_pfd_pw[0]
  PIN fz_pfd_pw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 230.468 0.292 230.512 ;
    END
  END fz_pfd_pw[1]
  PIN fz_pfd_pw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 230.018 0.292 230.062 ;
    END
  END fz_pfd_pw[2]
  PIN fz_skadj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 228.578 0.292 228.622 ;
    END
  END fz_skadj[3]
  PIN fz_nopfdpwrgate
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 231.098 0.292 231.142 ;
    END
  END fz_nopfdpwrgate
  PIN fz_lpfclksel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 231.728 0.292 231.772 ;
    END
  END fz_lpfclksel
  PIN fz_lockthresh[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 232.358 0.292 232.402 ;
    END
  END fz_lockthresh[1]
  PIN fz_lockthresh[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 231.908 0.292 231.952 ;
    END
  END fz_lockthresh[2]
  PIN fz_lockthresh[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 231.278 0.292 231.322 ;
    END
  END fz_lockthresh[3]
  PIN fz_lockstickyb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 232.538 0.292 232.582 ;
    END
  END fz_lockstickyb
  PIN fz_lockforce
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 233.168 0.292 233.212 ;
    END
  END fz_lockforce
  PIN fz_lockcnt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 234.248 0.292 234.292 ;
    END
  END fz_lockcnt[0]
  PIN fz_lockcnt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 233.798 0.292 233.842 ;
    END
  END fz_lockcnt[1]
  PIN fz_lockcnt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 233.618 0.292 233.662 ;
    END
  END fz_lockcnt[2]
  PIN fz_irefgen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 235.688 0.292 235.732 ;
    END
  END fz_irefgen[0]
  PIN fz_irefgen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 235.058 0.292 235.102 ;
    END
  END fz_irefgen[1]
  PIN fz_irefgen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 235.508 0.292 235.552 ;
    END
  END fz_irefgen[2]
  PIN fz_irefgen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 234.878 0.292 234.922 ;
    END
  END fz_irefgen[3]
  PIN fz_irefgen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 234.428 0.292 234.472 ;
    END
  END fz_irefgen[4]
  PIN fz_dca_ctrl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 238.028 0.292 238.072 ;
    END
  END fz_dca_ctrl[0]
  PIN fz_dca_ctrl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 237.398 0.292 237.442 ;
    END
  END fz_dca_ctrl[1]
  PIN fz_dca_ctrl[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 236.948 0.292 236.992 ;
    END
  END fz_dca_ctrl[2]
  PIN fz_dca_ctrl[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 236.318 0.292 236.362 ;
    END
  END fz_dca_ctrl[3]
  PIN fz_dca_ctrl[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 236.768 0.292 236.812 ;
    END
  END fz_dca_ctrl[4]
  PIN fz_dca_ctrl[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 236.138 0.292 236.182 ;
    END
  END fz_dca_ctrl[5]
  PIN fz_dca_cb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 237.578 0.292 237.622 ;
    END
  END fz_dca_cb[1]
  PIN fz_lockthresh[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 232.988 0.292 233.032 ;
    END
  END fz_lockthresh[0]
  PIN fz_cpnbias[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 239.288 0.292 239.332 ;
    END
  END fz_cpnbias[0]
  PIN fz_cpnbias[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 238.658 0.292 238.702 ;
    END
  END fz_cpnbias[1]
  PIN fz_cp2trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 240.548 0.292 240.592 ;
    END
  END fz_cp2trim[0]
  PIN fz_dca_cb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 238.208 0.292 238.252 ;
    END
  END fz_dca_cb[0]
  PIN fz_cp2trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 240.098 0.292 240.142 ;
    END
  END fz_cp2trim[1]
  PIN fz_cp2trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 239.468 0.292 239.512 ;
    END
  END fz_cp2trim[3]
  PIN fz_cp2trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 238.838 0.292 238.882 ;
    END
  END fz_cp2trim[4]
  PIN fz_cp1trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 242.438 0.292 242.482 ;
    END
  END fz_cp1trim[0]
  PIN fz_cp1trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 241.358 0.292 241.402 ;
    END
  END fz_cp1trim[1]
  PIN fz_cp1trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 241.808 0.292 241.852 ;
    END
  END fz_cp1trim[2]
  PIN fz_cp1trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 240.728 0.292 240.772 ;
    END
  END fz_cp1trim[3]
  PIN fz_cp1trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 241.178 0.292 241.222 ;
    END
  END fz_cp1trim[4]
  PIN fz_cp2trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 239.918 0.292 239.962 ;
    END
  END fz_cp2trim[2]
  PIN clkpll
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 190.328 0.292 190.372 ;
    END
  END clkpll
  PIN clkpll0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 189.878 0.292 189.922 ;
    END
  END clkpll0
  PIN clkpll1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 188.618 0.292 188.662 ;
    END
  END clkpll1
  PIN lock
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 210.488 0.292 210.532 ;
    END
  END lock
  PIN view_dig_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 209.678 0.292 209.722 ;
    END
  END view_dig_out[0]
  PIN view_dig_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 209.858 0.292 209.902 ;
    END
  END view_dig_out[1]
  PIN clkpostdist
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 191.138 0.292 191.182 ;
    END
  END clkpostdist
  PIN idvdisable_bo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 214.808 0.292 214.852 ;
    END
  END idvdisable_bo
  PIN idvfreqao
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 214.178 0.292 214.222 ;
    END
  END idvfreqao
  PIN idvfreqbo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 213.638 0.292 213.682 ;
    END
  END idvfreqbo
  PIN idvpulseo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 213.008 0.292 213.052 ;
    END
  END idvpulseo
  PIN idvtclko
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 213.458 0.292 213.502 ;
    END
  END idvtclko
  PIN idvtctrlo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 212.828 0.292 212.872 ;
    END
  END idvtctrlo
  PIN idvtdo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 212.378 0.292 212.422 ;
    END
  END idvtdo
  PIN idvtreso
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 211.658 0.292 211.702 ;
    END
  END idvtreso
  PIN tdo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 212.198 0.292 212.242 ;
    END
  END tdo
  PIN viewanabus[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 207.518 0.292 207.562 ;
    END
  END viewanabus[0]
  PIN viewanabus[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 207.788 0.292 207.832 ;
    END
  END viewanabus[1]
  PIN ssc_frac_step[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 257.108 0.292 257.152 ;
    END
  END ssc_frac_step[0]
  PIN ssc_frac_step[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 256.478 0.292 256.522 ;
    END
  END ssc_frac_step[1]
  PIN ssc_frac_step[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 256.928 0.292 256.972 ;
    END
  END ssc_frac_step[2]
  PIN ssc_frac_step[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 256.298 0.292 256.342 ;
    END
  END ssc_frac_step[3]
  PIN ssc_frac_step[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 255.848 0.292 255.892 ;
    END
  END ssc_frac_step[4]
  PIN ssc_frac_step[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 255.668 0.292 255.712 ;
    END
  END ssc_frac_step[6]
  PIN ssc_frac_step[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 255.038 0.292 255.082 ;
    END
  END ssc_frac_step[7]
  PIN ssc_frac_step[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 255.218 0.292 255.262 ;
    END
  END ssc_frac_step[5]
  PIN ssc_frac_step[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 253.958 0.292 254.002 ;
    END
  END ssc_frac_step[9]
  PIN ssc_frac_step[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 254.408 0.292 254.452 ;
    END
  END ssc_frac_step[10]
  PIN ssc_frac_step[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 253.778 0.292 253.822 ;
    END
  END ssc_frac_step[11]
  PIN ssc_frac_step[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 253.328 0.292 253.372 ;
    END
  END ssc_frac_step[12]
  PIN ssc_frac_step[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 252.698 0.292 252.742 ;
    END
  END ssc_frac_step[13]
  PIN ssc_frac_step[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 253.148 0.292 253.192 ;
    END
  END ssc_frac_step[14]
  PIN ssc_frac_step[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 252.518 0.292 252.562 ;
    END
  END ssc_frac_step[15]
  PIN ssc_frac_step[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 252.068 0.292 252.112 ;
    END
  END ssc_frac_step[16]
  PIN ssc_frac_step[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 251.438 0.292 251.482 ;
    END
  END ssc_frac_step[17]
  PIN ssc_frac_step[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 251.888 0.292 251.932 ;
    END
  END ssc_frac_step[18]
  PIN ssc_frac_step[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 254.588 0.292 254.632 ;
    END
  END ssc_frac_step[8]
  PIN ssc_frac_step[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 251.258 0.292 251.302 ;
    END
  END ssc_frac_step[19]
  PIN ssc_frac_step[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 250.178 0.292 250.222 ;
    END
  END ssc_frac_step[21]
  PIN ssc_frac_step[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 250.628 0.292 250.672 ;
    END
  END ssc_frac_step[22]
  PIN ssc_frac_step[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 249.998 0.292 250.042 ;
    END
  END ssc_frac_step[23]
  PIN ssc_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 257.558 0.292 257.602 ;
    END
  END ssc_en
  PIN ssc_cyc_to_peak_m1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 260.258 0.292 260.302 ;
    END
  END ssc_cyc_to_peak_m1[0]
  PIN ssc_cyc_to_peak_m1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 259.628 0.292 259.672 ;
    END
  END ssc_cyc_to_peak_m1[1]
  PIN ssc_cyc_to_peak_m1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 260.078 0.292 260.122 ;
    END
  END ssc_cyc_to_peak_m1[2]
  PIN ssc_cyc_to_peak_m1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 259.448 0.292 259.492 ;
    END
  END ssc_cyc_to_peak_m1[3]
  PIN ssc_cyc_to_peak_m1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 258.998 0.292 259.042 ;
    END
  END ssc_cyc_to_peak_m1[4]
  PIN ssc_frac_step[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 250.808 0.292 250.852 ;
    END
  END ssc_frac_step[20]
  PIN ssc_cyc_to_peak_m1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 258.818 0.292 258.862 ;
    END
  END ssc_cyc_to_peak_m1[5]
  PIN ssc_cyc_to_peak_m1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 258.188 0.292 258.232 ;
    END
  END ssc_cyc_to_peak_m1[7]
  PIN ssc_cyc_to_peak_m1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 257.738 0.292 257.782 ;
    END
  END ssc_cyc_to_peak_m1[8]
  PIN mash_order_plus_one
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 260.708 0.292 260.752 ;
    END
  END mash_order_plus_one
  PIN mdiv_ratio[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 262.598 0.292 262.642 ;
    END
  END mdiv_ratio[0]
  PIN ssc_cyc_to_peak_m1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 258.368 0.292 258.412 ;
    END
  END ssc_cyc_to_peak_m1[6]
  PIN mdiv_ratio[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 261.968 0.292 262.012 ;
    END
  END mdiv_ratio[2]
  PIN mdiv_ratio[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 261.518 0.292 261.562 ;
    END
  END mdiv_ratio[3]
  PIN mdiv_ratio[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 261.338 0.292 261.382 ;
    END
  END mdiv_ratio[4]
  PIN mdiv_ratio[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 260.888 0.292 260.932 ;
    END
  END mdiv_ratio[5]
  PIN mdiv_ratio[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 262.148 0.292 262.192 ;
    END
  END mdiv_ratio[1]
  PIN fraction[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 270.158 0.292 270.202 ;
    END
  END fraction[1]
  PIN fraction[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 269.078 0.292 269.122 ;
    END
  END fraction[2]
  PIN fraction[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 269.708 0.292 269.752 ;
    END
  END fraction[0]
  PIN fraction[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 268.448 0.292 268.492 ;
    END
  END fraction[4]
  PIN fraction[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 268.898 0.292 268.942 ;
    END
  END fraction[5]
  PIN fraction[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 269.528 0.292 269.572 ;
    END
  END fraction[3]
  PIN fraction[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 268.268 0.292 268.312 ;
    END
  END fraction[7]
  PIN fraction[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 267.188 0.292 267.232 ;
    END
  END fraction[8]
  PIN fraction[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 267.638 0.292 267.682 ;
    END
  END fraction[9]
  PIN fraction[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 266.558 0.292 266.602 ;
    END
  END fraction[10]
  PIN fraction[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 267.008 0.292 267.052 ;
    END
  END fraction[11]
  PIN fraction[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 265.928 0.292 265.972 ;
    END
  END fraction[12]
  PIN fraction[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 267.818 0.292 267.862 ;
    END
  END fraction[6]
  PIN fraction[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 265.298 0.292 265.342 ;
    END
  END fraction[14]
  PIN fraction[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 265.748 0.292 265.792 ;
    END
  END fraction[15]
  PIN fraction[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 264.668 0.292 264.712 ;
    END
  END fraction[16]
  PIN fraction[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 265.118 0.292 265.162 ;
    END
  END fraction[17]
  PIN fraction[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 264.038 0.292 264.082 ;
    END
  END fraction[18]
  PIN fraction[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 266.378 0.292 266.422 ;
    END
  END fraction[13]
  PIN fraction[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 263.408 0.292 263.452 ;
    END
  END fraction[20]
  PIN fraction[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 263.858 0.292 263.902 ;
    END
  END fraction[21]
  PIN fraction[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 262.778 0.292 262.822 ;
    END
  END fraction[22]
  PIN fraction[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 264.488 0.292 264.532 ;
    END
  END fraction[19]
  PIN fraction[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 263.228 0.292 263.272 ;
    END
  END fraction[23]
  PIN ratio[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 270.788 0.292 270.832 ;
    END
  END ratio[1]
  PIN ratio[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 270.968 0.292 271.012 ;
    END
  END ratio[2]
  PIN ratio[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 271.418 0.292 271.462 ;
    END
  END ratio[3]
  PIN ratio[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 271.598 0.292 271.642 ;
    END
  END ratio[4]
  PIN ratio[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 270.338 0.292 270.382 ;
    END
  END ratio[0]
  PIN ratio[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 272.048 0.292 272.092 ;
    END
  END ratio[5]
  PIN ratio[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 272.228 0.292 272.272 ;
    END
  END ratio[6]
  PIN ratio[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 272.858 0.292 272.902 ;
    END
  END ratio[8]
  PIN ratio[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 273.308 0.292 273.352 ;
    END
  END ratio[9]
  PIN ratio[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 272.678 0.292 272.722 ;
    END
  END ratio[7]
  PIN pllfwen_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 273.938 0.292 273.982 ;
    END
  END pllfwen_b
  PIN fz_vcotrim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 223.538 0.292 223.582 ;
    END
  END fz_vcotrim[0]
  PIN bypass
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 274.118 0.292 274.162 ;
    END
  END bypass
  PIN clkref
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 201.218 0.292 201.262 ;
    END
  END clkref
  PIN pllen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 273.488 0.292 273.532 ;
    END
  END pllen
  PIN tshiftdr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 215.528 0.292 215.572 ;
    END
  END tshiftdr
  PIN trst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 216.158 0.292 216.202 ;
    END
  END trst_n
  PIN treg_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 215.978 0.292 216.022 ;
    END
  END treg_en
  PIN tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 216.608 0.292 216.652 ;
    END
  END tdi
  PIN tupdatedr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 215.348 0.292 215.392 ;
    END
  END tupdatedr
  PIN idvtresi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 217.418 0.292 217.462 ;
    END
  END idvtresi
  PIN idvtdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 218.048 0.292 218.092 ;
    END
  END idvtdi
  PIN idvtctrli
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 218.498 0.292 218.542 ;
    END
  END idvtctrli
  PIN idvtclki
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 219.128 0.292 219.172 ;
    END
  END idvtclki
  PIN idvpulsei
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 218.678 0.292 218.722 ;
    END
  END idvpulsei
  PIN tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 217.868 0.292 217.912 ;
    END
  END tck
  PIN idvfreqbi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 219.308 0.292 219.352 ;
    END
  END idvfreqbi
  PIN idvfreqai
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 219.758 0.292 219.802 ;
    END
  END idvfreqai
  PIN idvdisable_bi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 220.388 0.292 220.432 ;
    END
  END idvdisable_bi
  PIN fz_vcotrim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 222.458 0.292 222.502 ;
    END
  END fz_vcotrim[2]
  PIN ldo_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 279.248 0.292 279.292 ;
    END
  END ldo_enable
  PIN fz_ldo_reftrim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 275.198 0.292 275.242 ;
    END
  END fz_ldo_reftrim[0]
  PIN fz_ldo_reftrim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 274.748 0.292 274.792 ;
    END
  END fz_ldo_reftrim[1]
  PIN fz_ldo_reftrim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 275.378 0.292 275.422 ;
    END
  END fz_ldo_reftrim[2]
  PIN fz_ldo_reftrim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 275.828 0.292 275.872 ;
    END
  END fz_ldo_reftrim[3]
  PIN fz_ldo_fbtrim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 276.458 0.292 276.502 ;
    END
  END fz_ldo_fbtrim[0]
  PIN fz_ldo_fbtrim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 276.008 0.292 276.052 ;
    END
  END fz_ldo_fbtrim[1]
  PIN fz_ldo_fbtrim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 276.638 0.292 276.682 ;
    END
  END fz_ldo_fbtrim[2]
  PIN fz_ldo_fbtrim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 277.088 0.292 277.132 ;
    END
  END fz_ldo_fbtrim[3]
  PIN ldo_vref
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 197.888 0.292 197.932 ;
    END
  END ldo_vref
  PIN fz_ldo_faststart
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 277.268 0.292 277.312 ;
    END
  END fz_ldo_faststart
  PIN fz_ldo_extrefsel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 277.718 0.292 277.762 ;
    END
  END fz_ldo_extrefsel
  PIN fz_ldo_bypass
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 277.898 0.292 277.942 ;
    END
  END fz_ldo_bypass
  PIN fz_ldo_vinvoltsel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 278.348 0.292 278.392 ;
    END
  END fz_ldo_vinvoltsel[0]
  PIN fz_ldo_vinvoltsel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 278.528 0.292 278.572 ;
    END
  END fz_ldo_vinvoltsel[1]
  PIN zdiv1_ratio_p5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 241.988 0.292 242.032 ;
    END
  END zdiv1_ratio_p5
  PIN zdiv1_ratio[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 245.588 0.292 245.632 ;
    END
  END zdiv1_ratio[0]
  PIN zdiv1_ratio[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 245.138 0.292 245.182 ;
    END
  END zdiv1_ratio[1]
  PIN zdiv1_ratio[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 244.508 0.292 244.552 ;
    END
  END zdiv1_ratio[2]
  PIN zdiv1_ratio[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 244.958 0.292 245.002 ;
    END
  END zdiv1_ratio[3]
  PIN zdiv1_ratio[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 243.878 0.292 243.922 ;
    END
  END zdiv1_ratio[4]
  PIN zdiv1_ratio[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 244.328 0.292 244.372 ;
    END
  END zdiv1_ratio[5]
  PIN zdiv1_ratio[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 243.248 0.292 243.292 ;
    END
  END zdiv1_ratio[6]
  PIN zdiv1_ratio[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 243.698 0.292 243.742 ;
    END
  END zdiv1_ratio[7]
  PIN zdiv1_ratio[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 242.618 0.292 242.662 ;
    END
  END zdiv1_ratio[8]
  PIN zdiv1_ratio[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 243.068 0.292 243.112 ;
    END
  END zdiv1_ratio[9]
  PIN zdiv0_ratio_p5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 245.768 0.292 245.812 ;
    END
  END zdiv0_ratio_p5
  PIN zdiv0_ratio[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 249.368 0.292 249.412 ;
    END
  END zdiv0_ratio[0]
  PIN zdiv0_ratio[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 248.738 0.292 248.782 ;
    END
  END zdiv0_ratio[1]
  PIN zdiv0_ratio[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 248.288 0.292 248.332 ;
    END
  END zdiv0_ratio[2]
  PIN zdiv0_ratio[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 247.658 0.292 247.702 ;
    END
  END zdiv0_ratio[3]
  PIN zdiv0_ratio[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 248.108 0.292 248.152 ;
    END
  END zdiv0_ratio[4]
  PIN zdiv0_ratio[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 247.028 0.292 247.072 ;
    END
  END zdiv0_ratio[6]
  PIN zdiv0_ratio[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 246.398 0.292 246.442 ;
    END
  END zdiv0_ratio[7]
  PIN zdiv0_ratio[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 247.478 0.292 247.522 ;
    END
  END zdiv0_ratio[5]
  PIN zdiv0_ratio[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 246.848 0.292 246.892 ;
    END
  END zdiv0_ratio[8]
  PIN zdiv0_ratio[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 246.218 0.292 246.262 ;
    END
  END zdiv0_ratio[9]
  PIN vcodiv_ratio[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 249.548 0.292 249.592 ;
    END
  END vcodiv_ratio[0]
  PIN vcodiv_ratio[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 248.918 0.292 248.962 ;
    END
  END vcodiv_ratio[1]
  PIN idfx_fscan_sdi[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 204.998 0.292 205.042 ;
    END
  END idfx_fscan_sdi[2]
  PIN tcapturedr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 216.788 0.292 216.832 ;
    END
  END tcapturedr
  PIN vss
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.35 0.5175 1.53 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 0.63 0.5175 0.81 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 123.75 0.5175 123.93 189.8285 ;
    END
    PORT
      LAYER m7 ;
        RECT 124.47 0.5175 124.65 189.8285 ;
        RECT 125.19 0.5175 125.37 189.8285 ;
        RECT 125.91 0.5175 126.09 189.8285 ;
        RECT 126.63 0.5175 126.81 189.8285 ;
        RECT 127.35 0.5175 127.53 189.8285 ;
        RECT 128.07 0.5175 128.25 189.8285 ;
        RECT 128.79 0.5175 128.97 189.8285 ;
        RECT 129.51 0.5175 129.69 189.8285 ;
        RECT 130.23 0.5175 130.41 189.8285 ;
        RECT 130.95 0.5175 131.13 189.8285 ;
    END
    PORT
      LAYER m7 ;
        RECT 131.67 0.5175 131.85 189.8285 ;
        RECT 132.39 0.5175 132.57 189.8285 ;
        RECT 133.11 0.5175 133.29 189.8285 ;
        RECT 133.83 0.5175 134.01 189.8285 ;
        RECT 134.55 0.5175 134.73 189.8285 ;
        RECT 135.27 0.5175 135.45 189.8285 ;
    END
    PORT
      LAYER m7 ;
        RECT 153.27 0.5175 153.45 350.01 ;
        RECT 156.15 0.5175 156.33 350.01 ;
        RECT 159.03 0.5175 159.21 350.01 ;
        RECT 164.79 0.5175 164.97 350.01 ;
        RECT 167.67 0.5175 167.85 350.01 ;
        RECT 170.55 0.5175 170.73 350.01 ;
        RECT 176.31 0.5175 176.49 350.01 ;
        RECT 179.19 0.5175 179.37 350.01 ;
        RECT 182.07 0.5175 182.25 350.01 ;
        RECT 187.83 0.5175 188.01 350.01 ;
        RECT 190.71 0.5175 190.89 350.01 ;
        RECT 193.59 0.5175 193.77 350.01 ;
        RECT 199.35 0.5175 199.53 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 153.99 0.5175 154.17 350.01 ;
        RECT 156.87 0.5175 157.05 350.01 ;
        RECT 159.75 0.5175 159.93 350.01 ;
        RECT 165.51 0.5175 165.69 350.01 ;
        RECT 168.39 0.5175 168.57 350.01 ;
        RECT 171.27 0.5175 171.45 350.01 ;
        RECT 177.03 0.5175 177.21 350.01 ;
        RECT 179.91 0.5175 180.09 350.01 ;
        RECT 182.79 0.5175 182.97 350.01 ;
        RECT 188.55 0.5175 188.73 350.01 ;
        RECT 191.43 0.5175 191.61 350.01 ;
        RECT 194.31 0.5175 194.49 350.01 ;
        RECT 200.07 0.5175 200.25 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 189.99 0.5175 190.17 350.01 ;
        RECT 192.87 0.5175 193.05 350.01 ;
        RECT 198.63 0.5175 198.81 350.01 ;
        RECT 152.55 0.5175 152.73 350.01 ;
        RECT 155.43 0.5175 155.61 350.01 ;
        RECT 158.31 0.5175 158.49 350.01 ;
        RECT 164.07 0.5175 164.25 350.01 ;
        RECT 166.95 0.5175 167.13 350.01 ;
        RECT 169.83 0.5175 170.01 350.01 ;
        RECT 175.59 0.5175 175.77 350.01 ;
        RECT 178.47 0.5175 178.65 350.01 ;
        RECT 181.35 0.5175 181.53 350.01 ;
        RECT 187.11 0.5175 187.29 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 102.87 0.5175 103.05 350.01 ;
        RECT 103.59 0.5175 103.77 350.01 ;
        RECT 104.31 0.5175 104.49 350.01 ;
        RECT 105.03 0.5175 105.21 350.01 ;
        RECT 105.75 0.5175 105.93 350.01 ;
        RECT 106.47 0.5175 106.65 350.01 ;
        RECT 107.19 0.5175 107.37 350.01 ;
        RECT 107.91 0.5175 108.09 350.01 ;
        RECT 108.63 0.5175 108.81 350.01 ;
        RECT 109.35 0.5175 109.53 350.01 ;
        RECT 110.07 0.5175 110.25 350.01 ;
        RECT 110.79 0.5175 110.97 350.01 ;
        RECT 111.51 0.5175 111.69 350.01 ;
        RECT 112.23 0.5175 112.41 350.01 ;
        RECT 112.95 0.5175 113.13 350.01 ;
        RECT 113.67 0.5175 113.85 350.01 ;
        RECT 114.39 0.5175 114.57 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 143.19 0.5175 143.37 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 142.47 0.5175 142.65 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 141.75 0.5175 141.93 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 141.03 0.5175 141.21 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 143.91 0.5175 144.09 350.01 ;
        RECT 146.79 0.5175 146.97 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 144.63 0.5175 144.81 350.01 ;
        RECT 147.51 0.5175 147.69 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 146.07 0.5175 146.25 350.01 ;
        RECT 148.95 0.5175 149.13 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 145.35 0.5175 145.53 350.01 ;
        RECT 148.23 0.5175 148.41 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 183.51 0.5175 183.69 350.01 ;
        RECT 189.27 0.5175 189.45 350.01 ;
        RECT 192.15 0.5175 192.33 350.01 ;
        RECT 195.03 0.5175 195.21 350.01 ;
        RECT 200.79 0.5175 200.97 350.01 ;
        RECT 154.71 0.5175 154.89 350.01 ;
        RECT 157.59 0.5175 157.77 350.01 ;
        RECT 160.47 0.5175 160.65 350.01 ;
        RECT 166.23 0.5175 166.41 350.01 ;
        RECT 169.11 0.5175 169.29 350.01 ;
        RECT 171.99 0.5175 172.17 350.01 ;
        RECT 177.75 0.5175 177.93 350.01 ;
        RECT 180.63 0.5175 180.81 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 58.95 0.5175 59.13 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 59.67 0.5175 59.85 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 60.39 0.5175 60.57 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 61.11 0.5175 61.29 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 63.27 0.5175 63.45 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 63.99 0.5175 64.17 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 64.71 0.5175 64.89 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 65.43 0.5175 65.61 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 66.15 0.5175 66.33 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 66.87 0.5175 67.05 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 69.03 0.5175 69.21 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 69.75 0.5175 69.93 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 70.47 0.5175 70.65 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 71.19 0.5175 71.37 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 71.91 0.5175 72.09 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 72.63 0.5175 72.81 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 74.79 0.5175 74.97 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 75.51 0.5175 75.69 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 76.23 0.5175 76.41 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 76.95 0.5175 77.13 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 77.67 0.5175 77.85 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 78.39 0.5175 78.57 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 80.55 0.5175 80.73 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 81.27 0.5175 81.45 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 81.99 0.5175 82.17 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 82.71 0.5175 82.89 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 60.39 0.5175 60.57 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 61.11 0.5175 61.29 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 84.15 0.5175 84.33 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 83.43 0.5175 83.61 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 91.35 0.5175 91.53 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 94.23 0.5175 94.41 350.01 ;
        RECT 94.95 0.5175 95.13 350.01 ;
        RECT 95.67 0.5175 95.85 350.01 ;
        RECT 96.39 0.5175 96.57 350.01 ;
        RECT 97.11 0.5175 97.29 350.01 ;
        RECT 97.83 0.5175 98.01 350.01 ;
        RECT 98.55 0.5175 98.73 350.01 ;
        RECT 99.27 0.5175 99.45 350.01 ;
        RECT 99.99 0.5175 100.17 350.01 ;
        RECT 100.71 0.5175 100.89 350.01 ;
        RECT 101.43 0.5175 101.61 350.01 ;
        RECT 102.15 0.5175 102.33 350.01 ;
        RECT 92.07 0.5175 92.25 350.01 ;
        RECT 92.79 0.5175 92.97 350.01 ;
        RECT 93.51 0.5175 93.69 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 24.39 0.5175 24.57 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 23.67 0.5175 23.85 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 22.95 0.5175 23.13 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 20.79 0.5175 20.97 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 20.07 0.5175 20.25 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 19.35 0.5175 19.53 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 18.63 0.5175 18.81 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.91 0.5175 18.09 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.19 0.5175 17.37 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 38.07 0.5175 38.25 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 37.35 0.5175 37.53 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 36.63 0.5175 36.81 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 35.91 0.5175 36.09 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 35.19 0.5175 35.37 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 34.47 0.5175 34.65 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 32.31 0.5175 32.49 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 31.59 0.5175 31.77 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 40.23 0.5175 40.41 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 40.95 0.5175 41.13 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 41.67 0.5175 41.85 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 42.39 0.5175 42.57 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 43.11 0.5175 43.29 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 43.83 0.5175 44.01 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 45.99 0.5175 46.17 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 46.71 0.5175 46.89 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 47.43 0.5175 47.61 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 48.15 0.5175 48.33 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 48.87 0.5175 49.05 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 49.59 0.5175 49.77 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 51.75 0.5175 51.93 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 52.47 0.5175 52.65 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 53.19 0.5175 53.37 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 53.91 0.5175 54.09 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 54.63 0.5175 54.81 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 55.35 0.5175 55.53 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 57.51 0.5175 57.69 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 58.23 0.5175 58.41 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 4.95 0.5175 5.13 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 2.79 0.5175 2.97 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 2.07 0.5175 2.25 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 9.99 0.5175 10.17 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 7.11 0.5175 7.29 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 6.39 0.5175 6.57 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 5.67 0.5175 5.85 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 9.27 0.5175 9.45 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 10.71 0.5175 10.89 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 13.59 0.5175 13.77 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 14.31 0.5175 14.49 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 15.03 0.5175 15.21 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 12.87 0.5175 13.05 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 11.43 0.5175 11.61 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 30.87 0.5175 31.05 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 30.15 0.5175 30.33 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 29.43 0.5175 29.61 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 28.71 0.5175 28.89 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 26.55 0.5175 26.73 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 25.83 0.5175 26.01 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 25.11 0.5175 25.29 350.01 ;
    END
  END vss
  PIN idfx_fscan_sdi[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 205.178 0.292 205.222 ;
    END
  END idfx_fscan_sdi[1]
  PIN vccdist_nom
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 5.31 164.12 5.49 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 4.59 164.12 4.77 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 3.15 164.12 3.33 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 1.71 164.12 1.89 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 0.99 164.12 1.17 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 2.43 164.12 2.61 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 10.35 164.12 10.53 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 9.63 164.12 9.81 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 6.75 164.12 6.93 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 6.03 164.12 6.21 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 8.91 164.12 9.09 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 7.47 164.12 7.65 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 13.95 164.12 14.13 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 13.23 164.12 13.41 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 15.39 164.12 15.57 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 14.67 164.12 14.85 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 11.07 164.12 11.25 350.01 ;
    END
  END vccdist_nom
  PIN idfx_fscan_sdi[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 205.538 0.292 205.582 ;
    END
  END idfx_fscan_sdi[0]
  PIN odfx_fscan_sdo[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 202.658 0.292 202.702 ;
    END
  END odfx_fscan_sdo[1]
  PIN odfx_fscan_sdo[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 203.018 0.292 203.062 ;
    END
  END odfx_fscan_sdo[0]
  PIN vccldo_hv
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 144.27 272.66 144.45 350.01 ;
        RECT 147.15 272.66 147.33 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 144.99 272.66 145.17 350.01 ;
        RECT 147.87 272.66 148.05 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 152.91 272.66 153.09 350.01 ;
        RECT 155.79 272.66 155.97 350.01 ;
        RECT 158.67 272.66 158.85 350.01 ;
        RECT 164.43 272.66 164.61 350.01 ;
        RECT 167.31 272.66 167.49 350.01 ;
        RECT 170.19 272.66 170.37 350.01 ;
        RECT 175.95 272.66 176.13 350.01 ;
        RECT 178.83 272.66 179.01 350.01 ;
        RECT 181.71 272.66 181.89 350.01 ;
        RECT 187.47 272.66 187.65 350.01 ;
        RECT 190.35 272.66 190.53 350.01 ;
        RECT 193.23 272.66 193.41 350.01 ;
        RECT 198.99 272.66 199.17 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 153.63 272.66 153.81 350.01 ;
        RECT 156.51 272.66 156.69 350.01 ;
        RECT 159.39 272.66 159.57 350.01 ;
        RECT 165.15 272.66 165.33 350.01 ;
        RECT 168.03 272.66 168.21 350.01 ;
        RECT 170.91 272.66 171.09 350.01 ;
        RECT 176.67 272.66 176.85 350.01 ;
        RECT 179.55 272.66 179.73 350.01 ;
        RECT 182.43 272.66 182.61 350.01 ;
        RECT 188.19 272.66 188.37 350.01 ;
        RECT 191.07 272.66 191.25 350.01 ;
        RECT 193.95 272.66 194.13 350.01 ;
        RECT 199.71 272.66 199.89 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 171.63 272.66 171.81 350.01 ;
        RECT 177.39 272.66 177.57 350.01 ;
        RECT 180.27 272.66 180.45 350.01 ;
        RECT 183.15 272.66 183.33 350.01 ;
        RECT 188.91 272.66 189.09 350.01 ;
        RECT 191.79 272.66 191.97 350.01 ;
        RECT 194.67 272.66 194.85 350.01 ;
        RECT 200.43 272.66 200.61 350.01 ;
        RECT 154.35 272.66 154.53 350.01 ;
        RECT 157.23 272.66 157.41 350.01 ;
        RECT 160.11 272.66 160.29 350.01 ;
        RECT 165.87 272.66 166.05 350.01 ;
        RECT 168.75 272.66 168.93 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 141.39 272.66 141.57 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 142.11 272.66 142.29 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 142.83 272.66 143.01 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 145.71 272.66 145.89 350.01 ;
        RECT 148.59 272.66 148.77 350.01 ;
    END
  END vccldo_hv
  PIN odfx_fscan_sdo[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 202.478 0.292 202.522 ;
    END
  END odfx_fscan_sdo[2]
  PIN idfx_fscan_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 200.498 0.292 200.542 ;
    END
  END idfx_fscan_mode
  PIN idfx_fscan_shiften
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 200.138 0.292 200.182 ;
    END
  END idfx_fscan_shiften
  PIN idfx_fscan_rstbypen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 199.958 0.292 200.002 ;
    END
  END idfx_fscan_rstbypen
  PIN idfx_fscan_byprstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 197.618 0.292 197.662 ;
    END
  END idfx_fscan_byprstb
  PIN idfx_fscan_clkungate
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 197.438 0.292 197.482 ;
    END
  END idfx_fscan_clkungate
  PIN vnnaon_nom
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 84.87 184.16 85.05 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 85.59 184.16 85.77 350.01 ;
        RECT 86.31 184.16 86.49 350.01 ;
        RECT 87.03 184.16 87.21 350.01 ;
        RECT 87.75 184.16 87.93 350.01 ;
    END
  END vnnaon_nom
  PIN vccdig_nom
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 46.35 156.02 46.53 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 47.79 156.02 47.97 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 49.23 156.02 49.41 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 52.11 156.02 52.29 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 53.55 156.02 53.73 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 54.99 156.02 55.17 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 57.87 156.02 58.05 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 59.31 156.02 59.49 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 60.75 156.02 60.93 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 63.63 156.02 63.81 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 65.07 156.02 65.25 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 66.51 156.02 66.69 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 69.39 156.02 69.57 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 70.83 156.02 71.01 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 72.27 156.02 72.45 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 75.15 156.02 75.33 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 76.59 156.02 76.77 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 78.03 156.02 78.21 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 80.91 156.02 81.09 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 82.35 156.02 82.53 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 60.75 156.02 60.93 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 83.79 156.02 83.97 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 123.75 190.18 123.93 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 125.19 190.18 125.37 350.01 ;
        RECT 125.91 190.18 126.09 350.01 ;
        RECT 126.63 190.18 126.81 350.01 ;
        RECT 127.35 190.18 127.53 350.01 ;
        RECT 128.07 190.18 128.25 350.01 ;
        RECT 128.79 190.18 128.97 350.01 ;
        RECT 129.51 190.18 129.69 350.01 ;
        RECT 130.23 190.18 130.41 350.01 ;
        RECT 130.95 190.18 131.13 350.01 ;
        RECT 131.67 190.18 131.85 350.01 ;
        RECT 132.39 190.18 132.57 350.01 ;
        RECT 133.11 190.18 133.29 350.01 ;
        RECT 133.83 190.18 134.01 350.01 ;
        RECT 134.55 190.18 134.73 350.01 ;
        RECT 135.27 190.18 135.45 350.01 ;
        RECT 124.47 190.18 124.65 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 24.75 156.02 24.93 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 26.19 156.02 26.37 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 29.07 156.02 29.25 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 30.51 156.02 30.69 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 31.95 156.02 32.13 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 34.83 156.02 35.01 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 36.27 156.02 36.45 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 37.71 156.02 37.89 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 23.31 156.02 23.49 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 20.43 156.02 20.61 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 18.99 156.02 19.17 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.55 156.02 17.73 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 40.59 156.02 40.77 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 42.03 156.02 42.21 350.01 ;
    END
    PORT
      LAYER m7 ;
        RECT 43.47 156.02 43.65 350.01 ;
    END
  END vccdig_nom
  PIN powergood_vnn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 187.358 0.292 187.402 ;
    END
  END powergood_vnn
  OBS
    LAYER v6 ;
      RECT 0.62 118.26 0.82 118.38 ;
      RECT 1.34 118.26 1.54 118.38 ;
      RECT 7.1 118.26 7.3 118.38 ;
      RECT 5.66 118.26 5.86 118.38 ;
      RECT 2.78 118.26 2.98 118.38 ;
      RECT 0.62 121.498 0.82 121.618 ;
      RECT 1.34 121.498 1.54 121.618 ;
      RECT 2.06 121.498 2.26 121.618 ;
      RECT 2.78 121.498 2.98 121.618 ;
      RECT 4.94 121.498 5.14 121.618 ;
      RECT 5.66 121.498 5.86 121.618 ;
      RECT 6.38 121.498 6.58 121.618 ;
      RECT 7.1 121.498 7.3 121.618 ;
      RECT 6.38 121.02 6.58 121.14 ;
      RECT 7.1 121.02 7.3 121.14 ;
      RECT 1.34 121.02 1.54 121.14 ;
      RECT 4.94 121.02 5.14 121.14 ;
      RECT 0.62 120.78 0.82 120.9 ;
      RECT 2.78 120.78 2.98 120.9 ;
      RECT 5.66 120.78 5.86 120.9 ;
      RECT 0.62 124.018 0.82 124.138 ;
      RECT 1.34 124.018 1.54 124.138 ;
      RECT 2.06 124.018 2.26 124.138 ;
      RECT 2.78 124.018 2.98 124.138 ;
      RECT 4.94 124.018 5.14 124.138 ;
      RECT 5.66 124.018 5.86 124.138 ;
      RECT 6.38 124.018 6.58 124.138 ;
      RECT 7.1 124.018 7.3 124.138 ;
      RECT 1.34 123.54 1.54 123.66 ;
      RECT 4.94 123.54 5.14 123.66 ;
    LAYER m7 EXCEPTPGNET ;
      RECT 0 0 201.96 413.28 ;
    LAYER m6 SPACING 0 ;
      RECT 0 0 201.96 413.28 ;
    LAYER m5 ;
      RECT 0 0 201.96 413.28 ;
    LAYER m4 ;
      RECT 0 0 201.96 413.28 ;
    LAYER m3 ;
      RECT 0 0 201.96 413.28 ;
    LAYER m2 ;
      RECT 0 0 201.96 413.28 ;
    LAYER m1 ;
      RECT 0 0 201.96 413.28 ;
    LAYER v6 ;
      RECT 4.94 118.5 5.14 118.62 ;
      RECT 6.38 118.5 6.58 118.62 ;
      RECT 7.1 118.978 7.3 119.098 ;
      RECT 6.38 118.978 6.58 119.098 ;
      RECT 5.66 118.978 5.86 119.098 ;
      RECT 4.94 118.978 5.14 119.098 ;
      RECT 2.78 118.978 2.98 119.098 ;
      RECT 2.06 118.978 2.26 119.098 ;
      RECT 1.34 118.978 1.54 119.098 ;
      RECT 0.62 118.978 0.82 119.098 ;
      RECT 35.9 196.38 36.1 196.5 ;
      RECT 34.82 195.902 35.02 196.022 ;
      RECT 36.26 195.902 36.46 196.022 ;
      RECT 35.54 195.36 35.74 195.48 ;
      RECT 35.54 197.88 35.74 198 ;
      RECT 36.62 196.62 36.82 196.74 ;
      RECT 35.18 196.62 35.38 196.74 ;
      RECT 34.46 199.14 34.66 199.26 ;
      RECT 35.9 199.14 36.1 199.26 ;
      RECT 36.62 198.9 36.82 199.02 ;
      RECT 35.18 198.9 35.38 199.02 ;
      RECT 34.82 198.422 35.02 198.542 ;
      RECT 36.26 198.182 36.46 198.302 ;
      RECT 35.54 200.4 35.74 200.52 ;
      RECT 36.62 201.66 36.82 201.78 ;
      RECT 35.18 201.66 35.38 201.78 ;
      RECT 34.46 201.66 34.66 201.78 ;
      RECT 35.9 201.42 36.1 201.54 ;
      RECT 36.26 200.942 36.46 201.062 ;
      RECT 34.82 200.702 35.02 200.822 ;
      RECT 34.82 203.222 35.02 203.342 ;
      RECT 35.54 202.68 35.74 202.8 ;
      RECT 35.18 204.18 35.38 204.3 ;
      RECT 35.9 204.18 36.1 204.3 ;
      RECT 36.62 204.18 36.82 204.3 ;
      RECT 34.46 203.94 34.66 204.06 ;
      RECT 36.26 203.462 36.46 203.582 ;
      RECT 36.26 205.982 36.46 206.102 ;
      RECT 34.82 205.742 35.02 205.862 ;
      RECT 35.54 205.44 35.74 205.56 ;
      RECT 36.62 206.7 36.82 206.82 ;
      RECT 35.9 206.7 36.1 206.82 ;
      RECT 34.46 206.7 34.66 206.82 ;
      RECT 35.18 206.46 35.38 206.58 ;
      RECT 36.26 208.502 36.46 208.622 ;
      RECT 34.82 208.262 35.02 208.382 ;
      RECT 35.54 207.96 35.74 208.08 ;
      RECT 36.26 210.09 36.46 210.21 ;
      RECT 34.82 210.09 35.02 210.21 ;
      RECT 36.62 209.46 36.82 209.58 ;
      RECT 35.9 209.46 36.1 209.58 ;
      RECT 35.18 209.46 35.38 209.58 ;
      RECT 34.46 209.46 34.66 209.58 ;
      RECT 34.82 211.35 35.02 211.47 ;
      RECT 36.26 211.35 36.46 211.47 ;
      RECT 34.46 210.72 34.66 210.84 ;
      RECT 35.18 210.72 35.38 210.84 ;
      RECT 35.9 210.72 36.1 210.84 ;
      RECT 36.62 210.72 36.82 210.84 ;
      RECT 34.82 212.61 35.02 212.73 ;
      RECT 36.26 212.61 36.46 212.73 ;
      RECT 36.62 211.98 36.82 212.1 ;
      RECT 35.9 211.98 36.1 212.1 ;
      RECT 35.18 211.98 35.38 212.1 ;
      RECT 34.46 211.98 34.66 212.1 ;
      RECT 34.82 213.87 35.02 213.99 ;
      RECT 36.26 213.87 36.46 213.99 ;
      RECT 34.46 213.24 34.66 213.36 ;
      RECT 35.18 213.24 35.38 213.36 ;
      RECT 35.9 213.24 36.1 213.36 ;
      RECT 36.62 213.24 36.82 213.36 ;
      RECT 7.1 143.46 7.3 143.58 ;
      RECT 0.62 143.46 0.82 143.58 ;
      RECT 2.78 140.94 2.98 141.06 ;
      RECT 5.66 140.94 5.86 141.06 ;
      RECT 7.1 140.94 7.3 141.06 ;
      RECT 0.62 140.94 0.82 141.06 ;
      RECT 4.94 141.18 5.14 141.3 ;
      RECT 6.38 141.18 6.58 141.3 ;
      RECT 1.34 141.18 1.54 141.3 ;
      RECT 7.1 136.618 7.3 136.738 ;
      RECT 6.38 136.618 6.58 136.738 ;
      RECT 5.66 136.618 5.86 136.738 ;
      RECT 4.94 136.618 5.14 136.738 ;
      RECT 2.78 136.618 2.98 136.738 ;
      RECT 2.06 136.618 2.26 136.738 ;
      RECT 1.34 136.618 1.54 136.738 ;
      RECT 0.62 136.618 0.82 136.738 ;
      RECT 4.94 138.42 5.14 138.54 ;
      RECT 6.38 138.42 6.58 138.54 ;
      RECT 0.62 138.42 0.82 138.54 ;
      RECT 2.78 138.66 2.98 138.78 ;
      RECT 1.34 138.66 1.54 138.78 ;
      RECT 7.1 138.66 7.3 138.78 ;
      RECT 5.66 138.66 5.86 138.78 ;
      RECT 7.1 139.138 7.3 139.258 ;
      RECT 6.38 139.138 6.58 139.258 ;
      RECT 5.66 139.138 5.86 139.258 ;
      RECT 4.94 139.138 5.14 139.258 ;
      RECT 2.78 139.138 2.98 139.258 ;
      RECT 2.06 139.138 2.26 139.258 ;
      RECT 1.34 139.138 1.54 139.258 ;
      RECT 0.62 139.138 0.82 139.258 ;
      RECT 7.1 134.098 7.3 134.218 ;
      RECT 6.38 134.098 6.58 134.218 ;
      RECT 5.66 134.098 5.86 134.218 ;
      RECT 4.94 134.098 5.14 134.218 ;
      RECT 2.78 134.098 2.98 134.218 ;
      RECT 2.06 134.098 2.26 134.218 ;
      RECT 1.34 134.098 1.54 134.218 ;
      RECT 0.62 134.098 0.82 134.218 ;
      RECT 4.94 135.9 5.14 136.02 ;
      RECT 6.38 135.9 6.58 136.02 ;
      RECT 2.78 136.14 2.98 136.26 ;
      RECT 5.66 136.14 5.86 136.26 ;
      RECT 7.1 136.14 7.3 136.26 ;
      RECT 4.94 131.1 5.14 131.22 ;
      RECT 6.38 131.1 6.58 131.22 ;
      RECT 1.34 131.1 1.54 131.22 ;
      RECT 7.1 131.578 7.3 131.698 ;
      RECT 6.38 131.578 6.58 131.698 ;
      RECT 5.66 131.578 5.86 131.698 ;
      RECT 4.94 131.578 5.14 131.698 ;
      RECT 2.78 131.578 2.98 131.698 ;
      RECT 2.06 131.578 2.26 131.698 ;
      RECT 1.34 131.578 1.54 131.698 ;
      RECT 0.62 131.578 0.82 131.698 ;
      RECT 2.78 133.38 2.98 133.5 ;
      RECT 5.66 133.38 5.86 133.5 ;
      RECT 7.1 133.38 7.3 133.5 ;
      RECT 0.62 133.38 0.82 133.5 ;
      RECT 6.38 133.62 6.58 133.74 ;
      RECT 4.94 133.62 5.14 133.74 ;
      RECT 1.34 133.62 1.54 133.74 ;
      RECT 2.78 128.34 2.98 128.46 ;
      RECT 5.66 128.34 5.86 128.46 ;
      RECT 7.1 128.34 7.3 128.46 ;
      RECT 0.62 128.34 0.82 128.46 ;
      RECT 4.94 128.58 5.14 128.7 ;
      RECT 6.38 128.58 6.58 128.7 ;
      RECT 1.34 128.58 1.54 128.7 ;
      RECT 6.38 129.058 6.58 129.178 ;
      RECT 4.94 129.058 5.14 129.178 ;
      RECT 2.06 129.058 2.26 129.178 ;
      RECT 0.62 129.058 0.82 129.178 ;
      RECT 7.1 129.298 7.3 129.418 ;
      RECT 5.66 129.298 5.86 129.418 ;
      RECT 2.78 129.298 2.98 129.418 ;
      RECT 1.34 129.298 1.54 129.418 ;
      RECT 7.1 130.86 7.3 130.98 ;
      RECT 5.66 130.86 5.86 130.98 ;
      RECT 2.78 130.86 2.98 130.98 ;
      RECT 0.62 130.86 0.82 130.98 ;
      RECT 7.1 125.82 7.3 125.94 ;
      RECT 5.66 125.82 5.86 125.94 ;
      RECT 2.78 125.82 2.98 125.94 ;
      RECT 0.62 125.82 0.82 125.94 ;
      RECT 6.38 126.06 6.58 126.18 ;
      RECT 4.94 126.06 5.14 126.18 ;
      RECT 1.34 126.06 1.54 126.18 ;
      RECT 7.1 126.538 7.3 126.658 ;
      RECT 6.38 126.538 6.58 126.658 ;
      RECT 5.66 126.538 5.86 126.658 ;
      RECT 4.94 126.538 5.14 126.658 ;
      RECT 2.78 126.538 2.98 126.658 ;
      RECT 2.06 126.538 2.26 126.658 ;
      RECT 1.34 126.538 1.54 126.658 ;
      RECT 0.62 126.538 0.82 126.658 ;
      RECT 7.1 123.3 7.3 123.42 ;
      RECT 5.66 123.3 5.86 123.42 ;
      RECT 2.78 123.3 2.98 123.42 ;
      RECT 0.62 123.3 0.82 123.42 ;
      RECT 6.38 123.54 6.58 123.66 ;
      RECT 6.02 169.92 6.22 170.04 ;
      RECT 5.3 169.92 5.5 170.04 ;
      RECT 4.58 169.92 4.78 170.04 ;
      RECT 3.14 169.92 3.34 170.04 ;
      RECT 2.42 169.92 2.62 170.04 ;
      RECT 1.7 169.92 1.9 170.04 ;
      RECT 0.98 169.92 1.18 170.04 ;
      RECT 1.34 171.18 1.54 171.3 ;
      RECT 4.94 171.18 5.14 171.3 ;
      RECT 6.38 171.18 6.58 171.3 ;
      RECT 2.78 171.42 2.98 171.54 ;
      RECT 5.66 171.42 5.86 171.54 ;
      RECT 7.1 171.42 7.3 171.54 ;
      RECT 2.06 171.42 2.26 171.54 ;
      RECT 0.62 171.42 0.82 171.54 ;
      RECT 7.46 167.4 7.66 167.52 ;
      RECT 6.74 167.4 6.94 167.52 ;
      RECT 6.02 167.4 6.22 167.52 ;
      RECT 5.3 167.4 5.5 167.52 ;
      RECT 4.58 167.4 4.78 167.52 ;
      RECT 3.14 167.4 3.34 167.52 ;
      RECT 2.42 167.4 2.62 167.52 ;
      RECT 1.7 167.4 1.9 167.52 ;
      RECT 0.98 167.4 1.18 167.52 ;
      RECT 6.38 168.66 6.58 168.78 ;
      RECT 2.78 168.66 2.98 168.78 ;
      RECT 1.34 168.66 1.54 168.78 ;
      RECT 0.62 168.9 0.82 169.02 ;
      RECT 2.06 168.9 2.26 169.02 ;
      RECT 4.94 168.9 5.14 169.02 ;
      RECT 5.66 168.9 5.86 169.02 ;
      RECT 7.1 168.9 7.3 169.02 ;
      RECT 1.34 163.86 1.54 163.98 ;
      RECT 2.06 163.86 2.26 163.98 ;
      RECT 2.78 163.86 2.98 163.98 ;
      RECT 4.94 163.86 5.14 163.98 ;
      RECT 6.38 163.86 6.58 163.98 ;
      RECT 7.46 164.88 7.66 165 ;
      RECT 6.74 164.88 6.94 165 ;
      RECT 6.02 164.88 6.22 165 ;
      RECT 5.3 164.88 5.5 165 ;
      RECT 4.58 164.88 4.78 165 ;
      RECT 3.14 164.88 3.34 165 ;
      RECT 2.42 164.88 2.62 165 ;
      RECT 1.7 164.88 1.9 165 ;
      RECT 0.98 164.88 1.18 165 ;
      RECT 1.34 166.14 1.54 166.26 ;
      RECT 0.62 166.38 0.82 166.5 ;
      RECT 2.06 166.38 2.26 166.5 ;
      RECT 2.78 166.38 2.98 166.5 ;
      RECT 4.94 166.38 5.14 166.5 ;
      RECT 5.66 166.38 5.86 166.5 ;
      RECT 6.38 166.38 6.58 166.5 ;
      RECT 7.1 166.38 7.3 166.5 ;
      RECT 7.1 163.62 7.3 163.74 ;
      RECT 5.66 163.62 5.86 163.74 ;
      RECT 0.62 163.62 0.82 163.74 ;
      RECT 1.34 158.58 1.54 158.7 ;
      RECT 2.78 158.58 2.98 158.7 ;
      RECT 5.66 158.58 5.86 158.7 ;
      RECT 7.1 158.82 7.3 158.94 ;
      RECT 6.38 158.82 6.58 158.94 ;
      RECT 4.94 158.82 5.14 158.94 ;
      RECT 2.06 158.82 2.26 158.94 ;
      RECT 0.62 158.82 0.82 158.94 ;
      RECT 1.34 156.06 1.54 156.18 ;
      RECT 4.94 156.06 5.14 156.18 ;
      RECT 6.38 156.06 6.58 156.18 ;
      RECT 2.78 156.3 2.98 156.42 ;
      RECT 2.06 156.3 2.26 156.42 ;
      RECT 0.62 156.3 0.82 156.42 ;
      RECT 7.1 156.3 7.3 156.42 ;
      RECT 5.66 156.3 5.86 156.42 ;
      RECT 1.34 153.54 1.54 153.66 ;
      RECT 2.78 153.54 2.98 153.66 ;
      RECT 6.38 153.54 6.58 153.66 ;
      RECT 7.1 153.78 7.3 153.9 ;
      RECT 5.66 153.78 5.86 153.9 ;
      RECT 4.94 153.78 5.14 153.9 ;
      RECT 2.06 153.78 2.26 153.9 ;
      RECT 0.62 153.78 0.82 153.9 ;
      RECT 1.34 148.5 1.54 148.62 ;
      RECT 4.94 148.5 5.14 148.62 ;
      RECT 6.38 148.5 6.58 148.62 ;
      RECT 7.1 148.74 7.3 148.86 ;
      RECT 5.66 148.74 5.86 148.86 ;
      RECT 2.78 148.74 2.98 148.86 ;
      RECT 2.06 148.74 2.26 148.86 ;
      RECT 0.62 148.74 0.82 148.86 ;
      RECT 7.1 145.98 7.3 146.1 ;
      RECT 6.38 145.98 6.58 146.1 ;
      RECT 5.66 145.98 5.86 146.1 ;
      RECT 4.94 145.98 5.14 146.1 ;
      RECT 2.78 145.98 2.98 146.1 ;
      RECT 2.06 145.98 2.26 146.1 ;
      RECT 1.34 145.98 1.54 146.1 ;
      RECT 0.62 145.98 0.82 146.1 ;
      RECT 4.94 143.7 5.14 143.82 ;
      RECT 6.38 143.7 6.58 143.82 ;
      RECT 1.34 143.7 1.54 143.82 ;
      RECT 2.78 143.46 2.98 143.58 ;
      RECT 5.66 143.46 5.86 143.58 ;
      RECT 7.46 169.92 7.66 170.04 ;
      RECT 6.74 169.92 6.94 170.04 ;
      RECT 1.34 178.74 1.54 178.86 ;
      RECT 2.78 178.74 2.98 178.86 ;
      RECT 5.66 178.74 5.86 178.86 ;
      RECT 7.1 178.74 7.3 178.86 ;
      RECT 6.38 178.98 6.58 179.1 ;
      RECT 4.94 178.98 5.14 179.1 ;
      RECT 2.06 178.98 2.26 179.1 ;
      RECT 0.62 178.98 0.82 179.1 ;
      RECT 7.46 180 7.66 180.12 ;
      RECT 6.74 180 6.94 180.12 ;
      RECT 6.02 180 6.22 180.12 ;
      RECT 5.3 180 5.5 180.12 ;
      RECT 4.58 180 4.78 180.12 ;
      RECT 3.14 180 3.34 180.12 ;
      RECT 2.42 180 2.62 180.12 ;
      RECT 1.7 180 1.9 180.12 ;
      RECT 0.98 180 1.18 180.12 ;
      RECT 7.46 174.96 7.66 175.08 ;
      RECT 6.74 174.96 6.94 175.08 ;
      RECT 6.02 174.96 6.22 175.08 ;
      RECT 5.3 174.96 5.5 175.08 ;
      RECT 4.58 174.96 4.78 175.08 ;
      RECT 3.14 174.96 3.34 175.08 ;
      RECT 2.42 174.96 2.62 175.08 ;
      RECT 1.7 174.96 1.9 175.08 ;
      RECT 0.98 174.96 1.18 175.08 ;
      RECT 1.34 176.22 1.54 176.34 ;
      RECT 2.78 176.22 2.98 176.34 ;
      RECT 5.66 176.22 5.86 176.34 ;
      RECT 7.1 176.22 7.3 176.34 ;
      RECT 0.62 176.46 0.82 176.58 ;
      RECT 2.06 176.46 2.26 176.58 ;
      RECT 4.94 176.46 5.14 176.58 ;
      RECT 6.38 176.46 6.58 176.58 ;
      RECT 7.46 177.48 7.66 177.6 ;
      RECT 6.74 177.48 6.94 177.6 ;
      RECT 6.02 177.48 6.22 177.6 ;
      RECT 5.3 177.48 5.5 177.6 ;
      RECT 4.58 177.48 4.78 177.6 ;
      RECT 3.14 177.48 3.34 177.6 ;
      RECT 2.42 177.48 2.62 177.6 ;
      RECT 1.7 177.48 1.9 177.6 ;
      RECT 0.98 177.48 1.18 177.6 ;
      RECT 7.46 172.44 7.66 172.56 ;
      RECT 6.74 172.44 6.94 172.56 ;
      RECT 6.02 172.44 6.22 172.56 ;
      RECT 5.3 172.44 5.5 172.56 ;
      RECT 4.58 172.44 4.78 172.56 ;
      RECT 3.14 172.44 3.34 172.56 ;
      RECT 2.42 172.44 2.62 172.56 ;
      RECT 1.7 172.44 1.9 172.56 ;
      RECT 0.98 172.44 1.18 172.56 ;
      RECT 1.34 173.7 1.54 173.82 ;
      RECT 2.78 173.7 2.98 173.82 ;
      RECT 5.66 173.7 5.86 173.82 ;
      RECT 0.62 173.94 0.82 174.06 ;
      RECT 4.94 173.94 5.14 174.06 ;
      RECT 2.06 173.94 2.26 174.06 ;
      RECT 6.38 173.94 6.58 174.06 ;
      RECT 7.1 173.94 7.3 174.06 ;
      RECT 6.38 196.62 6.58 196.74 ;
      RECT 7.46 196.922 7.66 197.042 ;
      RECT 6.74 196.922 6.94 197.042 ;
      RECT 6.02 196.922 6.22 197.042 ;
      RECT 5.3 196.922 5.5 197.042 ;
      RECT 4.58 196.922 4.78 197.042 ;
      RECT 6.38 198.9 6.58 199.02 ;
      RECT 2.78 198.9 2.98 199.02 ;
      RECT 1.34 198.9 1.54 199.02 ;
      RECT 7.1 199.14 7.3 199.26 ;
      RECT 5.66 199.14 5.86 199.26 ;
      RECT 4.94 199.14 5.14 199.26 ;
      RECT 2.06 199.14 2.26 199.26 ;
      RECT 0.62 199.14 0.82 199.26 ;
      RECT 7.1 196.38 7.3 196.5 ;
      RECT 5.66 196.38 5.86 196.5 ;
      RECT 2.78 196.38 2.98 196.5 ;
      RECT 1.34 196.38 1.54 196.5 ;
      RECT 0.62 194.1 0.82 194.22 ;
      RECT 2.06 194.1 2.26 194.22 ;
      RECT 4.94 194.1 5.14 194.22 ;
      RECT 5.66 194.1 5.86 194.22 ;
      RECT 7.1 194.1 7.3 194.22 ;
      RECT 6.38 191.34 6.58 191.46 ;
      RECT 2.06 191.34 2.26 191.46 ;
      RECT 0.62 191.58 0.82 191.7 ;
      RECT 1.34 191.58 1.54 191.7 ;
      RECT 2.78 191.58 2.98 191.7 ;
      RECT 4.94 191.58 5.14 191.7 ;
      RECT 5.66 191.58 5.86 191.7 ;
      RECT 7.1 191.58 7.3 191.7 ;
      RECT 6.38 193.86 6.58 193.98 ;
      RECT 2.78 193.86 2.98 193.98 ;
      RECT 1.34 193.86 1.54 193.98 ;
      RECT 1.34 188.82 1.54 188.94 ;
      RECT 2.78 188.82 2.98 188.94 ;
      RECT 6.38 188.82 6.58 188.94 ;
      RECT 0.62 189.06 0.82 189.18 ;
      RECT 2.06 189.06 2.26 189.18 ;
      RECT 4.94 189.06 5.14 189.18 ;
      RECT 5.66 189.06 5.86 189.18 ;
      RECT 7.1 189.06 7.3 189.18 ;
      RECT 5.3 189.362 5.5 189.482 ;
      RECT 6.74 189.362 6.94 189.482 ;
      RECT 3.14 189.362 3.34 189.482 ;
      RECT 1.7 189.362 1.9 189.482 ;
      RECT 4.58 189.602 4.78 189.722 ;
      RECT 6.02 189.602 6.22 189.722 ;
      RECT 7.46 189.602 7.66 189.722 ;
      RECT 2.42 189.602 2.62 189.722 ;
      RECT 0.98 189.602 1.18 189.722 ;
      RECT 7.1 186.3 7.3 186.42 ;
      RECT 4.94 186.3 5.14 186.42 ;
      RECT 1.34 186.3 1.54 186.42 ;
      RECT 0.62 186.54 0.82 186.66 ;
      RECT 2.06 186.54 2.26 186.66 ;
      RECT 2.78 186.54 2.98 186.66 ;
      RECT 5.66 186.54 5.86 186.66 ;
      RECT 6.38 186.54 6.58 186.66 ;
      RECT 5.3 188.102 5.5 188.222 ;
      RECT 6.74 188.102 6.94 188.222 ;
      RECT 1.7 188.102 1.9 188.222 ;
      RECT 3.14 188.102 3.34 188.222 ;
      RECT 4.58 188.342 4.78 188.462 ;
      RECT 6.02 188.342 6.22 188.462 ;
      RECT 7.46 188.342 7.66 188.462 ;
      RECT 0.98 188.342 1.18 188.462 ;
      RECT 2.42 188.342 2.62 188.462 ;
      RECT 0.62 183.78 0.82 183.9 ;
      RECT 2.06 183.78 2.26 183.9 ;
      RECT 5.66 183.78 5.86 183.9 ;
      RECT 1.34 184.02 1.54 184.14 ;
      RECT 2.78 184.02 2.98 184.14 ;
      RECT 4.94 184.02 5.14 184.14 ;
      RECT 6.38 184.02 6.58 184.14 ;
      RECT 7.1 184.02 7.3 184.14 ;
      RECT 7.46 185.04 7.66 185.16 ;
      RECT 6.74 185.04 6.94 185.16 ;
      RECT 6.02 185.04 6.22 185.16 ;
      RECT 5.3 185.04 5.5 185.16 ;
      RECT 4.58 185.04 4.78 185.16 ;
      RECT 3.14 185.04 3.34 185.16 ;
      RECT 2.42 185.04 2.62 185.16 ;
      RECT 1.7 185.04 1.9 185.16 ;
      RECT 0.98 185.04 1.18 185.16 ;
      RECT 2.06 181.26 2.26 181.38 ;
      RECT 4.94 181.26 5.14 181.38 ;
      RECT 7.1 181.5 7.3 181.62 ;
      RECT 6.38 181.5 6.58 181.62 ;
      RECT 5.66 181.5 5.86 181.62 ;
      RECT 2.78 181.5 2.98 181.62 ;
      RECT 1.34 181.5 1.54 181.62 ;
      RECT 0.62 181.5 0.82 181.62 ;
      RECT 7.46 182.52 7.66 182.64 ;
      RECT 6.74 182.52 6.94 182.64 ;
      RECT 6.02 182.52 6.22 182.64 ;
      RECT 5.3 182.52 5.5 182.64 ;
      RECT 4.58 182.52 4.78 182.64 ;
      RECT 3.14 182.52 3.34 182.64 ;
      RECT 2.42 182.52 2.62 182.64 ;
      RECT 1.7 182.52 1.9 182.64 ;
      RECT 0.98 182.52 1.18 182.64 ;
      RECT 1.34 217.02 1.54 217.14 ;
      RECT 2.06 217.02 2.26 217.14 ;
      RECT 2.78 217.02 2.98 217.14 ;
      RECT 4.94 217.02 5.14 217.14 ;
      RECT 5.66 217.02 5.86 217.14 ;
      RECT 6.38 217.02 6.58 217.14 ;
      RECT 7.1 217.02 7.3 217.14 ;
      RECT 7.1 218.28 7.3 218.4 ;
      RECT 6.38 218.28 6.58 218.4 ;
      RECT 5.66 218.28 5.86 218.4 ;
      RECT 4.94 218.28 5.14 218.4 ;
      RECT 2.78 218.28 2.98 218.4 ;
      RECT 2.06 218.28 2.26 218.4 ;
      RECT 1.34 218.28 1.54 218.4 ;
      RECT 0.62 218.28 0.82 218.4 ;
      RECT 7.1 213.24 7.3 213.36 ;
      RECT 6.38 213.24 6.58 213.36 ;
      RECT 5.66 213.24 5.86 213.36 ;
      RECT 4.94 213.24 5.14 213.36 ;
      RECT 2.78 213.24 2.98 213.36 ;
      RECT 2.06 213.24 2.26 213.36 ;
      RECT 1.34 213.24 1.54 213.36 ;
      RECT 0.62 213.24 0.82 213.36 ;
      RECT 0.62 214.5 0.82 214.62 ;
      RECT 1.34 214.5 1.54 214.62 ;
      RECT 2.06 214.5 2.26 214.62 ;
      RECT 2.78 214.5 2.98 214.62 ;
      RECT 4.94 214.5 5.14 214.62 ;
      RECT 5.66 214.5 5.86 214.62 ;
      RECT 6.38 214.5 6.58 214.62 ;
      RECT 7.1 214.5 7.3 214.62 ;
      RECT 0.62 210.72 0.82 210.84 ;
      RECT 1.34 210.72 1.54 210.84 ;
      RECT 2.06 210.72 2.26 210.84 ;
      RECT 2.78 210.72 2.98 210.84 ;
      RECT 4.94 210.72 5.14 210.84 ;
      RECT 5.66 210.72 5.86 210.84 ;
      RECT 6.38 210.72 6.58 210.84 ;
      RECT 7.1 210.72 7.3 210.84 ;
      RECT 0.62 211.98 0.82 212.1 ;
      RECT 1.34 211.98 1.54 212.1 ;
      RECT 2.06 211.98 2.26 212.1 ;
      RECT 2.78 211.98 2.98 212.1 ;
      RECT 4.94 211.98 5.14 212.1 ;
      RECT 5.66 211.98 5.86 212.1 ;
      RECT 6.38 211.98 6.58 212.1 ;
      RECT 7.1 211.98 7.3 212.1 ;
      RECT 0.62 209.46 0.82 209.58 ;
      RECT 1.34 209.46 1.54 209.58 ;
      RECT 2.06 209.46 2.26 209.58 ;
      RECT 2.78 209.46 2.98 209.58 ;
      RECT 4.94 209.46 5.14 209.58 ;
      RECT 5.66 209.46 5.86 209.58 ;
      RECT 6.38 209.46 6.58 209.58 ;
      RECT 7.1 209.46 7.3 209.58 ;
      RECT 1.34 206.46 1.54 206.58 ;
      RECT 2.78 206.46 2.98 206.58 ;
      RECT 5.66 206.46 5.86 206.58 ;
      RECT 7.1 206.46 7.3 206.58 ;
      RECT 0.62 206.7 0.82 206.82 ;
      RECT 2.06 206.7 2.26 206.82 ;
      RECT 4.94 206.7 5.14 206.82 ;
      RECT 6.38 206.7 6.58 206.82 ;
      RECT 7.46 207.002 7.66 207.122 ;
      RECT 6.74 207.002 6.94 207.122 ;
      RECT 6.02 207.002 6.22 207.122 ;
      RECT 5.3 207.002 5.5 207.122 ;
      RECT 4.58 207.002 4.78 207.122 ;
      RECT 1.34 203.94 1.54 204.06 ;
      RECT 2.78 203.94 2.98 204.06 ;
      RECT 5.66 203.94 5.86 204.06 ;
      RECT 7.1 203.94 7.3 204.06 ;
      RECT 6.38 204.18 6.58 204.3 ;
      RECT 4.94 204.18 5.14 204.3 ;
      RECT 2.06 204.18 2.26 204.3 ;
      RECT 0.62 204.18 0.82 204.3 ;
      RECT 7.46 204.482 7.66 204.602 ;
      RECT 6.74 204.482 6.94 204.602 ;
      RECT 6.02 204.482 6.22 204.602 ;
      RECT 5.3 204.482 5.5 204.602 ;
      RECT 4.58 204.482 4.78 204.602 ;
      RECT 7.46 199.442 7.66 199.562 ;
      RECT 6.74 199.442 6.94 199.562 ;
      RECT 6.02 199.442 6.22 199.562 ;
      RECT 5.3 199.442 5.5 199.562 ;
      RECT 4.58 199.442 4.78 199.562 ;
      RECT 7.1 201.42 7.3 201.54 ;
      RECT 5.66 201.42 5.86 201.54 ;
      RECT 2.78 201.42 2.98 201.54 ;
      RECT 1.34 201.42 1.54 201.54 ;
      RECT 0.62 201.66 0.82 201.78 ;
      RECT 2.06 201.66 2.26 201.78 ;
      RECT 4.94 201.66 5.14 201.78 ;
      RECT 6.38 201.66 6.58 201.78 ;
      RECT 7.46 201.962 7.66 202.082 ;
      RECT 6.74 201.962 6.94 202.082 ;
      RECT 6.02 201.962 6.22 202.082 ;
      RECT 5.3 201.962 5.5 202.082 ;
      RECT 4.58 201.962 4.78 202.082 ;
      RECT 0.62 196.62 0.82 196.74 ;
      RECT 2.06 196.62 2.26 196.74 ;
      RECT 4.94 196.62 5.14 196.74 ;
      RECT 2.78 233.4 2.98 233.52 ;
      RECT 4.94 233.4 5.14 233.52 ;
      RECT 5.66 233.4 5.86 233.52 ;
      RECT 6.38 233.4 6.58 233.52 ;
      RECT 7.1 233.4 7.3 233.52 ;
      RECT 0.62 234.66 0.82 234.78 ;
      RECT 1.34 234.66 1.54 234.78 ;
      RECT 2.06 234.66 2.26 234.78 ;
      RECT 2.78 234.66 2.98 234.78 ;
      RECT 4.94 234.66 5.14 234.78 ;
      RECT 5.66 234.66 5.86 234.78 ;
      RECT 6.38 234.66 6.58 234.78 ;
      RECT 7.1 234.66 7.3 234.78 ;
      RECT 2.78 229.62 2.98 229.74 ;
      RECT 4.94 229.62 5.14 229.74 ;
      RECT 5.66 229.62 5.86 229.74 ;
      RECT 6.38 229.62 6.58 229.74 ;
      RECT 7.1 229.62 7.3 229.74 ;
      RECT 2.06 229.62 2.26 229.74 ;
      RECT 1.34 229.62 1.54 229.74 ;
      RECT 0.62 229.62 0.82 229.74 ;
      RECT 0.62 230.88 0.82 231 ;
      RECT 1.34 230.88 1.54 231 ;
      RECT 2.06 230.88 2.26 231 ;
      RECT 2.78 230.88 2.98 231 ;
      RECT 4.94 230.88 5.14 231 ;
      RECT 5.66 230.88 5.86 231 ;
      RECT 6.38 230.88 6.58 231 ;
      RECT 7.1 230.88 7.3 231 ;
      RECT 7.1 227.1 7.3 227.22 ;
      RECT 6.38 227.1 6.58 227.22 ;
      RECT 5.66 227.1 5.86 227.22 ;
      RECT 4.94 227.1 5.14 227.22 ;
      RECT 2.78 227.1 2.98 227.22 ;
      RECT 2.06 227.1 2.26 227.22 ;
      RECT 1.34 227.1 1.54 227.22 ;
      RECT 0.62 227.1 0.82 227.22 ;
      RECT 7.1 228.36 7.3 228.48 ;
      RECT 6.38 228.36 6.58 228.48 ;
      RECT 5.66 228.36 5.86 228.48 ;
      RECT 4.94 228.36 5.14 228.48 ;
      RECT 2.78 228.36 2.98 228.48 ;
      RECT 2.06 228.36 2.26 228.48 ;
      RECT 1.34 228.36 1.54 228.48 ;
      RECT 0.62 228.36 0.82 228.48 ;
      RECT 7.1 224.58 7.3 224.7 ;
      RECT 6.38 224.58 6.58 224.7 ;
      RECT 5.66 224.58 5.86 224.7 ;
      RECT 4.94 224.58 5.14 224.7 ;
      RECT 2.78 224.58 2.98 224.7 ;
      RECT 2.06 224.58 2.26 224.7 ;
      RECT 1.34 224.58 1.54 224.7 ;
      RECT 0.62 224.58 0.82 224.7 ;
      RECT 7.1 225.84 7.3 225.96 ;
      RECT 6.38 225.84 6.58 225.96 ;
      RECT 5.66 225.84 5.86 225.96 ;
      RECT 4.94 225.84 5.14 225.96 ;
      RECT 2.78 225.84 2.98 225.96 ;
      RECT 2.06 225.84 2.26 225.96 ;
      RECT 1.34 225.84 1.54 225.96 ;
      RECT 0.62 225.84 0.82 225.96 ;
      RECT 0.62 222.06 0.82 222.18 ;
      RECT 7.1 222.06 7.3 222.18 ;
      RECT 6.38 222.06 6.58 222.18 ;
      RECT 5.66 222.06 5.86 222.18 ;
      RECT 4.94 222.06 5.14 222.18 ;
      RECT 2.78 222.06 2.98 222.18 ;
      RECT 2.06 222.06 2.26 222.18 ;
      RECT 1.34 222.06 1.54 222.18 ;
      RECT 7.1 223.32 7.3 223.44 ;
      RECT 6.38 223.32 6.58 223.44 ;
      RECT 5.66 223.32 5.86 223.44 ;
      RECT 4.94 223.32 5.14 223.44 ;
      RECT 2.78 223.32 2.98 223.44 ;
      RECT 2.06 223.32 2.26 223.44 ;
      RECT 1.34 223.32 1.54 223.44 ;
      RECT 0.62 223.32 0.82 223.44 ;
      RECT 0.62 219.54 0.82 219.66 ;
      RECT 1.34 219.54 1.54 219.66 ;
      RECT 2.06 219.54 2.26 219.66 ;
      RECT 2.78 219.54 2.98 219.66 ;
      RECT 4.94 219.54 5.14 219.66 ;
      RECT 5.66 219.54 5.86 219.66 ;
      RECT 6.38 219.54 6.58 219.66 ;
      RECT 7.1 219.54 7.3 219.66 ;
      RECT 7.1 220.8 7.3 220.92 ;
      RECT 6.38 220.8 6.58 220.92 ;
      RECT 5.66 220.8 5.86 220.92 ;
      RECT 4.94 220.8 5.14 220.92 ;
      RECT 2.78 220.8 2.98 220.92 ;
      RECT 2.06 220.8 2.26 220.92 ;
      RECT 1.34 220.8 1.54 220.92 ;
      RECT 0.62 220.8 0.82 220.92 ;
      RECT 7.1 215.76 7.3 215.88 ;
      RECT 6.38 215.76 6.58 215.88 ;
      RECT 5.66 215.76 5.86 215.88 ;
      RECT 4.94 215.76 5.14 215.88 ;
      RECT 2.78 215.76 2.98 215.88 ;
      RECT 2.06 215.76 2.26 215.88 ;
      RECT 1.34 215.76 1.54 215.88 ;
      RECT 0.62 215.76 0.82 215.88 ;
      RECT 0.62 217.02 0.82 217.14 ;
      RECT 4.94 249.78 5.14 249.9 ;
      RECT 5.66 249.78 5.86 249.9 ;
      RECT 6.38 249.78 6.58 249.9 ;
      RECT 0.62 251.04 0.82 251.16 ;
      RECT 1.34 251.04 1.54 251.16 ;
      RECT 2.06 251.04 2.26 251.16 ;
      RECT 2.78 251.04 2.98 251.16 ;
      RECT 4.94 251.04 5.14 251.16 ;
      RECT 7.1 251.04 7.3 251.16 ;
      RECT 6.38 251.04 6.58 251.16 ;
      RECT 5.66 251.04 5.86 251.16 ;
      RECT 0.62 247.26 0.82 247.38 ;
      RECT 1.34 247.26 1.54 247.38 ;
      RECT 2.06 247.26 2.26 247.38 ;
      RECT 2.78 247.26 2.98 247.38 ;
      RECT 4.94 247.26 5.14 247.38 ;
      RECT 5.66 247.26 5.86 247.38 ;
      RECT 6.38 247.26 6.58 247.38 ;
      RECT 7.1 247.26 7.3 247.38 ;
      RECT 7.1 246 7.3 246.12 ;
      RECT 6.38 246 6.58 246.12 ;
      RECT 5.66 246 5.86 246.12 ;
      RECT 4.94 246 5.14 246.12 ;
      RECT 2.78 246 2.98 246.12 ;
      RECT 2.06 246 2.26 246.12 ;
      RECT 1.34 246 1.54 246.12 ;
      RECT 0.62 246 0.82 246.12 ;
      RECT 0.62 243.48 0.82 243.6 ;
      RECT 1.34 243.48 1.54 243.6 ;
      RECT 2.06 243.48 2.26 243.6 ;
      RECT 7.1 243.48 7.3 243.6 ;
      RECT 2.78 243.48 2.98 243.6 ;
      RECT 4.94 243.48 5.14 243.6 ;
      RECT 5.66 243.48 5.86 243.6 ;
      RECT 6.38 243.48 6.58 243.6 ;
      RECT 7.1 244.74 7.3 244.86 ;
      RECT 0.62 244.74 0.82 244.86 ;
      RECT 1.34 244.74 1.54 244.86 ;
      RECT 2.06 244.74 2.26 244.86 ;
      RECT 2.78 244.74 2.98 244.86 ;
      RECT 4.94 244.74 5.14 244.86 ;
      RECT 5.66 244.74 5.86 244.86 ;
      RECT 6.38 244.74 6.58 244.86 ;
      RECT 7.1 240.96 7.3 241.08 ;
      RECT 6.38 240.96 6.58 241.08 ;
      RECT 5.66 240.96 5.86 241.08 ;
      RECT 4.94 240.96 5.14 241.08 ;
      RECT 2.78 240.96 2.98 241.08 ;
      RECT 2.06 240.96 2.26 241.08 ;
      RECT 1.34 240.96 1.54 241.08 ;
      RECT 0.62 240.96 0.82 241.08 ;
      RECT 2.78 242.22 2.98 242.34 ;
      RECT 4.94 242.22 5.14 242.34 ;
      RECT 5.66 242.22 5.86 242.34 ;
      RECT 6.38 242.22 6.58 242.34 ;
      RECT 2.06 242.22 2.26 242.34 ;
      RECT 1.34 242.22 1.54 242.34 ;
      RECT 0.62 242.22 0.82 242.34 ;
      RECT 7.1 242.22 7.3 242.34 ;
      RECT 7.1 238.44 7.3 238.56 ;
      RECT 6.38 238.44 6.58 238.56 ;
      RECT 5.66 238.44 5.86 238.56 ;
      RECT 4.94 238.44 5.14 238.56 ;
      RECT 2.78 238.44 2.98 238.56 ;
      RECT 2.06 238.44 2.26 238.56 ;
      RECT 1.34 238.44 1.54 238.56 ;
      RECT 0.62 238.44 0.82 238.56 ;
      RECT 0.62 239.7 0.82 239.82 ;
      RECT 1.34 239.7 1.54 239.82 ;
      RECT 2.06 239.7 2.26 239.82 ;
      RECT 2.78 239.7 2.98 239.82 ;
      RECT 4.94 239.7 5.14 239.82 ;
      RECT 5.66 239.7 5.86 239.82 ;
      RECT 6.38 239.7 6.58 239.82 ;
      RECT 7.1 239.7 7.3 239.82 ;
      RECT 0.62 235.92 0.82 236.04 ;
      RECT 1.34 235.92 1.54 236.04 ;
      RECT 2.06 235.92 2.26 236.04 ;
      RECT 2.78 235.92 2.98 236.04 ;
      RECT 4.94 235.92 5.14 236.04 ;
      RECT 5.66 235.92 5.86 236.04 ;
      RECT 6.38 235.92 6.58 236.04 ;
      RECT 7.1 235.92 7.3 236.04 ;
      RECT 7.1 237.18 7.3 237.3 ;
      RECT 6.38 237.18 6.58 237.3 ;
      RECT 5.66 237.18 5.86 237.3 ;
      RECT 4.94 237.18 5.14 237.3 ;
      RECT 2.78 237.18 2.98 237.3 ;
      RECT 2.06 237.18 2.26 237.3 ;
      RECT 1.34 237.18 1.54 237.3 ;
      RECT 0.62 237.18 0.82 237.3 ;
      RECT 0.62 232.14 0.82 232.26 ;
      RECT 1.34 232.14 1.54 232.26 ;
      RECT 2.06 232.14 2.26 232.26 ;
      RECT 2.78 232.14 2.98 232.26 ;
      RECT 4.94 232.14 5.14 232.26 ;
      RECT 5.66 232.14 5.86 232.26 ;
      RECT 6.38 232.14 6.58 232.26 ;
      RECT 7.1 232.14 7.3 232.26 ;
      RECT 0.62 233.4 0.82 233.52 ;
      RECT 1.34 233.4 1.54 233.52 ;
      RECT 2.06 233.4 2.26 233.52 ;
      RECT 5.66 266.16 5.86 266.28 ;
      RECT 0.62 267.42 0.82 267.54 ;
      RECT 1.34 267.42 1.54 267.54 ;
      RECT 2.06 267.42 2.26 267.54 ;
      RECT 2.78 267.42 2.98 267.54 ;
      RECT 4.94 267.42 5.14 267.54 ;
      RECT 5.66 267.42 5.86 267.54 ;
      RECT 6.38 267.42 6.58 267.54 ;
      RECT 7.1 267.42 7.3 267.54 ;
      RECT 0.62 262.38 0.82 262.5 ;
      RECT 1.34 262.38 1.54 262.5 ;
      RECT 2.06 262.38 2.26 262.5 ;
      RECT 2.78 262.38 2.98 262.5 ;
      RECT 4.94 262.38 5.14 262.5 ;
      RECT 5.66 262.38 5.86 262.5 ;
      RECT 6.38 262.38 6.58 262.5 ;
      RECT 7.1 262.38 7.3 262.5 ;
      RECT 0.62 263.64 0.82 263.76 ;
      RECT 1.34 263.64 1.54 263.76 ;
      RECT 2.06 263.64 2.26 263.76 ;
      RECT 2.78 263.64 2.98 263.76 ;
      RECT 4.94 263.64 5.14 263.76 ;
      RECT 5.66 263.64 5.86 263.76 ;
      RECT 6.38 263.64 6.58 263.76 ;
      RECT 7.1 263.64 7.3 263.76 ;
      RECT 6.38 259.86 6.58 259.98 ;
      RECT 7.1 259.86 7.3 259.98 ;
      RECT 0.62 259.86 0.82 259.98 ;
      RECT 1.34 259.86 1.54 259.98 ;
      RECT 2.06 259.86 2.26 259.98 ;
      RECT 2.78 259.86 2.98 259.98 ;
      RECT 4.94 259.86 5.14 259.98 ;
      RECT 5.66 259.86 5.86 259.98 ;
      RECT 0.62 261.12 0.82 261.24 ;
      RECT 1.34 261.12 1.54 261.24 ;
      RECT 2.06 261.12 2.26 261.24 ;
      RECT 2.78 261.12 2.98 261.24 ;
      RECT 4.94 261.12 5.14 261.24 ;
      RECT 5.66 261.12 5.86 261.24 ;
      RECT 6.38 261.12 6.58 261.24 ;
      RECT 7.1 261.12 7.3 261.24 ;
      RECT 0.62 257.34 0.82 257.46 ;
      RECT 1.34 257.34 1.54 257.46 ;
      RECT 2.06 257.34 2.26 257.46 ;
      RECT 2.78 257.34 2.98 257.46 ;
      RECT 4.94 257.34 5.14 257.46 ;
      RECT 5.66 257.34 5.86 257.46 ;
      RECT 6.38 257.34 6.58 257.46 ;
      RECT 7.1 257.34 7.3 257.46 ;
      RECT 0.62 258.6 0.82 258.72 ;
      RECT 1.34 258.6 1.54 258.72 ;
      RECT 2.06 258.6 2.26 258.72 ;
      RECT 2.78 258.6 2.98 258.72 ;
      RECT 4.94 258.6 5.14 258.72 ;
      RECT 5.66 258.6 5.86 258.72 ;
      RECT 6.38 258.6 6.58 258.72 ;
      RECT 7.1 258.6 7.3 258.72 ;
      RECT 0.62 254.82 0.82 254.94 ;
      RECT 1.34 254.82 1.54 254.94 ;
      RECT 2.06 254.82 2.26 254.94 ;
      RECT 2.78 254.82 2.98 254.94 ;
      RECT 4.94 254.82 5.14 254.94 ;
      RECT 5.66 254.82 5.86 254.94 ;
      RECT 6.38 254.82 6.58 254.94 ;
      RECT 7.1 254.82 7.3 254.94 ;
      RECT 6.38 256.08 6.58 256.2 ;
      RECT 7.1 256.08 7.3 256.2 ;
      RECT 0.62 256.08 0.82 256.2 ;
      RECT 1.34 256.08 1.54 256.2 ;
      RECT 2.06 256.08 2.26 256.2 ;
      RECT 5.66 256.08 5.86 256.2 ;
      RECT 4.94 256.08 5.14 256.2 ;
      RECT 2.78 256.08 2.98 256.2 ;
      RECT 0.62 252.3 0.82 252.42 ;
      RECT 1.34 252.3 1.54 252.42 ;
      RECT 2.06 252.3 2.26 252.42 ;
      RECT 2.78 252.3 2.98 252.42 ;
      RECT 4.94 252.3 5.14 252.42 ;
      RECT 5.66 252.3 5.86 252.42 ;
      RECT 6.38 252.3 6.58 252.42 ;
      RECT 7.1 252.3 7.3 252.42 ;
      RECT 0.62 253.56 0.82 253.68 ;
      RECT 1.34 253.56 1.54 253.68 ;
      RECT 2.06 253.56 2.26 253.68 ;
      RECT 2.78 253.56 2.98 253.68 ;
      RECT 4.94 253.56 5.14 253.68 ;
      RECT 5.66 253.56 5.86 253.68 ;
      RECT 6.38 253.56 6.58 253.68 ;
      RECT 7.1 253.56 7.3 253.68 ;
      RECT 0.62 248.52 0.82 248.64 ;
      RECT 1.34 248.52 1.54 248.64 ;
      RECT 2.06 248.52 2.26 248.64 ;
      RECT 2.78 248.52 2.98 248.64 ;
      RECT 4.94 248.52 5.14 248.64 ;
      RECT 5.66 248.52 5.86 248.64 ;
      RECT 6.38 248.52 6.58 248.64 ;
      RECT 7.1 248.52 7.3 248.64 ;
      RECT 7.1 249.78 7.3 249.9 ;
      RECT 0.62 249.78 0.82 249.9 ;
      RECT 1.34 249.78 1.54 249.9 ;
      RECT 2.06 249.78 2.26 249.9 ;
      RECT 2.78 249.78 2.98 249.9 ;
      RECT 1.34 305.967 1.54 306.087 ;
      RECT 2.06 305.967 2.26 306.087 ;
      RECT 2.78 305.967 2.98 306.087 ;
      RECT 4.94 305.967 5.14 306.087 ;
      RECT 5.66 305.967 5.86 306.087 ;
      RECT 6.38 305.967 6.58 306.087 ;
      RECT 7.1 305.967 7.3 306.087 ;
      RECT 0.62 283.087 0.82 283.207 ;
      RECT 1.34 283.087 1.54 283.207 ;
      RECT 2.06 283.087 2.26 283.207 ;
      RECT 2.78 283.087 2.98 283.207 ;
      RECT 4.94 283.087 5.14 283.207 ;
      RECT 5.66 283.087 5.86 283.207 ;
      RECT 6.38 283.087 6.58 283.207 ;
      RECT 7.1 283.087 7.3 283.207 ;
      RECT 7.1 278.76 7.3 278.88 ;
      RECT 0.62 278.76 0.82 278.88 ;
      RECT 1.34 278.76 1.54 278.88 ;
      RECT 2.06 278.76 2.26 278.88 ;
      RECT 2.78 278.76 2.98 278.88 ;
      RECT 4.94 278.76 5.14 278.88 ;
      RECT 5.66 278.76 5.86 278.88 ;
      RECT 6.38 278.76 6.58 278.88 ;
      RECT 0.62 276.24 0.82 276.36 ;
      RECT 1.34 276.24 1.54 276.36 ;
      RECT 2.06 276.24 2.26 276.36 ;
      RECT 2.78 276.24 2.98 276.36 ;
      RECT 4.94 276.24 5.14 276.36 ;
      RECT 5.66 276.24 5.86 276.36 ;
      RECT 6.38 276.24 6.58 276.36 ;
      RECT 7.1 276.24 7.3 276.36 ;
      RECT 0.62 277.5 0.82 277.62 ;
      RECT 1.34 277.5 1.54 277.62 ;
      RECT 2.06 277.5 2.26 277.62 ;
      RECT 2.78 277.5 2.98 277.62 ;
      RECT 4.94 277.5 5.14 277.62 ;
      RECT 5.66 277.5 5.86 277.62 ;
      RECT 6.38 277.5 6.58 277.62 ;
      RECT 7.1 277.5 7.3 277.62 ;
      RECT 5.66 273.72 5.86 273.84 ;
      RECT 6.38 273.72 6.58 273.84 ;
      RECT 7.1 273.72 7.3 273.84 ;
      RECT 0.62 273.72 0.82 273.84 ;
      RECT 1.34 273.72 1.54 273.84 ;
      RECT 2.06 273.72 2.26 273.84 ;
      RECT 2.78 273.72 2.98 273.84 ;
      RECT 4.94 273.72 5.14 273.84 ;
      RECT 0.62 274.98 0.82 275.1 ;
      RECT 1.34 274.98 1.54 275.1 ;
      RECT 2.06 274.98 2.26 275.1 ;
      RECT 2.78 274.98 2.98 275.1 ;
      RECT 5.66 274.98 5.86 275.1 ;
      RECT 4.94 274.98 5.14 275.1 ;
      RECT 7.1 274.98 7.3 275.1 ;
      RECT 6.38 274.98 6.58 275.1 ;
      RECT 0.62 272.46 0.82 272.58 ;
      RECT 1.34 272.46 1.54 272.58 ;
      RECT 2.06 272.46 2.26 272.58 ;
      RECT 2.78 272.46 2.98 272.58 ;
      RECT 4.94 272.46 5.14 272.58 ;
      RECT 5.66 272.46 5.86 272.58 ;
      RECT 6.38 272.46 6.58 272.58 ;
      RECT 7.1 272.46 7.3 272.58 ;
      RECT 0.62 271.2 0.82 271.32 ;
      RECT 1.34 271.2 1.54 271.32 ;
      RECT 2.06 271.2 2.26 271.32 ;
      RECT 2.78 271.2 2.98 271.32 ;
      RECT 4.94 271.2 5.14 271.32 ;
      RECT 5.66 271.2 5.86 271.32 ;
      RECT 6.38 271.2 6.58 271.32 ;
      RECT 7.1 271.2 7.3 271.32 ;
      RECT 6.38 268.68 6.58 268.8 ;
      RECT 7.1 268.68 7.3 268.8 ;
      RECT 0.62 268.68 0.82 268.8 ;
      RECT 1.34 268.68 1.54 268.8 ;
      RECT 2.06 268.68 2.26 268.8 ;
      RECT 2.78 268.68 2.98 268.8 ;
      RECT 4.94 268.68 5.14 268.8 ;
      RECT 5.66 268.68 5.86 268.8 ;
      RECT 0.62 269.94 0.82 270.06 ;
      RECT 1.34 269.94 1.54 270.06 ;
      RECT 2.06 269.94 2.26 270.06 ;
      RECT 2.78 269.94 2.98 270.06 ;
      RECT 4.94 269.94 5.14 270.06 ;
      RECT 5.66 269.94 5.86 270.06 ;
      RECT 6.38 269.94 6.58 270.06 ;
      RECT 7.1 269.94 7.3 270.06 ;
      RECT 0.62 264.9 0.82 265.02 ;
      RECT 1.34 264.9 1.54 265.02 ;
      RECT 2.06 264.9 2.26 265.02 ;
      RECT 2.78 264.9 2.98 265.02 ;
      RECT 4.94 264.9 5.14 265.02 ;
      RECT 5.66 264.9 5.86 265.02 ;
      RECT 6.38 264.9 6.58 265.02 ;
      RECT 7.1 264.9 7.3 265.02 ;
      RECT 7.1 266.16 7.3 266.28 ;
      RECT 6.38 266.16 6.58 266.28 ;
      RECT 0.62 266.16 0.82 266.28 ;
      RECT 1.34 266.16 1.54 266.28 ;
      RECT 2.06 266.16 2.26 266.28 ;
      RECT 2.78 266.16 2.98 266.28 ;
      RECT 4.94 266.16 5.14 266.28 ;
      RECT 9.26 131.578 9.46 131.698 ;
      RECT 9.98 133.38 10.18 133.5 ;
      RECT 13.58 133.38 13.78 133.5 ;
      RECT 15.02 133.38 15.22 133.5 ;
      RECT 14.3 133.62 14.5 133.74 ;
      RECT 12.86 133.62 13.06 133.74 ;
      RECT 11.42 133.62 11.62 133.74 ;
      RECT 10.7 133.62 10.9 133.74 ;
      RECT 9.26 133.62 9.46 133.74 ;
      RECT 11.42 128.34 11.62 128.46 ;
      RECT 13.58 128.34 13.78 128.46 ;
      RECT 15.02 128.34 15.22 128.46 ;
      RECT 9.98 128.34 10.18 128.46 ;
      RECT 9.26 128.58 9.46 128.7 ;
      RECT 10.7 128.58 10.9 128.7 ;
      RECT 12.86 128.58 13.06 128.7 ;
      RECT 14.3 128.58 14.5 128.7 ;
      RECT 14.3 129.058 14.5 129.178 ;
      RECT 12.86 129.058 13.06 129.178 ;
      RECT 10.7 129.058 10.9 129.178 ;
      RECT 9.26 129.058 9.46 129.178 ;
      RECT 15.02 129.298 15.22 129.418 ;
      RECT 13.58 129.298 13.78 129.418 ;
      RECT 11.42 129.298 11.62 129.418 ;
      RECT 9.98 129.298 10.18 129.418 ;
      RECT 15.02 130.86 15.22 130.98 ;
      RECT 13.58 130.86 13.78 130.98 ;
      RECT 11.42 130.86 11.62 130.98 ;
      RECT 9.98 130.86 10.18 130.98 ;
      RECT 14.3 125.82 14.5 125.94 ;
      RECT 12.86 125.82 13.06 125.94 ;
      RECT 9.98 125.82 10.18 125.94 ;
      RECT 15.02 126.06 15.22 126.18 ;
      RECT 13.58 126.06 13.78 126.18 ;
      RECT 11.42 126.06 11.62 126.18 ;
      RECT 10.7 126.06 10.9 126.18 ;
      RECT 9.26 126.06 9.46 126.18 ;
      RECT 15.02 126.538 15.22 126.658 ;
      RECT 14.3 126.538 14.5 126.658 ;
      RECT 13.58 126.538 13.78 126.658 ;
      RECT 12.86 126.538 13.06 126.658 ;
      RECT 11.42 126.538 11.62 126.658 ;
      RECT 10.7 126.538 10.9 126.658 ;
      RECT 9.98 126.538 10.18 126.658 ;
      RECT 9.26 126.538 9.46 126.658 ;
      RECT 15.02 123.3 15.22 123.42 ;
      RECT 12.86 123.3 13.06 123.42 ;
      RECT 10.7 123.3 10.9 123.42 ;
      RECT 14.3 123.54 14.5 123.66 ;
      RECT 13.58 123.54 13.78 123.66 ;
      RECT 11.42 123.54 11.62 123.66 ;
      RECT 9.98 123.54 10.18 123.66 ;
      RECT 9.26 123.54 9.46 123.66 ;
      RECT 15.02 124.018 15.22 124.138 ;
      RECT 14.3 124.018 14.5 124.138 ;
      RECT 13.58 124.018 13.78 124.138 ;
      RECT 12.86 124.018 13.06 124.138 ;
      RECT 11.42 124.018 11.62 124.138 ;
      RECT 10.7 124.018 10.9 124.138 ;
      RECT 9.98 124.018 10.18 124.138 ;
      RECT 9.26 124.018 9.46 124.138 ;
      RECT 13.58 120.78 13.78 120.9 ;
      RECT 9.98 120.78 10.18 120.9 ;
      RECT 14.3 120.78 14.5 120.9 ;
      RECT 11.42 121.02 11.62 121.14 ;
      RECT 10.7 121.02 10.9 121.14 ;
      RECT 9.26 121.02 9.46 121.14 ;
      RECT 15.02 121.02 15.22 121.14 ;
      RECT 12.86 121.02 13.06 121.14 ;
      RECT 15.02 121.498 15.22 121.618 ;
      RECT 14.3 121.498 14.5 121.618 ;
      RECT 13.58 121.498 13.78 121.618 ;
      RECT 12.86 121.498 13.06 121.618 ;
      RECT 11.42 121.498 11.62 121.618 ;
      RECT 10.7 121.498 10.9 121.618 ;
      RECT 9.98 121.498 10.18 121.618 ;
      RECT 9.26 121.498 9.46 121.618 ;
      RECT 9.98 118.26 10.18 118.38 ;
      RECT 11.42 118.26 11.62 118.38 ;
      RECT 13.58 118.26 13.78 118.38 ;
      RECT 15.02 118.26 15.22 118.38 ;
      RECT 9.26 118.5 9.46 118.62 ;
      RECT 10.7 118.5 10.9 118.62 ;
      RECT 12.86 118.5 13.06 118.62 ;
      RECT 14.3 118.5 14.5 118.62 ;
      RECT 15.02 118.978 15.22 119.098 ;
      RECT 14.3 118.978 14.5 119.098 ;
      RECT 13.58 118.978 13.78 119.098 ;
      RECT 12.86 118.978 13.06 119.098 ;
      RECT 11.42 118.978 11.62 119.098 ;
      RECT 10.7 118.978 10.9 119.098 ;
      RECT 9.98 118.978 10.18 119.098 ;
      RECT 9.26 118.978 9.46 119.098 ;
      RECT 7.1 325.9425 7.3 326.0625 ;
      RECT 6.38 325.9425 6.58 326.0625 ;
      RECT 5.66 325.9425 5.86 326.0625 ;
      RECT 4.94 325.9425 5.14 326.0625 ;
      RECT 2.78 325.9425 2.98 326.0625 ;
      RECT 2.06 325.9425 2.26 326.0625 ;
      RECT 1.34 325.9425 1.54 326.0625 ;
      RECT 0.62 325.9425 0.82 326.0625 ;
      RECT 0.62 305.967 0.82 306.087 ;
      RECT 10.7 158.82 10.9 158.94 ;
      RECT 9.98 158.82 10.18 158.94 ;
      RECT 14.3 158.82 14.5 158.94 ;
      RECT 9.26 156.06 9.46 156.18 ;
      RECT 10.7 156.06 10.9 156.18 ;
      RECT 12.86 156.06 13.06 156.18 ;
      RECT 14.3 156.06 14.5 156.18 ;
      RECT 15.02 156.3 15.22 156.42 ;
      RECT 13.58 156.3 13.78 156.42 ;
      RECT 11.42 156.3 11.62 156.42 ;
      RECT 9.98 156.3 10.18 156.42 ;
      RECT 9.26 153.54 9.46 153.66 ;
      RECT 10.7 153.54 10.9 153.66 ;
      RECT 14.3 153.54 14.5 153.66 ;
      RECT 15.02 153.78 15.22 153.9 ;
      RECT 13.58 153.78 13.78 153.9 ;
      RECT 12.86 153.78 13.06 153.9 ;
      RECT 11.42 153.78 11.62 153.9 ;
      RECT 9.98 153.78 10.18 153.9 ;
      RECT 10.7 148.5 10.9 148.62 ;
      RECT 11.42 148.5 11.62 148.62 ;
      RECT 15.02 148.5 15.22 148.62 ;
      RECT 14.3 148.74 14.5 148.86 ;
      RECT 13.58 148.74 13.78 148.86 ;
      RECT 12.86 148.74 13.06 148.86 ;
      RECT 9.98 148.74 10.18 148.86 ;
      RECT 9.26 148.74 9.46 148.86 ;
      RECT 15.02 145.98 15.22 146.1 ;
      RECT 14.3 145.98 14.5 146.1 ;
      RECT 13.58 145.98 13.78 146.1 ;
      RECT 12.86 145.98 13.06 146.1 ;
      RECT 11.42 145.98 11.62 146.1 ;
      RECT 10.7 145.98 10.9 146.1 ;
      RECT 9.98 145.98 10.18 146.1 ;
      RECT 9.26 145.98 9.46 146.1 ;
      RECT 9.26 143.7 9.46 143.82 ;
      RECT 10.7 143.7 10.9 143.82 ;
      RECT 12.86 143.7 13.06 143.82 ;
      RECT 14.3 143.7 14.5 143.82 ;
      RECT 9.98 143.46 10.18 143.58 ;
      RECT 11.42 143.46 11.62 143.58 ;
      RECT 13.58 143.46 13.78 143.58 ;
      RECT 15.02 143.46 15.22 143.58 ;
      RECT 9.98 140.94 10.18 141.06 ;
      RECT 15.02 140.94 15.22 141.06 ;
      RECT 11.42 140.94 11.62 141.06 ;
      RECT 9.26 141.18 9.46 141.3 ;
      RECT 10.7 141.18 10.9 141.3 ;
      RECT 12.86 141.18 13.06 141.3 ;
      RECT 13.58 141.18 13.78 141.3 ;
      RECT 14.3 141.18 14.5 141.3 ;
      RECT 15.02 136.618 15.22 136.738 ;
      RECT 14.3 136.618 14.5 136.738 ;
      RECT 13.58 136.618 13.78 136.738 ;
      RECT 12.86 136.618 13.06 136.738 ;
      RECT 11.42 136.618 11.62 136.738 ;
      RECT 10.7 136.618 10.9 136.738 ;
      RECT 9.98 136.618 10.18 136.738 ;
      RECT 9.26 136.618 9.46 136.738 ;
      RECT 9.26 138.42 9.46 138.54 ;
      RECT 10.7 138.42 10.9 138.54 ;
      RECT 12.86 138.42 13.06 138.54 ;
      RECT 14.3 138.42 14.5 138.54 ;
      RECT 15.02 138.66 15.22 138.78 ;
      RECT 13.58 138.66 13.78 138.78 ;
      RECT 11.42 138.66 11.62 138.78 ;
      RECT 9.98 138.66 10.18 138.78 ;
      RECT 15.02 139.138 15.22 139.258 ;
      RECT 14.3 139.138 14.5 139.258 ;
      RECT 13.58 139.138 13.78 139.258 ;
      RECT 12.86 139.138 13.06 139.258 ;
      RECT 11.42 139.138 11.62 139.258 ;
      RECT 10.7 139.138 10.9 139.258 ;
      RECT 9.98 139.138 10.18 139.258 ;
      RECT 9.26 139.138 9.46 139.258 ;
      RECT 15.02 134.098 15.22 134.218 ;
      RECT 14.3 134.098 14.5 134.218 ;
      RECT 13.58 134.098 13.78 134.218 ;
      RECT 12.86 134.098 13.06 134.218 ;
      RECT 11.42 134.098 11.62 134.218 ;
      RECT 10.7 134.098 10.9 134.218 ;
      RECT 9.98 134.098 10.18 134.218 ;
      RECT 9.26 134.098 9.46 134.218 ;
      RECT 9.98 135.9 10.18 136.02 ;
      RECT 11.42 135.9 11.62 136.02 ;
      RECT 13.58 135.9 13.78 136.02 ;
      RECT 15.02 135.9 15.22 136.02 ;
      RECT 9.26 136.14 9.46 136.26 ;
      RECT 10.7 136.14 10.9 136.26 ;
      RECT 12.86 136.14 13.06 136.26 ;
      RECT 14.3 136.14 14.5 136.26 ;
      RECT 9.26 131.1 9.46 131.22 ;
      RECT 10.7 131.1 10.9 131.22 ;
      RECT 12.86 131.1 13.06 131.22 ;
      RECT 14.3 131.1 14.5 131.22 ;
      RECT 15.02 131.578 15.22 131.698 ;
      RECT 14.3 131.578 14.5 131.698 ;
      RECT 13.58 131.578 13.78 131.698 ;
      RECT 12.86 131.578 13.06 131.698 ;
      RECT 11.42 131.578 11.62 131.698 ;
      RECT 10.7 131.578 10.9 131.698 ;
      RECT 9.98 131.578 10.18 131.698 ;
      RECT 8.9 180 9.1 180.12 ;
      RECT 15.38 174.96 15.58 175.08 ;
      RECT 14.66 174.96 14.86 175.08 ;
      RECT 13.94 174.96 14.14 175.08 ;
      RECT 13.22 174.96 13.42 175.08 ;
      RECT 11.06 174.96 11.26 175.08 ;
      RECT 10.34 174.96 10.54 175.08 ;
      RECT 9.62 174.96 9.82 175.08 ;
      RECT 8.9 174.96 9.1 175.08 ;
      RECT 9.98 176.22 10.18 176.34 ;
      RECT 11.42 176.22 11.62 176.34 ;
      RECT 13.58 176.22 13.78 176.34 ;
      RECT 9.26 176.46 9.46 176.58 ;
      RECT 10.7 176.46 10.9 176.58 ;
      RECT 12.86 176.46 13.06 176.58 ;
      RECT 14.3 176.46 14.5 176.58 ;
      RECT 15.02 176.46 15.22 176.58 ;
      RECT 15.38 177.48 15.58 177.6 ;
      RECT 14.66 177.48 14.86 177.6 ;
      RECT 13.94 177.48 14.14 177.6 ;
      RECT 13.22 177.48 13.42 177.6 ;
      RECT 11.06 177.48 11.26 177.6 ;
      RECT 10.34 177.48 10.54 177.6 ;
      RECT 9.62 177.48 9.82 177.6 ;
      RECT 8.9 177.48 9.1 177.6 ;
      RECT 15.38 172.44 15.58 172.56 ;
      RECT 14.66 172.44 14.86 172.56 ;
      RECT 13.94 172.44 14.14 172.56 ;
      RECT 13.22 172.44 13.42 172.56 ;
      RECT 11.06 172.44 11.26 172.56 ;
      RECT 10.34 172.44 10.54 172.56 ;
      RECT 9.62 172.44 9.82 172.56 ;
      RECT 8.9 172.44 9.1 172.56 ;
      RECT 9.98 173.7 10.18 173.82 ;
      RECT 12.86 173.7 13.06 173.82 ;
      RECT 9.26 173.94 9.46 174.06 ;
      RECT 10.7 173.94 10.9 174.06 ;
      RECT 11.42 173.94 11.62 174.06 ;
      RECT 13.58 173.94 13.78 174.06 ;
      RECT 14.3 173.94 14.5 174.06 ;
      RECT 15.02 173.94 15.22 174.06 ;
      RECT 15.38 169.92 15.58 170.04 ;
      RECT 14.66 169.92 14.86 170.04 ;
      RECT 13.94 169.92 14.14 170.04 ;
      RECT 13.22 169.92 13.42 170.04 ;
      RECT 11.06 169.92 11.26 170.04 ;
      RECT 10.34 169.92 10.54 170.04 ;
      RECT 9.62 169.92 9.82 170.04 ;
      RECT 8.9 169.92 9.1 170.04 ;
      RECT 15.02 171.18 15.22 171.3 ;
      RECT 11.42 171.18 11.62 171.3 ;
      RECT 9.98 171.18 10.18 171.3 ;
      RECT 9.26 171.42 9.46 171.54 ;
      RECT 10.7 171.42 10.9 171.54 ;
      RECT 12.86 171.42 13.06 171.54 ;
      RECT 13.58 171.42 13.78 171.54 ;
      RECT 14.3 171.42 14.5 171.54 ;
      RECT 15.38 167.4 15.58 167.52 ;
      RECT 14.66 167.4 14.86 167.52 ;
      RECT 13.94 167.4 14.14 167.52 ;
      RECT 13.22 167.4 13.42 167.52 ;
      RECT 11.06 167.4 11.26 167.52 ;
      RECT 10.34 167.4 10.54 167.52 ;
      RECT 9.62 167.4 9.82 167.52 ;
      RECT 8.9 167.4 9.1 167.52 ;
      RECT 13.58 168.66 13.78 168.78 ;
      RECT 9.26 168.66 9.46 168.78 ;
      RECT 9.98 168.9 10.18 169.02 ;
      RECT 10.7 168.9 10.9 169.02 ;
      RECT 11.42 168.9 11.62 169.02 ;
      RECT 12.86 168.9 13.06 169.02 ;
      RECT 14.3 168.9 14.5 169.02 ;
      RECT 15.02 168.9 15.22 169.02 ;
      RECT 9.26 163.86 9.46 163.98 ;
      RECT 10.7 163.86 10.9 163.98 ;
      RECT 11.42 163.86 11.62 163.98 ;
      RECT 13.58 163.86 13.78 163.98 ;
      RECT 15.02 163.86 15.22 163.98 ;
      RECT 15.38 164.88 15.58 165 ;
      RECT 14.66 164.88 14.86 165 ;
      RECT 13.94 164.88 14.14 165 ;
      RECT 13.22 164.88 13.42 165 ;
      RECT 11.06 164.88 11.26 165 ;
      RECT 10.34 164.88 10.54 165 ;
      RECT 9.62 164.88 9.82 165 ;
      RECT 8.9 164.88 9.1 165 ;
      RECT 9.98 166.14 10.18 166.26 ;
      RECT 12.86 166.14 13.06 166.26 ;
      RECT 14.3 166.14 14.5 166.26 ;
      RECT 9.26 166.38 9.46 166.5 ;
      RECT 10.7 166.38 10.9 166.5 ;
      RECT 11.42 166.38 11.62 166.5 ;
      RECT 13.58 166.38 13.78 166.5 ;
      RECT 15.02 166.38 15.22 166.5 ;
      RECT 14.3 163.62 14.5 163.74 ;
      RECT 12.86 163.62 13.06 163.74 ;
      RECT 9.98 163.62 10.18 163.74 ;
      RECT 9.26 158.58 9.46 158.7 ;
      RECT 11.42 158.58 11.62 158.7 ;
      RECT 13.58 158.58 13.78 158.7 ;
      RECT 15.02 158.58 15.22 158.7 ;
      RECT 12.86 158.82 13.06 158.94 ;
      RECT 14.3 199.14 14.5 199.26 ;
      RECT 13.58 199.14 13.78 199.26 ;
      RECT 11.42 199.14 11.62 199.26 ;
      RECT 9.98 199.14 10.18 199.26 ;
      RECT 13.58 196.38 13.78 196.5 ;
      RECT 11.42 196.38 11.62 196.5 ;
      RECT 9.98 196.38 10.18 196.5 ;
      RECT 9.26 194.1 9.46 194.22 ;
      RECT 10.7 194.1 10.9 194.22 ;
      RECT 12.86 194.1 13.06 194.22 ;
      RECT 14.3 194.1 14.5 194.22 ;
      RECT 13.58 191.34 13.78 191.46 ;
      RECT 10.7 191.34 10.9 191.46 ;
      RECT 9.26 191.34 9.46 191.46 ;
      RECT 9.98 191.58 10.18 191.7 ;
      RECT 11.42 191.58 11.62 191.7 ;
      RECT 12.86 191.58 13.06 191.7 ;
      RECT 14.3 191.58 14.5 191.7 ;
      RECT 15.02 191.58 15.22 191.7 ;
      RECT 15.02 193.86 15.22 193.98 ;
      RECT 13.58 193.86 13.78 193.98 ;
      RECT 11.42 193.86 11.62 193.98 ;
      RECT 9.98 193.86 10.18 193.98 ;
      RECT 9.26 188.82 9.46 188.94 ;
      RECT 10.7 188.82 10.9 188.94 ;
      RECT 12.86 188.82 13.06 188.94 ;
      RECT 15.02 188.82 15.22 188.94 ;
      RECT 9.98 189.06 10.18 189.18 ;
      RECT 11.42 189.06 11.62 189.18 ;
      RECT 13.58 189.06 13.78 189.18 ;
      RECT 14.3 189.06 14.5 189.18 ;
      RECT 13.22 189.362 13.42 189.482 ;
      RECT 14.66 189.362 14.86 189.482 ;
      RECT 9.62 189.362 9.82 189.482 ;
      RECT 11.06 189.362 11.26 189.482 ;
      RECT 13.94 189.602 14.14 189.722 ;
      RECT 15.38 189.602 15.58 189.722 ;
      RECT 8.9 189.602 9.1 189.722 ;
      RECT 10.34 189.602 10.54 189.722 ;
      RECT 15.02 186.3 15.22 186.42 ;
      RECT 11.42 186.3 11.62 186.42 ;
      RECT 9.98 186.3 10.18 186.42 ;
      RECT 9.26 186.54 9.46 186.66 ;
      RECT 10.7 186.54 10.9 186.66 ;
      RECT 12.86 186.54 13.06 186.66 ;
      RECT 13.58 186.54 13.78 186.66 ;
      RECT 14.3 186.54 14.5 186.66 ;
      RECT 14.66 188.102 14.86 188.222 ;
      RECT 13.22 188.102 13.42 188.222 ;
      RECT 9.62 188.102 9.82 188.222 ;
      RECT 11.06 188.102 11.26 188.222 ;
      RECT 15.38 188.342 15.58 188.462 ;
      RECT 13.94 188.342 14.14 188.462 ;
      RECT 8.9 188.342 9.1 188.462 ;
      RECT 10.34 188.342 10.54 188.462 ;
      RECT 9.26 183.78 9.46 183.9 ;
      RECT 10.7 183.78 10.9 183.9 ;
      RECT 14.3 183.78 14.5 183.9 ;
      RECT 9.98 184.02 10.18 184.14 ;
      RECT 11.42 184.02 11.62 184.14 ;
      RECT 12.86 184.02 13.06 184.14 ;
      RECT 13.58 184.02 13.78 184.14 ;
      RECT 15.02 184.02 15.22 184.14 ;
      RECT 15.38 185.04 15.58 185.16 ;
      RECT 14.66 185.04 14.86 185.16 ;
      RECT 13.94 185.04 14.14 185.16 ;
      RECT 13.22 185.04 13.42 185.16 ;
      RECT 11.06 185.04 11.26 185.16 ;
      RECT 10.34 185.04 10.54 185.16 ;
      RECT 9.62 185.04 9.82 185.16 ;
      RECT 8.9 185.04 9.1 185.16 ;
      RECT 9.26 181.26 9.46 181.38 ;
      RECT 11.42 181.26 11.62 181.38 ;
      RECT 13.58 181.26 13.78 181.38 ;
      RECT 15.02 181.26 15.22 181.38 ;
      RECT 14.3 181.5 14.5 181.62 ;
      RECT 12.86 181.5 13.06 181.62 ;
      RECT 10.7 181.5 10.9 181.62 ;
      RECT 9.98 181.5 10.18 181.62 ;
      RECT 15.38 182.52 15.58 182.64 ;
      RECT 14.66 182.52 14.86 182.64 ;
      RECT 13.94 182.52 14.14 182.64 ;
      RECT 13.22 182.52 13.42 182.64 ;
      RECT 11.06 182.52 11.26 182.64 ;
      RECT 10.34 182.52 10.54 182.64 ;
      RECT 9.62 182.52 9.82 182.64 ;
      RECT 8.9 182.52 9.1 182.64 ;
      RECT 9.98 178.74 10.18 178.86 ;
      RECT 11.42 178.74 11.62 178.86 ;
      RECT 13.58 178.74 13.78 178.86 ;
      RECT 9.26 178.98 9.46 179.1 ;
      RECT 15.02 178.98 15.22 179.1 ;
      RECT 14.3 178.98 14.5 179.1 ;
      RECT 12.86 178.98 13.06 179.1 ;
      RECT 10.7 178.98 10.9 179.1 ;
      RECT 15.38 180 15.58 180.12 ;
      RECT 14.66 180 14.86 180.12 ;
      RECT 13.94 180 14.14 180.12 ;
      RECT 13.22 180 13.42 180.12 ;
      RECT 11.06 180 11.26 180.12 ;
      RECT 10.34 180 10.54 180.12 ;
      RECT 9.62 180 9.82 180.12 ;
      RECT 11.42 214.5 11.62 214.62 ;
      RECT 12.86 214.5 13.06 214.62 ;
      RECT 13.58 214.5 13.78 214.62 ;
      RECT 14.3 214.5 14.5 214.62 ;
      RECT 15.02 214.5 15.22 214.62 ;
      RECT 9.26 210.72 9.46 210.84 ;
      RECT 9.98 210.72 10.18 210.84 ;
      RECT 10.7 210.72 10.9 210.84 ;
      RECT 11.42 210.72 11.62 210.84 ;
      RECT 12.86 210.72 13.06 210.84 ;
      RECT 13.58 210.72 13.78 210.84 ;
      RECT 14.3 210.72 14.5 210.84 ;
      RECT 15.02 210.72 15.22 210.84 ;
      RECT 9.26 211.98 9.46 212.1 ;
      RECT 9.98 211.98 10.18 212.1 ;
      RECT 10.7 211.98 10.9 212.1 ;
      RECT 11.42 211.98 11.62 212.1 ;
      RECT 12.86 211.98 13.06 212.1 ;
      RECT 13.58 211.98 13.78 212.1 ;
      RECT 14.3 211.98 14.5 212.1 ;
      RECT 15.02 211.98 15.22 212.1 ;
      RECT 9.26 209.46 9.46 209.58 ;
      RECT 9.98 209.46 10.18 209.58 ;
      RECT 10.7 209.46 10.9 209.58 ;
      RECT 11.42 209.46 11.62 209.58 ;
      RECT 12.86 209.46 13.06 209.58 ;
      RECT 13.58 209.46 13.78 209.58 ;
      RECT 14.3 209.46 14.5 209.58 ;
      RECT 15.02 209.46 15.22 209.58 ;
      RECT 9.98 206.46 10.18 206.58 ;
      RECT 11.42 206.46 11.62 206.58 ;
      RECT 13.58 206.46 13.78 206.58 ;
      RECT 15.02 206.46 15.22 206.58 ;
      RECT 9.26 206.7 9.46 206.82 ;
      RECT 10.7 206.7 10.9 206.82 ;
      RECT 12.86 206.7 13.06 206.82 ;
      RECT 14.3 206.7 14.5 206.82 ;
      RECT 15.38 207.002 15.58 207.122 ;
      RECT 14.66 207.002 14.86 207.122 ;
      RECT 13.94 207.002 14.14 207.122 ;
      RECT 13.22 207.002 13.42 207.122 ;
      RECT 11.06 207.002 11.26 207.122 ;
      RECT 10.34 207.002 10.54 207.122 ;
      RECT 9.62 207.002 9.82 207.122 ;
      RECT 8.9 207.002 9.1 207.122 ;
      RECT 9.98 203.94 10.18 204.06 ;
      RECT 11.42 203.94 11.62 204.06 ;
      RECT 13.58 203.94 13.78 204.06 ;
      RECT 15.02 203.94 15.22 204.06 ;
      RECT 14.3 204.18 14.5 204.3 ;
      RECT 12.86 204.18 13.06 204.3 ;
      RECT 10.7 204.18 10.9 204.3 ;
      RECT 9.26 204.18 9.46 204.3 ;
      RECT 15.38 204.482 15.58 204.602 ;
      RECT 14.66 204.482 14.86 204.602 ;
      RECT 13.94 204.482 14.14 204.602 ;
      RECT 13.22 204.482 13.42 204.602 ;
      RECT 11.06 204.482 11.26 204.602 ;
      RECT 10.34 204.482 10.54 204.602 ;
      RECT 9.62 204.482 9.82 204.602 ;
      RECT 8.9 204.482 9.1 204.602 ;
      RECT 15.38 199.442 15.58 199.562 ;
      RECT 14.66 199.442 14.86 199.562 ;
      RECT 13.94 199.442 14.14 199.562 ;
      RECT 13.22 199.442 13.42 199.562 ;
      RECT 11.06 199.442 11.26 199.562 ;
      RECT 10.34 199.442 10.54 199.562 ;
      RECT 9.62 199.442 9.82 199.562 ;
      RECT 8.9 199.442 9.1 199.562 ;
      RECT 15.02 201.42 15.22 201.54 ;
      RECT 13.58 201.42 13.78 201.54 ;
      RECT 11.42 201.42 11.62 201.54 ;
      RECT 9.98 201.42 10.18 201.54 ;
      RECT 9.26 201.66 9.46 201.78 ;
      RECT 10.7 201.66 10.9 201.78 ;
      RECT 12.86 201.66 13.06 201.78 ;
      RECT 14.3 201.66 14.5 201.78 ;
      RECT 15.38 201.962 15.58 202.082 ;
      RECT 14.66 201.962 14.86 202.082 ;
      RECT 13.94 201.962 14.14 202.082 ;
      RECT 13.22 201.962 13.42 202.082 ;
      RECT 11.06 201.962 11.26 202.082 ;
      RECT 10.34 201.962 10.54 202.082 ;
      RECT 9.62 201.962 9.82 202.082 ;
      RECT 8.9 201.962 9.1 202.082 ;
      RECT 9.26 196.62 9.46 196.74 ;
      RECT 10.7 196.62 10.9 196.74 ;
      RECT 12.86 196.62 13.06 196.74 ;
      RECT 14.3 196.62 14.5 196.74 ;
      RECT 15.02 196.62 15.22 196.74 ;
      RECT 15.38 196.922 15.58 197.042 ;
      RECT 14.66 196.922 14.86 197.042 ;
      RECT 13.94 196.922 14.14 197.042 ;
      RECT 13.22 196.922 13.42 197.042 ;
      RECT 11.06 196.922 11.26 197.042 ;
      RECT 10.34 196.922 10.54 197.042 ;
      RECT 9.62 196.922 9.82 197.042 ;
      RECT 8.9 196.922 9.1 197.042 ;
      RECT 15.02 198.9 15.22 199.02 ;
      RECT 12.86 198.9 13.06 199.02 ;
      RECT 10.7 198.9 10.9 199.02 ;
      RECT 9.26 198.9 9.46 199.02 ;
      RECT 13.58 230.88 13.78 231 ;
      RECT 14.3 230.88 14.5 231 ;
      RECT 15.02 230.88 15.22 231 ;
      RECT 15.02 227.1 15.22 227.22 ;
      RECT 14.3 227.1 14.5 227.22 ;
      RECT 13.58 227.1 13.78 227.22 ;
      RECT 12.86 227.1 13.06 227.22 ;
      RECT 11.42 227.1 11.62 227.22 ;
      RECT 10.7 227.1 10.9 227.22 ;
      RECT 9.98 227.1 10.18 227.22 ;
      RECT 9.26 227.1 9.46 227.22 ;
      RECT 15.02 228.36 15.22 228.48 ;
      RECT 14.3 228.36 14.5 228.48 ;
      RECT 13.58 228.36 13.78 228.48 ;
      RECT 12.86 228.36 13.06 228.48 ;
      RECT 11.42 228.36 11.62 228.48 ;
      RECT 10.7 228.36 10.9 228.48 ;
      RECT 9.98 228.36 10.18 228.48 ;
      RECT 9.26 228.36 9.46 228.48 ;
      RECT 15.02 224.58 15.22 224.7 ;
      RECT 14.3 224.58 14.5 224.7 ;
      RECT 13.58 224.58 13.78 224.7 ;
      RECT 12.86 224.58 13.06 224.7 ;
      RECT 11.42 224.58 11.62 224.7 ;
      RECT 10.7 224.58 10.9 224.7 ;
      RECT 9.98 224.58 10.18 224.7 ;
      RECT 9.26 224.58 9.46 224.7 ;
      RECT 15.02 225.84 15.22 225.96 ;
      RECT 14.3 225.84 14.5 225.96 ;
      RECT 13.58 225.84 13.78 225.96 ;
      RECT 12.86 225.84 13.06 225.96 ;
      RECT 11.42 225.84 11.62 225.96 ;
      RECT 10.7 225.84 10.9 225.96 ;
      RECT 9.98 225.84 10.18 225.96 ;
      RECT 9.26 225.84 9.46 225.96 ;
      RECT 15.02 222.06 15.22 222.18 ;
      RECT 14.3 222.06 14.5 222.18 ;
      RECT 13.58 222.06 13.78 222.18 ;
      RECT 12.86 222.06 13.06 222.18 ;
      RECT 11.42 222.06 11.62 222.18 ;
      RECT 10.7 222.06 10.9 222.18 ;
      RECT 9.98 222.06 10.18 222.18 ;
      RECT 9.26 222.06 9.46 222.18 ;
      RECT 9.98 223.32 10.18 223.44 ;
      RECT 9.26 223.32 9.46 223.44 ;
      RECT 15.02 223.32 15.22 223.44 ;
      RECT 14.3 223.32 14.5 223.44 ;
      RECT 13.58 223.32 13.78 223.44 ;
      RECT 12.86 223.32 13.06 223.44 ;
      RECT 11.42 223.32 11.62 223.44 ;
      RECT 10.7 223.32 10.9 223.44 ;
      RECT 9.26 219.54 9.46 219.66 ;
      RECT 9.98 219.54 10.18 219.66 ;
      RECT 10.7 219.54 10.9 219.66 ;
      RECT 11.42 219.54 11.62 219.66 ;
      RECT 12.86 219.54 13.06 219.66 ;
      RECT 13.58 219.54 13.78 219.66 ;
      RECT 14.3 219.54 14.5 219.66 ;
      RECT 15.02 219.54 15.22 219.66 ;
      RECT 15.02 220.8 15.22 220.92 ;
      RECT 14.3 220.8 14.5 220.92 ;
      RECT 13.58 220.8 13.78 220.92 ;
      RECT 12.86 220.8 13.06 220.92 ;
      RECT 11.42 220.8 11.62 220.92 ;
      RECT 10.7 220.8 10.9 220.92 ;
      RECT 9.98 220.8 10.18 220.92 ;
      RECT 9.26 220.8 9.46 220.92 ;
      RECT 15.02 215.76 15.22 215.88 ;
      RECT 14.3 215.76 14.5 215.88 ;
      RECT 13.58 215.76 13.78 215.88 ;
      RECT 12.86 215.76 13.06 215.88 ;
      RECT 11.42 215.76 11.62 215.88 ;
      RECT 10.7 215.76 10.9 215.88 ;
      RECT 9.98 215.76 10.18 215.88 ;
      RECT 9.26 215.76 9.46 215.88 ;
      RECT 9.26 217.02 9.46 217.14 ;
      RECT 9.98 217.02 10.18 217.14 ;
      RECT 10.7 217.02 10.9 217.14 ;
      RECT 11.42 217.02 11.62 217.14 ;
      RECT 12.86 217.02 13.06 217.14 ;
      RECT 13.58 217.02 13.78 217.14 ;
      RECT 14.3 217.02 14.5 217.14 ;
      RECT 15.02 217.02 15.22 217.14 ;
      RECT 15.02 218.28 15.22 218.4 ;
      RECT 14.3 218.28 14.5 218.4 ;
      RECT 13.58 218.28 13.78 218.4 ;
      RECT 12.86 218.28 13.06 218.4 ;
      RECT 11.42 218.28 11.62 218.4 ;
      RECT 10.7 218.28 10.9 218.4 ;
      RECT 9.98 218.28 10.18 218.4 ;
      RECT 9.26 218.28 9.46 218.4 ;
      RECT 15.02 213.24 15.22 213.36 ;
      RECT 14.3 213.24 14.5 213.36 ;
      RECT 13.58 213.24 13.78 213.36 ;
      RECT 12.86 213.24 13.06 213.36 ;
      RECT 11.42 213.24 11.62 213.36 ;
      RECT 10.7 213.24 10.9 213.36 ;
      RECT 9.98 213.24 10.18 213.36 ;
      RECT 9.26 213.24 9.46 213.36 ;
      RECT 9.26 214.5 9.46 214.62 ;
      RECT 9.98 214.5 10.18 214.62 ;
      RECT 10.7 214.5 10.9 214.62 ;
      RECT 13.58 246 13.78 246.12 ;
      RECT 9.26 243.48 9.46 243.6 ;
      RECT 9.98 243.48 10.18 243.6 ;
      RECT 10.7 243.48 10.9 243.6 ;
      RECT 11.42 243.48 11.62 243.6 ;
      RECT 12.86 243.48 13.06 243.6 ;
      RECT 13.58 243.48 13.78 243.6 ;
      RECT 14.3 243.48 14.5 243.6 ;
      RECT 15.02 243.48 15.22 243.6 ;
      RECT 9.98 244.74 10.18 244.86 ;
      RECT 9.26 244.74 9.46 244.86 ;
      RECT 10.7 244.74 10.9 244.86 ;
      RECT 11.42 244.74 11.62 244.86 ;
      RECT 12.86 244.74 13.06 244.86 ;
      RECT 13.58 244.74 13.78 244.86 ;
      RECT 14.3 244.74 14.5 244.86 ;
      RECT 15.02 244.74 15.22 244.86 ;
      RECT 9.26 240.96 9.46 241.08 ;
      RECT 9.98 240.96 10.18 241.08 ;
      RECT 10.7 240.96 10.9 241.08 ;
      RECT 11.42 240.96 11.62 241.08 ;
      RECT 12.86 240.96 13.06 241.08 ;
      RECT 13.58 240.96 13.78 241.08 ;
      RECT 14.3 240.96 14.5 241.08 ;
      RECT 15.02 240.96 15.22 241.08 ;
      RECT 15.02 242.22 15.22 242.34 ;
      RECT 9.26 242.22 9.46 242.34 ;
      RECT 9.98 242.22 10.18 242.34 ;
      RECT 10.7 242.22 10.9 242.34 ;
      RECT 14.3 242.22 14.5 242.34 ;
      RECT 13.58 242.22 13.78 242.34 ;
      RECT 12.86 242.22 13.06 242.34 ;
      RECT 11.42 242.22 11.62 242.34 ;
      RECT 15.02 238.44 15.22 238.56 ;
      RECT 14.3 238.44 14.5 238.56 ;
      RECT 13.58 238.44 13.78 238.56 ;
      RECT 12.86 238.44 13.06 238.56 ;
      RECT 11.42 238.44 11.62 238.56 ;
      RECT 10.7 238.44 10.9 238.56 ;
      RECT 9.98 238.44 10.18 238.56 ;
      RECT 9.26 238.44 9.46 238.56 ;
      RECT 12.86 239.7 13.06 239.82 ;
      RECT 13.58 239.7 13.78 239.82 ;
      RECT 14.3 239.7 14.5 239.82 ;
      RECT 15.02 239.7 15.22 239.82 ;
      RECT 11.42 239.7 11.62 239.82 ;
      RECT 10.7 239.7 10.9 239.82 ;
      RECT 9.98 239.7 10.18 239.82 ;
      RECT 9.26 239.7 9.46 239.82 ;
      RECT 9.26 235.92 9.46 236.04 ;
      RECT 9.98 235.92 10.18 236.04 ;
      RECT 10.7 235.92 10.9 236.04 ;
      RECT 11.42 235.92 11.62 236.04 ;
      RECT 12.86 235.92 13.06 236.04 ;
      RECT 13.58 235.92 13.78 236.04 ;
      RECT 14.3 235.92 14.5 236.04 ;
      RECT 15.02 235.92 15.22 236.04 ;
      RECT 15.02 237.18 15.22 237.3 ;
      RECT 14.3 237.18 14.5 237.3 ;
      RECT 13.58 237.18 13.78 237.3 ;
      RECT 12.86 237.18 13.06 237.3 ;
      RECT 10.7 237.18 10.9 237.3 ;
      RECT 11.42 237.18 11.62 237.3 ;
      RECT 9.98 237.18 10.18 237.3 ;
      RECT 9.26 237.18 9.46 237.3 ;
      RECT 9.26 232.14 9.46 232.26 ;
      RECT 9.98 232.14 10.18 232.26 ;
      RECT 10.7 232.14 10.9 232.26 ;
      RECT 11.42 232.14 11.62 232.26 ;
      RECT 12.86 232.14 13.06 232.26 ;
      RECT 13.58 232.14 13.78 232.26 ;
      RECT 14.3 232.14 14.5 232.26 ;
      RECT 15.02 232.14 15.22 232.26 ;
      RECT 9.26 233.4 9.46 233.52 ;
      RECT 9.98 233.4 10.18 233.52 ;
      RECT 10.7 233.4 10.9 233.52 ;
      RECT 11.42 233.4 11.62 233.52 ;
      RECT 12.86 233.4 13.06 233.52 ;
      RECT 13.58 233.4 13.78 233.52 ;
      RECT 14.3 233.4 14.5 233.52 ;
      RECT 15.02 233.4 15.22 233.52 ;
      RECT 9.26 234.66 9.46 234.78 ;
      RECT 9.98 234.66 10.18 234.78 ;
      RECT 10.7 234.66 10.9 234.78 ;
      RECT 11.42 234.66 11.62 234.78 ;
      RECT 12.86 234.66 13.06 234.78 ;
      RECT 13.58 234.66 13.78 234.78 ;
      RECT 14.3 234.66 14.5 234.78 ;
      RECT 15.02 234.66 15.22 234.78 ;
      RECT 12.86 229.62 13.06 229.74 ;
      RECT 13.58 229.62 13.78 229.74 ;
      RECT 14.3 229.62 14.5 229.74 ;
      RECT 15.02 229.62 15.22 229.74 ;
      RECT 9.26 229.62 9.46 229.74 ;
      RECT 9.98 229.62 10.18 229.74 ;
      RECT 10.7 229.62 10.9 229.74 ;
      RECT 11.42 229.62 11.62 229.74 ;
      RECT 9.26 230.88 9.46 231 ;
      RECT 9.98 230.88 10.18 231 ;
      RECT 10.7 230.88 10.9 231 ;
      RECT 11.42 230.88 11.62 231 ;
      RECT 12.86 230.88 13.06 231 ;
      RECT 9.98 259.86 10.18 259.98 ;
      RECT 10.7 259.86 10.9 259.98 ;
      RECT 11.42 259.86 11.62 259.98 ;
      RECT 12.86 259.86 13.06 259.98 ;
      RECT 13.58 259.86 13.78 259.98 ;
      RECT 14.3 259.86 14.5 259.98 ;
      RECT 15.02 259.86 15.22 259.98 ;
      RECT 9.26 261.12 9.46 261.24 ;
      RECT 9.98 261.12 10.18 261.24 ;
      RECT 10.7 261.12 10.9 261.24 ;
      RECT 11.42 261.12 11.62 261.24 ;
      RECT 12.86 261.12 13.06 261.24 ;
      RECT 13.58 261.12 13.78 261.24 ;
      RECT 14.3 261.12 14.5 261.24 ;
      RECT 15.02 261.12 15.22 261.24 ;
      RECT 9.26 257.34 9.46 257.46 ;
      RECT 9.98 257.34 10.18 257.46 ;
      RECT 10.7 257.34 10.9 257.46 ;
      RECT 11.42 257.34 11.62 257.46 ;
      RECT 12.86 257.34 13.06 257.46 ;
      RECT 13.58 257.34 13.78 257.46 ;
      RECT 14.3 257.34 14.5 257.46 ;
      RECT 15.02 257.34 15.22 257.46 ;
      RECT 10.7 258.6 10.9 258.72 ;
      RECT 9.98 258.6 10.18 258.72 ;
      RECT 11.42 258.6 11.62 258.72 ;
      RECT 15.02 258.6 15.22 258.72 ;
      RECT 9.26 258.6 9.46 258.72 ;
      RECT 12.86 258.6 13.06 258.72 ;
      RECT 13.58 258.6 13.78 258.72 ;
      RECT 14.3 258.6 14.5 258.72 ;
      RECT 15.02 254.82 15.22 254.94 ;
      RECT 9.26 254.82 9.46 254.94 ;
      RECT 9.98 254.82 10.18 254.94 ;
      RECT 10.7 254.82 10.9 254.94 ;
      RECT 11.42 254.82 11.62 254.94 ;
      RECT 12.86 254.82 13.06 254.94 ;
      RECT 13.58 254.82 13.78 254.94 ;
      RECT 14.3 254.82 14.5 254.94 ;
      RECT 9.26 256.08 9.46 256.2 ;
      RECT 9.98 256.08 10.18 256.2 ;
      RECT 10.7 256.08 10.9 256.2 ;
      RECT 11.42 256.08 11.62 256.2 ;
      RECT 12.86 256.08 13.06 256.2 ;
      RECT 13.58 256.08 13.78 256.2 ;
      RECT 14.3 256.08 14.5 256.2 ;
      RECT 15.02 256.08 15.22 256.2 ;
      RECT 14.3 252.3 14.5 252.42 ;
      RECT 13.58 252.3 13.78 252.42 ;
      RECT 15.02 252.3 15.22 252.42 ;
      RECT 9.26 252.3 9.46 252.42 ;
      RECT 9.98 252.3 10.18 252.42 ;
      RECT 10.7 252.3 10.9 252.42 ;
      RECT 11.42 252.3 11.62 252.42 ;
      RECT 12.86 252.3 13.06 252.42 ;
      RECT 9.26 253.56 9.46 253.68 ;
      RECT 9.98 253.56 10.18 253.68 ;
      RECT 10.7 253.56 10.9 253.68 ;
      RECT 11.42 253.56 11.62 253.68 ;
      RECT 12.86 253.56 13.06 253.68 ;
      RECT 13.58 253.56 13.78 253.68 ;
      RECT 14.3 253.56 14.5 253.68 ;
      RECT 15.02 253.56 15.22 253.68 ;
      RECT 9.26 248.52 9.46 248.64 ;
      RECT 9.98 248.52 10.18 248.64 ;
      RECT 10.7 248.52 10.9 248.64 ;
      RECT 11.42 248.52 11.62 248.64 ;
      RECT 12.86 248.52 13.06 248.64 ;
      RECT 13.58 248.52 13.78 248.64 ;
      RECT 14.3 248.52 14.5 248.64 ;
      RECT 15.02 248.52 15.22 248.64 ;
      RECT 9.26 249.78 9.46 249.9 ;
      RECT 9.98 249.78 10.18 249.9 ;
      RECT 10.7 249.78 10.9 249.9 ;
      RECT 11.42 249.78 11.62 249.9 ;
      RECT 12.86 249.78 13.06 249.9 ;
      RECT 13.58 249.78 13.78 249.9 ;
      RECT 14.3 249.78 14.5 249.9 ;
      RECT 15.02 249.78 15.22 249.9 ;
      RECT 9.26 251.04 9.46 251.16 ;
      RECT 9.98 251.04 10.18 251.16 ;
      RECT 10.7 251.04 10.9 251.16 ;
      RECT 11.42 251.04 11.62 251.16 ;
      RECT 12.86 251.04 13.06 251.16 ;
      RECT 13.58 251.04 13.78 251.16 ;
      RECT 14.3 251.04 14.5 251.16 ;
      RECT 15.02 251.04 15.22 251.16 ;
      RECT 10.7 247.26 10.9 247.38 ;
      RECT 11.42 247.26 11.62 247.38 ;
      RECT 12.86 247.26 13.06 247.38 ;
      RECT 13.58 247.26 13.78 247.38 ;
      RECT 14.3 247.26 14.5 247.38 ;
      RECT 15.02 247.26 15.22 247.38 ;
      RECT 9.26 247.26 9.46 247.38 ;
      RECT 9.98 247.26 10.18 247.38 ;
      RECT 9.26 246 9.46 246.12 ;
      RECT 9.98 246 10.18 246.12 ;
      RECT 10.7 246 10.9 246.12 ;
      RECT 11.42 246 11.62 246.12 ;
      RECT 12.86 246 13.06 246.12 ;
      RECT 15.02 246 15.22 246.12 ;
      RECT 14.3 246 14.5 246.12 ;
      RECT 11.42 276.24 11.62 276.36 ;
      RECT 12.86 276.24 13.06 276.36 ;
      RECT 13.58 276.24 13.78 276.36 ;
      RECT 14.3 276.24 14.5 276.36 ;
      RECT 15.02 276.24 15.22 276.36 ;
      RECT 9.26 277.5 9.46 277.62 ;
      RECT 9.98 277.5 10.18 277.62 ;
      RECT 10.7 277.5 10.9 277.62 ;
      RECT 11.42 277.5 11.62 277.62 ;
      RECT 12.86 277.5 13.06 277.62 ;
      RECT 13.58 277.5 13.78 277.62 ;
      RECT 14.3 277.5 14.5 277.62 ;
      RECT 15.02 277.5 15.22 277.62 ;
      RECT 9.26 273.72 9.46 273.84 ;
      RECT 9.98 273.72 10.18 273.84 ;
      RECT 10.7 273.72 10.9 273.84 ;
      RECT 11.42 273.72 11.62 273.84 ;
      RECT 12.86 273.72 13.06 273.84 ;
      RECT 13.58 273.72 13.78 273.84 ;
      RECT 14.3 273.72 14.5 273.84 ;
      RECT 15.02 273.72 15.22 273.84 ;
      RECT 9.26 274.98 9.46 275.1 ;
      RECT 9.98 274.98 10.18 275.1 ;
      RECT 10.7 274.98 10.9 275.1 ;
      RECT 11.42 274.98 11.62 275.1 ;
      RECT 12.86 274.98 13.06 275.1 ;
      RECT 13.58 274.98 13.78 275.1 ;
      RECT 14.3 274.98 14.5 275.1 ;
      RECT 15.02 274.98 15.22 275.1 ;
      RECT 9.26 272.46 9.46 272.58 ;
      RECT 9.98 272.46 10.18 272.58 ;
      RECT 10.7 272.46 10.9 272.58 ;
      RECT 11.42 272.46 11.62 272.58 ;
      RECT 12.86 272.46 13.06 272.58 ;
      RECT 13.58 272.46 13.78 272.58 ;
      RECT 14.3 272.46 14.5 272.58 ;
      RECT 15.02 272.46 15.22 272.58 ;
      RECT 9.26 271.2 9.46 271.32 ;
      RECT 9.98 271.2 10.18 271.32 ;
      RECT 10.7 271.2 10.9 271.32 ;
      RECT 11.42 271.2 11.62 271.32 ;
      RECT 12.86 271.2 13.06 271.32 ;
      RECT 13.58 271.2 13.78 271.32 ;
      RECT 14.3 271.2 14.5 271.32 ;
      RECT 15.02 271.2 15.22 271.32 ;
      RECT 9.26 268.68 9.46 268.8 ;
      RECT 9.98 268.68 10.18 268.8 ;
      RECT 10.7 268.68 10.9 268.8 ;
      RECT 11.42 268.68 11.62 268.8 ;
      RECT 12.86 268.68 13.06 268.8 ;
      RECT 13.58 268.68 13.78 268.8 ;
      RECT 14.3 268.68 14.5 268.8 ;
      RECT 15.02 268.68 15.22 268.8 ;
      RECT 15.02 269.94 15.22 270.06 ;
      RECT 14.3 269.94 14.5 270.06 ;
      RECT 9.26 269.94 9.46 270.06 ;
      RECT 9.98 269.94 10.18 270.06 ;
      RECT 10.7 269.94 10.9 270.06 ;
      RECT 11.42 269.94 11.62 270.06 ;
      RECT 12.86 269.94 13.06 270.06 ;
      RECT 13.58 269.94 13.78 270.06 ;
      RECT 9.26 264.9 9.46 265.02 ;
      RECT 9.98 264.9 10.18 265.02 ;
      RECT 10.7 264.9 10.9 265.02 ;
      RECT 11.42 264.9 11.62 265.02 ;
      RECT 12.86 264.9 13.06 265.02 ;
      RECT 13.58 264.9 13.78 265.02 ;
      RECT 14.3 264.9 14.5 265.02 ;
      RECT 15.02 264.9 15.22 265.02 ;
      RECT 9.26 266.16 9.46 266.28 ;
      RECT 9.98 266.16 10.18 266.28 ;
      RECT 10.7 266.16 10.9 266.28 ;
      RECT 11.42 266.16 11.62 266.28 ;
      RECT 12.86 266.16 13.06 266.28 ;
      RECT 13.58 266.16 13.78 266.28 ;
      RECT 14.3 266.16 14.5 266.28 ;
      RECT 15.02 266.16 15.22 266.28 ;
      RECT 9.26 267.42 9.46 267.54 ;
      RECT 9.98 267.42 10.18 267.54 ;
      RECT 10.7 267.42 10.9 267.54 ;
      RECT 11.42 267.42 11.62 267.54 ;
      RECT 12.86 267.42 13.06 267.54 ;
      RECT 13.58 267.42 13.78 267.54 ;
      RECT 14.3 267.42 14.5 267.54 ;
      RECT 15.02 267.42 15.22 267.54 ;
      RECT 9.26 262.38 9.46 262.5 ;
      RECT 9.98 262.38 10.18 262.5 ;
      RECT 10.7 262.38 10.9 262.5 ;
      RECT 11.42 262.38 11.62 262.5 ;
      RECT 12.86 262.38 13.06 262.5 ;
      RECT 13.58 262.38 13.78 262.5 ;
      RECT 14.3 262.38 14.5 262.5 ;
      RECT 15.02 262.38 15.22 262.5 ;
      RECT 9.26 263.64 9.46 263.76 ;
      RECT 9.98 263.64 10.18 263.76 ;
      RECT 10.7 263.64 10.9 263.76 ;
      RECT 11.42 263.64 11.62 263.76 ;
      RECT 12.86 263.64 13.06 263.76 ;
      RECT 13.58 263.64 13.78 263.76 ;
      RECT 14.3 263.64 14.5 263.76 ;
      RECT 15.02 263.64 15.22 263.76 ;
      RECT 9.26 259.86 9.46 259.98 ;
      RECT 19.34 131.578 19.54 131.698 ;
      RECT 20.06 131.578 20.26 131.698 ;
      RECT 17.9 131.1 18.1 131.22 ;
      RECT 17.18 131.1 17.38 131.22 ;
      RECT 19.34 131.1 19.54 131.22 ;
      RECT 18.62 130.86 18.82 130.98 ;
      RECT 20.06 130.86 20.26 130.98 ;
      RECT 18.26 129.84 18.46 129.96 ;
      RECT 19.7 129.6 19.9 129.72 ;
      RECT 17.18 129.298 17.38 129.418 ;
      RECT 18.62 129.298 18.82 129.418 ;
      RECT 20.06 129.298 20.26 129.418 ;
      RECT 17.9 129.058 18.1 129.178 ;
      RECT 19.34 129.058 19.54 129.178 ;
      RECT 18.62 128.58 18.82 128.7 ;
      RECT 17.9 128.58 18.1 128.7 ;
      RECT 17.18 128.58 17.38 128.7 ;
      RECT 20.06 128.34 20.26 128.46 ;
      RECT 19.34 128.34 19.54 128.46 ;
      RECT 18.26 127.32 18.46 127.44 ;
      RECT 19.7 127.08 19.9 127.2 ;
      RECT 17.18 126.538 17.38 126.658 ;
      RECT 17.9 126.538 18.1 126.658 ;
      RECT 18.62 126.538 18.82 126.658 ;
      RECT 19.34 126.538 19.54 126.658 ;
      RECT 20.06 126.538 20.26 126.658 ;
      RECT 17.18 126.06 17.38 126.18 ;
      RECT 19.34 126.06 19.54 126.18 ;
      RECT 17.9 125.82 18.1 125.94 ;
      RECT 18.62 125.82 18.82 125.94 ;
      RECT 20.06 125.82 20.26 125.94 ;
      RECT 18.26 124.8 18.46 124.92 ;
      RECT 19.7 124.56 19.9 124.68 ;
      RECT 17.18 124.018 17.38 124.138 ;
      RECT 17.9 124.018 18.1 124.138 ;
      RECT 18.62 124.018 18.82 124.138 ;
      RECT 19.34 124.018 19.54 124.138 ;
      RECT 20.06 124.018 20.26 124.138 ;
      RECT 17.9 123.54 18.1 123.66 ;
      RECT 19.34 123.54 19.54 123.66 ;
      RECT 20.06 123.54 20.26 123.66 ;
      RECT 17.18 123.3 17.38 123.42 ;
      RECT 18.62 123.3 18.82 123.42 ;
      RECT 18.26 122.28 18.46 122.4 ;
      RECT 19.7 122.04 19.9 122.16 ;
      RECT 17.18 121.498 17.38 121.618 ;
      RECT 17.9 121.498 18.1 121.618 ;
      RECT 18.62 121.498 18.82 121.618 ;
      RECT 19.34 121.498 19.54 121.618 ;
      RECT 20.06 121.498 20.26 121.618 ;
      RECT 17.18 121.02 17.38 121.14 ;
      RECT 17.9 121.02 18.1 121.14 ;
      RECT 19.34 121.02 19.54 121.14 ;
      RECT 18.62 120.78 18.82 120.9 ;
      RECT 20.06 120.78 20.26 120.9 ;
      RECT 18.26 119.76 18.46 119.88 ;
      RECT 19.7 119.52 19.9 119.64 ;
      RECT 17.18 118.978 17.38 119.098 ;
      RECT 17.9 118.978 18.1 119.098 ;
      RECT 18.62 118.978 18.82 119.098 ;
      RECT 19.34 118.978 19.54 119.098 ;
      RECT 20.06 118.978 20.26 119.098 ;
      RECT 20.06 118.5 20.26 118.62 ;
      RECT 18.62 118.5 18.82 118.62 ;
      RECT 17.18 118.5 17.38 118.62 ;
      RECT 19.34 118.26 19.54 118.38 ;
      RECT 17.9 118.26 18.1 118.38 ;
      RECT 15.02 325.9425 15.22 326.0625 ;
      RECT 14.3 325.9425 14.5 326.0625 ;
      RECT 13.58 325.9425 13.78 326.0625 ;
      RECT 12.86 325.9425 13.06 326.0625 ;
      RECT 11.42 325.9425 11.62 326.0625 ;
      RECT 10.7 325.9425 10.9 326.0625 ;
      RECT 9.98 325.9425 10.18 326.0625 ;
      RECT 9.26 325.9425 9.46 326.0625 ;
      RECT 9.26 305.967 9.46 306.087 ;
      RECT 9.98 305.967 10.18 306.087 ;
      RECT 10.7 305.967 10.9 306.087 ;
      RECT 11.42 305.967 11.62 306.087 ;
      RECT 12.86 305.967 13.06 306.087 ;
      RECT 13.58 305.967 13.78 306.087 ;
      RECT 14.3 305.967 14.5 306.087 ;
      RECT 15.02 305.967 15.22 306.087 ;
      RECT 9.26 283.087 9.46 283.207 ;
      RECT 9.98 283.087 10.18 283.207 ;
      RECT 10.7 283.087 10.9 283.207 ;
      RECT 11.42 283.087 11.62 283.207 ;
      RECT 12.86 283.087 13.06 283.207 ;
      RECT 13.58 283.087 13.78 283.207 ;
      RECT 14.3 283.087 14.5 283.207 ;
      RECT 15.02 283.087 15.22 283.207 ;
      RECT 9.26 278.76 9.46 278.88 ;
      RECT 9.98 278.76 10.18 278.88 ;
      RECT 10.7 278.76 10.9 278.88 ;
      RECT 11.42 278.76 11.62 278.88 ;
      RECT 12.86 278.76 13.06 278.88 ;
      RECT 13.58 278.76 13.78 278.88 ;
      RECT 14.3 278.76 14.5 278.88 ;
      RECT 15.02 278.76 15.22 278.88 ;
      RECT 9.26 276.24 9.46 276.36 ;
      RECT 9.98 276.24 10.18 276.36 ;
      RECT 10.7 276.24 10.9 276.36 ;
      RECT 19.7 164.88 19.9 165 ;
      RECT 20.06 163.86 20.26 163.98 ;
      RECT 19.34 163.86 19.54 163.98 ;
      RECT 17.9 163.86 18.1 163.98 ;
      RECT 17.18 163.86 17.38 163.98 ;
      RECT 18.62 163.62 18.82 163.74 ;
      RECT 19.7 162.6 19.9 162.72 ;
      RECT 18.26 162.6 18.46 162.72 ;
      RECT 19.7 160.08 19.9 160.2 ;
      RECT 18.26 159.84 18.46 159.96 ;
      RECT 17.18 158.82 17.38 158.94 ;
      RECT 18.62 158.82 18.82 158.94 ;
      RECT 19.34 158.82 19.54 158.94 ;
      RECT 20.06 158.58 20.26 158.7 ;
      RECT 17.9 158.58 18.1 158.7 ;
      RECT 20.42 158.278 20.62 158.398 ;
      RECT 17.54 158.278 17.74 158.398 ;
      RECT 18.98 158.038 19.18 158.158 ;
      RECT 19.7 157.56 19.9 157.68 ;
      RECT 18.26 157.32 18.46 157.44 ;
      RECT 18.98 156.842 19.18 156.962 ;
      RECT 17.54 156.842 17.74 156.962 ;
      RECT 20.42 156.602 20.62 156.722 ;
      RECT 17.9 156.3 18.1 156.42 ;
      RECT 19.34 156.3 19.54 156.42 ;
      RECT 20.06 156.3 20.26 156.42 ;
      RECT 17.18 156.06 17.38 156.18 ;
      RECT 18.62 156.06 18.82 156.18 ;
      RECT 19.7 155.04 19.9 155.16 ;
      RECT 18.26 155.04 18.46 155.16 ;
      RECT 17.18 153.78 17.38 153.9 ;
      RECT 18.62 153.78 18.82 153.9 ;
      RECT 20.06 153.78 20.26 153.9 ;
      RECT 19.34 153.54 19.54 153.66 ;
      RECT 17.9 153.54 18.1 153.66 ;
      RECT 19.7 152.52 19.9 152.64 ;
      RECT 18.26 152.28 18.46 152.4 ;
      RECT 17.18 148.74 17.38 148.86 ;
      RECT 18.62 148.74 18.82 148.86 ;
      RECT 20.06 148.74 20.26 148.86 ;
      RECT 19.34 148.5 19.54 148.62 ;
      RECT 17.9 148.5 18.1 148.62 ;
      RECT 17.18 145.98 17.38 146.1 ;
      RECT 17.9 145.98 18.1 146.1 ;
      RECT 18.62 145.98 18.82 146.1 ;
      RECT 19.34 145.98 19.54 146.1 ;
      RECT 20.06 145.98 20.26 146.1 ;
      RECT 18.26 144.96 18.46 145.08 ;
      RECT 19.7 144.72 19.9 144.84 ;
      RECT 20.06 143.46 20.26 143.58 ;
      RECT 17.9 143.46 18.1 143.58 ;
      RECT 19.34 143.7 19.54 143.82 ;
      RECT 18.62 143.7 18.82 143.82 ;
      RECT 17.18 143.7 17.38 143.82 ;
      RECT 18.26 142.44 18.46 142.56 ;
      RECT 19.7 142.2 19.9 142.32 ;
      RECT 19.34 141.18 19.54 141.3 ;
      RECT 17.9 141.18 18.1 141.3 ;
      RECT 17.18 141.18 17.38 141.3 ;
      RECT 18.62 140.94 18.82 141.06 ;
      RECT 20.06 140.94 20.26 141.06 ;
      RECT 19.7 139.92 19.9 140.04 ;
      RECT 18.26 139.68 18.46 139.8 ;
      RECT 17.18 139.138 17.38 139.258 ;
      RECT 17.9 139.138 18.1 139.258 ;
      RECT 18.62 139.138 18.82 139.258 ;
      RECT 19.34 139.138 19.54 139.258 ;
      RECT 20.06 139.138 20.26 139.258 ;
      RECT 17.9 138.66 18.1 138.78 ;
      RECT 18.62 138.66 18.82 138.78 ;
      RECT 20.06 138.66 20.26 138.78 ;
      RECT 19.34 138.42 19.54 138.54 ;
      RECT 17.18 138.42 17.38 138.54 ;
      RECT 19.7 137.4 19.9 137.52 ;
      RECT 18.26 137.16 18.46 137.28 ;
      RECT 17.18 136.618 17.38 136.738 ;
      RECT 17.9 136.618 18.1 136.738 ;
      RECT 18.62 136.618 18.82 136.738 ;
      RECT 19.34 136.618 19.54 136.738 ;
      RECT 20.06 136.618 20.26 136.738 ;
      RECT 19.34 136.14 19.54 136.26 ;
      RECT 17.9 136.14 18.1 136.26 ;
      RECT 17.18 136.14 17.38 136.26 ;
      RECT 20.06 135.9 20.26 136.02 ;
      RECT 18.62 135.9 18.82 136.02 ;
      RECT 19.7 134.88 19.9 135 ;
      RECT 18.26 134.64 18.46 134.76 ;
      RECT 17.18 134.098 17.38 134.218 ;
      RECT 17.9 134.098 18.1 134.218 ;
      RECT 18.62 134.098 18.82 134.218 ;
      RECT 19.34 134.098 19.54 134.218 ;
      RECT 20.06 134.098 20.26 134.218 ;
      RECT 17.18 133.62 17.38 133.74 ;
      RECT 17.9 133.62 18.1 133.74 ;
      RECT 18.62 133.62 18.82 133.74 ;
      RECT 20.06 133.62 20.26 133.74 ;
      RECT 19.34 133.38 19.54 133.5 ;
      RECT 18.26 132.36 18.46 132.48 ;
      RECT 19.7 132.12 19.9 132.24 ;
      RECT 17.18 131.578 17.38 131.698 ;
      RECT 17.9 131.578 18.1 131.698 ;
      RECT 18.62 131.578 18.82 131.698 ;
      RECT 20.06 198.9 20.26 199.02 ;
      RECT 17.54 198.422 17.74 198.542 ;
      RECT 20.42 198.422 20.62 198.542 ;
      RECT 18.98 198.182 19.18 198.302 ;
      RECT 19.7 197.88 19.9 198 ;
      RECT 18.26 197.64 18.46 197.76 ;
      RECT 19.34 196.62 19.54 196.74 ;
      RECT 17.9 196.62 18.1 196.74 ;
      RECT 17.18 196.62 17.38 196.74 ;
      RECT 18.62 196.38 18.82 196.5 ;
      RECT 20.06 196.38 20.26 196.5 ;
      RECT 20.42 195.902 20.62 196.022 ;
      RECT 17.54 195.902 17.74 196.022 ;
      RECT 18.98 195.662 19.18 195.782 ;
      RECT 19.7 195.36 19.9 195.48 ;
      RECT 18.26 195.12 18.46 195.24 ;
      RECT 20.06 193.86 20.26 193.98 ;
      RECT 18.62 193.86 18.82 193.98 ;
      RECT 17.18 194.1 17.38 194.22 ;
      RECT 17.9 194.1 18.1 194.22 ;
      RECT 19.34 194.1 19.54 194.22 ;
      RECT 18.98 194.402 19.18 194.522 ;
      RECT 17.54 194.642 17.74 194.762 ;
      RECT 20.42 194.642 20.62 194.762 ;
      RECT 18.26 192.84 18.46 192.96 ;
      RECT 19.7 192.84 19.9 192.96 ;
      RECT 20.42 193.142 20.62 193.262 ;
      RECT 18.98 193.382 19.18 193.502 ;
      RECT 17.54 193.382 17.74 193.502 ;
      RECT 18.62 191.34 18.82 191.46 ;
      RECT 17.18 191.34 17.38 191.46 ;
      RECT 17.9 191.58 18.1 191.7 ;
      RECT 19.34 191.58 19.54 191.7 ;
      RECT 20.06 191.58 20.26 191.7 ;
      RECT 18.98 191.882 19.18 192.002 ;
      RECT 20.42 192.122 20.62 192.242 ;
      RECT 17.54 192.122 17.74 192.242 ;
      RECT 19.7 190.08 19.9 190.2 ;
      RECT 18.26 190.32 18.46 190.44 ;
      RECT 17.54 190.622 17.74 190.742 ;
      RECT 20.42 190.862 20.62 190.982 ;
      RECT 18.98 190.862 19.18 190.982 ;
      RECT 18.62 188.82 18.82 188.94 ;
      RECT 17.18 189.06 17.38 189.18 ;
      RECT 20.06 189.06 20.26 189.18 ;
      RECT 19.34 189.06 19.54 189.18 ;
      RECT 17.9 189.06 18.1 189.18 ;
      RECT 19.7 187.56 19.9 187.68 ;
      RECT 18.26 187.8 18.46 187.92 ;
      RECT 20.06 186.3 20.26 186.42 ;
      RECT 17.9 186.3 18.1 186.42 ;
      RECT 17.18 186.54 17.38 186.66 ;
      RECT 18.62 186.54 18.82 186.66 ;
      RECT 19.34 186.54 19.54 186.66 ;
      RECT 19.7 185.04 19.9 185.16 ;
      RECT 17.18 183.78 17.38 183.9 ;
      RECT 18.62 183.78 18.82 183.9 ;
      RECT 17.9 184.02 18.1 184.14 ;
      RECT 19.34 184.02 19.54 184.14 ;
      RECT 20.06 184.02 20.26 184.14 ;
      RECT 19.7 182.52 19.9 182.64 ;
      RECT 19.7 180.24 19.9 180.36 ;
      RECT 17.9 181.26 18.1 181.38 ;
      RECT 19.34 181.26 19.54 181.38 ;
      RECT 20.06 181.5 20.26 181.62 ;
      RECT 18.62 181.5 18.82 181.62 ;
      RECT 17.18 181.5 17.38 181.62 ;
      RECT 20.06 178.98 20.26 179.1 ;
      RECT 18.62 178.98 18.82 179.1 ;
      RECT 17.9 178.98 18.1 179.1 ;
      RECT 19.7 177.48 19.9 177.6 ;
      RECT 17.18 178.74 17.38 178.86 ;
      RECT 19.34 178.74 19.54 178.86 ;
      RECT 17.18 176.22 17.38 176.34 ;
      RECT 19.34 176.22 19.54 176.34 ;
      RECT 17.9 176.46 18.1 176.58 ;
      RECT 18.62 176.46 18.82 176.58 ;
      RECT 20.06 176.46 20.26 176.58 ;
      RECT 19.7 174.96 19.9 175.08 ;
      RECT 17.9 173.7 18.1 173.82 ;
      RECT 20.06 173.7 20.26 173.82 ;
      RECT 19.34 173.94 19.54 174.06 ;
      RECT 17.18 173.94 17.38 174.06 ;
      RECT 18.62 173.94 18.82 174.06 ;
      RECT 19.7 172.44 19.9 172.56 ;
      RECT 17.18 171.42 17.38 171.54 ;
      RECT 17.9 171.42 18.1 171.54 ;
      RECT 18.62 171.42 18.82 171.54 ;
      RECT 19.34 171.42 19.54 171.54 ;
      RECT 20.06 171.42 20.26 171.54 ;
      RECT 19.7 169.92 19.9 170.04 ;
      RECT 19.34 168.9 19.54 169.02 ;
      RECT 18.62 168.9 18.82 169.02 ;
      RECT 17.18 168.9 17.38 169.02 ;
      RECT 17.9 168.66 18.1 168.78 ;
      RECT 20.06 168.66 20.26 168.78 ;
      RECT 19.7 167.64 19.9 167.76 ;
      RECT 20.06 166.38 20.26 166.5 ;
      RECT 18.62 166.38 18.82 166.5 ;
      RECT 17.9 166.38 18.1 166.5 ;
      RECT 17.18 166.38 17.38 166.5 ;
      RECT 19.34 166.14 19.54 166.26 ;
      RECT 18.98 218.91 19.18 219.03 ;
      RECT 20.42 218.91 20.62 219.03 ;
      RECT 17.18 218.28 17.38 218.4 ;
      RECT 17.9 218.28 18.1 218.4 ;
      RECT 20.06 218.28 20.26 218.4 ;
      RECT 19.34 218.28 19.54 218.4 ;
      RECT 18.62 218.28 18.82 218.4 ;
      RECT 17.54 217.65 17.74 217.77 ;
      RECT 18.98 217.65 19.18 217.77 ;
      RECT 20.42 217.65 20.62 217.77 ;
      RECT 18.62 217.02 18.82 217.14 ;
      RECT 19.34 217.02 19.54 217.14 ;
      RECT 20.06 217.02 20.26 217.14 ;
      RECT 17.9 217.02 18.1 217.14 ;
      RECT 17.18 217.02 17.38 217.14 ;
      RECT 20.42 216.39 20.62 216.51 ;
      RECT 18.98 216.39 19.18 216.51 ;
      RECT 17.54 216.39 17.74 216.51 ;
      RECT 17.18 215.76 17.38 215.88 ;
      RECT 17.9 215.76 18.1 215.88 ;
      RECT 18.62 215.76 18.82 215.88 ;
      RECT 19.34 215.76 19.54 215.88 ;
      RECT 20.06 215.76 20.26 215.88 ;
      RECT 17.54 215.13 17.74 215.25 ;
      RECT 18.98 215.13 19.18 215.25 ;
      RECT 20.42 215.13 20.62 215.25 ;
      RECT 20.06 214.5 20.26 214.62 ;
      RECT 19.34 214.5 19.54 214.62 ;
      RECT 18.62 214.5 18.82 214.62 ;
      RECT 17.9 214.5 18.1 214.62 ;
      RECT 17.18 214.5 17.38 214.62 ;
      RECT 17.54 213.87 17.74 213.99 ;
      RECT 18.98 213.87 19.18 213.99 ;
      RECT 20.42 213.87 20.62 213.99 ;
      RECT 17.18 213.24 17.38 213.36 ;
      RECT 17.9 213.24 18.1 213.36 ;
      RECT 18.62 213.24 18.82 213.36 ;
      RECT 19.34 213.24 19.54 213.36 ;
      RECT 20.06 213.24 20.26 213.36 ;
      RECT 17.54 212.61 17.74 212.73 ;
      RECT 18.98 212.61 19.18 212.73 ;
      RECT 20.42 212.61 20.62 212.73 ;
      RECT 20.06 211.98 20.26 212.1 ;
      RECT 19.34 211.98 19.54 212.1 ;
      RECT 18.62 211.98 18.82 212.1 ;
      RECT 17.9 211.98 18.1 212.1 ;
      RECT 17.18 211.98 17.38 212.1 ;
      RECT 17.54 211.35 17.74 211.47 ;
      RECT 18.98 211.35 19.18 211.47 ;
      RECT 20.42 211.35 20.62 211.47 ;
      RECT 17.18 210.72 17.38 210.84 ;
      RECT 17.9 210.72 18.1 210.84 ;
      RECT 18.62 210.72 18.82 210.84 ;
      RECT 19.34 210.72 19.54 210.84 ;
      RECT 20.06 210.72 20.26 210.84 ;
      RECT 20.42 210.09 20.62 210.21 ;
      RECT 18.98 210.09 19.18 210.21 ;
      RECT 17.54 210.09 17.74 210.21 ;
      RECT 20.06 209.46 20.26 209.58 ;
      RECT 19.34 209.46 19.54 209.58 ;
      RECT 18.62 209.46 18.82 209.58 ;
      RECT 17.9 209.46 18.1 209.58 ;
      RECT 17.18 209.46 17.38 209.58 ;
      RECT 17.54 208.502 17.74 208.622 ;
      RECT 20.42 208.502 20.62 208.622 ;
      RECT 18.98 208.262 19.18 208.382 ;
      RECT 19.7 207.96 19.9 208.08 ;
      RECT 18.26 207.72 18.46 207.84 ;
      RECT 20.06 206.7 20.26 206.82 ;
      RECT 18.62 206.7 18.82 206.82 ;
      RECT 17.18 206.7 17.38 206.82 ;
      RECT 19.34 206.46 19.54 206.58 ;
      RECT 17.9 206.46 18.1 206.58 ;
      RECT 17.54 205.982 17.74 206.102 ;
      RECT 20.42 205.982 20.62 206.102 ;
      RECT 18.98 205.742 19.18 205.862 ;
      RECT 19.7 205.44 19.9 205.56 ;
      RECT 18.26 205.2 18.46 205.32 ;
      RECT 17.18 204.18 17.38 204.3 ;
      RECT 18.62 204.18 18.82 204.3 ;
      RECT 20.06 204.18 20.26 204.3 ;
      RECT 19.34 203.94 19.54 204.06 ;
      RECT 17.9 203.94 18.1 204.06 ;
      RECT 20.42 203.462 20.62 203.582 ;
      RECT 17.54 203.462 17.74 203.582 ;
      RECT 18.98 203.222 19.18 203.342 ;
      RECT 19.7 202.92 19.9 203.04 ;
      RECT 18.26 202.68 18.46 202.8 ;
      RECT 20.06 201.66 20.26 201.78 ;
      RECT 18.62 201.66 18.82 201.78 ;
      RECT 17.9 201.66 18.1 201.78 ;
      RECT 17.18 201.66 17.38 201.78 ;
      RECT 19.34 201.42 19.54 201.54 ;
      RECT 20.42 200.942 20.62 201.062 ;
      RECT 17.54 200.942 17.74 201.062 ;
      RECT 18.98 200.702 19.18 200.822 ;
      RECT 19.7 200.4 19.9 200.52 ;
      RECT 18.26 200.16 18.46 200.28 ;
      RECT 17.18 199.14 17.38 199.26 ;
      RECT 17.9 199.14 18.1 199.26 ;
      RECT 18.62 199.14 18.82 199.26 ;
      RECT 19.34 199.14 19.54 199.26 ;
      RECT 20.06 234.66 20.26 234.78 ;
      RECT 19.34 234.66 19.54 234.78 ;
      RECT 18.62 234.66 18.82 234.78 ;
      RECT 17.9 234.66 18.1 234.78 ;
      RECT 17.18 234.66 17.38 234.78 ;
      RECT 17.54 234.03 17.74 234.15 ;
      RECT 18.98 234.03 19.18 234.15 ;
      RECT 20.42 234.03 20.62 234.15 ;
      RECT 20.06 233.4 20.26 233.52 ;
      RECT 19.34 233.4 19.54 233.52 ;
      RECT 18.62 233.4 18.82 233.52 ;
      RECT 17.9 233.4 18.1 233.52 ;
      RECT 17.18 233.4 17.38 233.52 ;
      RECT 20.42 232.77 20.62 232.89 ;
      RECT 18.98 232.77 19.18 232.89 ;
      RECT 17.54 232.77 17.74 232.89 ;
      RECT 20.06 232.14 20.26 232.26 ;
      RECT 19.34 232.14 19.54 232.26 ;
      RECT 18.62 232.14 18.82 232.26 ;
      RECT 17.9 232.14 18.1 232.26 ;
      RECT 17.18 232.14 17.38 232.26 ;
      RECT 20.42 231.51 20.62 231.63 ;
      RECT 18.98 231.51 19.18 231.63 ;
      RECT 17.54 231.51 17.74 231.63 ;
      RECT 20.06 230.88 20.26 231 ;
      RECT 19.34 230.88 19.54 231 ;
      RECT 18.62 230.88 18.82 231 ;
      RECT 17.9 230.88 18.1 231 ;
      RECT 17.18 230.88 17.38 231 ;
      RECT 20.42 230.25 20.62 230.37 ;
      RECT 18.98 230.25 19.18 230.37 ;
      RECT 17.54 230.25 17.74 230.37 ;
      RECT 20.06 229.62 20.26 229.74 ;
      RECT 19.34 229.62 19.54 229.74 ;
      RECT 18.62 229.62 18.82 229.74 ;
      RECT 17.9 229.62 18.1 229.74 ;
      RECT 17.18 229.62 17.38 229.74 ;
      RECT 17.54 228.99 17.74 229.11 ;
      RECT 18.98 228.99 19.18 229.11 ;
      RECT 20.42 228.99 20.62 229.11 ;
      RECT 17.18 228.36 17.38 228.48 ;
      RECT 17.9 228.36 18.1 228.48 ;
      RECT 18.62 228.36 18.82 228.48 ;
      RECT 19.34 228.36 19.54 228.48 ;
      RECT 20.06 228.36 20.26 228.48 ;
      RECT 17.54 227.73 17.74 227.85 ;
      RECT 18.98 227.73 19.18 227.85 ;
      RECT 20.42 227.73 20.62 227.85 ;
      RECT 17.18 227.1 17.38 227.22 ;
      RECT 17.9 227.1 18.1 227.22 ;
      RECT 18.62 227.1 18.82 227.22 ;
      RECT 19.34 227.1 19.54 227.22 ;
      RECT 20.06 227.1 20.26 227.22 ;
      RECT 17.54 226.47 17.74 226.59 ;
      RECT 18.98 226.47 19.18 226.59 ;
      RECT 20.42 226.47 20.62 226.59 ;
      RECT 17.18 225.84 17.38 225.96 ;
      RECT 17.9 225.84 18.1 225.96 ;
      RECT 18.62 225.84 18.82 225.96 ;
      RECT 19.34 225.84 19.54 225.96 ;
      RECT 20.06 225.84 20.26 225.96 ;
      RECT 17.54 225.21 17.74 225.33 ;
      RECT 18.98 225.21 19.18 225.33 ;
      RECT 20.42 225.21 20.62 225.33 ;
      RECT 17.18 224.58 17.38 224.7 ;
      RECT 17.9 224.58 18.1 224.7 ;
      RECT 18.62 224.58 18.82 224.7 ;
      RECT 19.34 224.58 19.54 224.7 ;
      RECT 20.06 224.58 20.26 224.7 ;
      RECT 17.54 223.95 17.74 224.07 ;
      RECT 18.98 223.95 19.18 224.07 ;
      RECT 20.42 223.95 20.62 224.07 ;
      RECT 17.18 223.32 17.38 223.44 ;
      RECT 17.9 223.32 18.1 223.44 ;
      RECT 18.62 223.32 18.82 223.44 ;
      RECT 19.34 223.32 19.54 223.44 ;
      RECT 20.06 223.32 20.26 223.44 ;
      RECT 17.54 222.69 17.74 222.81 ;
      RECT 18.98 222.69 19.18 222.81 ;
      RECT 20.42 222.69 20.62 222.81 ;
      RECT 17.18 222.06 17.38 222.18 ;
      RECT 17.9 222.06 18.1 222.18 ;
      RECT 18.62 222.06 18.82 222.18 ;
      RECT 19.34 222.06 19.54 222.18 ;
      RECT 20.06 222.06 20.26 222.18 ;
      RECT 17.54 221.43 17.74 221.55 ;
      RECT 18.98 221.43 19.18 221.55 ;
      RECT 20.42 221.43 20.62 221.55 ;
      RECT 17.18 220.8 17.38 220.92 ;
      RECT 17.9 220.8 18.1 220.92 ;
      RECT 18.62 220.8 18.82 220.92 ;
      RECT 19.34 220.8 19.54 220.92 ;
      RECT 20.06 220.8 20.26 220.92 ;
      RECT 20.42 220.17 20.62 220.29 ;
      RECT 18.98 220.17 19.18 220.29 ;
      RECT 17.54 220.17 17.74 220.29 ;
      RECT 20.06 219.54 20.26 219.66 ;
      RECT 19.34 219.54 19.54 219.66 ;
      RECT 18.62 219.54 18.82 219.66 ;
      RECT 17.9 219.54 18.1 219.66 ;
      RECT 17.18 219.54 17.38 219.66 ;
      RECT 17.54 218.91 17.74 219.03 ;
      RECT 18.62 251.04 18.82 251.16 ;
      RECT 17.9 251.04 18.1 251.16 ;
      RECT 17.18 251.04 17.38 251.16 ;
      RECT 20.42 250.41 20.62 250.53 ;
      RECT 18.98 250.41 19.18 250.53 ;
      RECT 17.54 250.41 17.74 250.53 ;
      RECT 17.18 249.78 17.38 249.9 ;
      RECT 17.9 249.78 18.1 249.9 ;
      RECT 18.62 249.78 18.82 249.9 ;
      RECT 20.06 249.78 20.26 249.9 ;
      RECT 19.34 249.78 19.54 249.9 ;
      RECT 20.42 249.15 20.62 249.27 ;
      RECT 18.98 249.15 19.18 249.27 ;
      RECT 17.54 249.15 17.74 249.27 ;
      RECT 20.06 248.52 20.26 248.64 ;
      RECT 19.34 248.52 19.54 248.64 ;
      RECT 18.62 248.52 18.82 248.64 ;
      RECT 17.9 248.52 18.1 248.64 ;
      RECT 17.18 248.52 17.38 248.64 ;
      RECT 20.42 247.89 20.62 248.01 ;
      RECT 18.98 247.89 19.18 248.01 ;
      RECT 17.54 247.89 17.74 248.01 ;
      RECT 20.06 247.26 20.26 247.38 ;
      RECT 19.34 247.26 19.54 247.38 ;
      RECT 18.62 247.26 18.82 247.38 ;
      RECT 17.9 247.26 18.1 247.38 ;
      RECT 17.18 247.26 17.38 247.38 ;
      RECT 17.18 246 17.38 246.12 ;
      RECT 17.9 246 18.1 246.12 ;
      RECT 20.06 246 20.26 246.12 ;
      RECT 18.62 246 18.82 246.12 ;
      RECT 19.34 246 19.54 246.12 ;
      RECT 17.54 246.63 17.74 246.75 ;
      RECT 18.98 246.63 19.18 246.75 ;
      RECT 20.42 246.63 20.62 246.75 ;
      RECT 17.54 245.37 17.74 245.49 ;
      RECT 18.98 245.37 19.18 245.49 ;
      RECT 20.42 245.37 20.62 245.49 ;
      RECT 18.62 244.74 18.82 244.86 ;
      RECT 17.9 244.74 18.1 244.86 ;
      RECT 17.18 244.74 17.38 244.86 ;
      RECT 20.06 244.74 20.26 244.86 ;
      RECT 19.34 244.74 19.54 244.86 ;
      RECT 20.42 244.11 20.62 244.23 ;
      RECT 18.98 244.11 19.18 244.23 ;
      RECT 17.54 244.11 17.74 244.23 ;
      RECT 20.06 243.48 20.26 243.6 ;
      RECT 19.34 243.48 19.54 243.6 ;
      RECT 18.62 243.48 18.82 243.6 ;
      RECT 17.9 243.48 18.1 243.6 ;
      RECT 17.18 243.48 17.38 243.6 ;
      RECT 20.42 242.85 20.62 242.97 ;
      RECT 18.98 242.85 19.18 242.97 ;
      RECT 17.54 242.85 17.74 242.97 ;
      RECT 19.34 242.22 19.54 242.34 ;
      RECT 20.06 242.22 20.26 242.34 ;
      RECT 18.62 242.22 18.82 242.34 ;
      RECT 17.9 242.22 18.1 242.34 ;
      RECT 17.18 242.22 17.38 242.34 ;
      RECT 20.42 241.59 20.62 241.71 ;
      RECT 17.54 241.59 17.74 241.71 ;
      RECT 18.98 241.59 19.18 241.71 ;
      RECT 20.06 240.96 20.26 241.08 ;
      RECT 19.34 240.96 19.54 241.08 ;
      RECT 18.62 240.96 18.82 241.08 ;
      RECT 17.9 240.96 18.1 241.08 ;
      RECT 17.18 240.96 17.38 241.08 ;
      RECT 20.42 240.33 20.62 240.45 ;
      RECT 18.98 240.33 19.18 240.45 ;
      RECT 17.54 240.33 17.74 240.45 ;
      RECT 20.06 239.7 20.26 239.82 ;
      RECT 19.34 239.7 19.54 239.82 ;
      RECT 18.62 239.7 18.82 239.82 ;
      RECT 17.9 239.7 18.1 239.82 ;
      RECT 17.18 239.7 17.38 239.82 ;
      RECT 20.42 239.07 20.62 239.19 ;
      RECT 18.98 239.07 19.18 239.19 ;
      RECT 17.54 239.07 17.74 239.19 ;
      RECT 17.18 238.44 17.38 238.56 ;
      RECT 17.9 238.44 18.1 238.56 ;
      RECT 18.62 238.44 18.82 238.56 ;
      RECT 19.34 238.44 19.54 238.56 ;
      RECT 20.06 238.44 20.26 238.56 ;
      RECT 17.54 237.81 17.74 237.93 ;
      RECT 18.98 237.81 19.18 237.93 ;
      RECT 20.42 237.81 20.62 237.93 ;
      RECT 17.18 237.18 17.38 237.3 ;
      RECT 17.9 237.18 18.1 237.3 ;
      RECT 18.62 237.18 18.82 237.3 ;
      RECT 19.34 237.18 19.54 237.3 ;
      RECT 20.06 237.18 20.26 237.3 ;
      RECT 20.42 236.55 20.62 236.67 ;
      RECT 18.98 236.55 19.18 236.67 ;
      RECT 17.54 236.55 17.74 236.67 ;
      RECT 20.06 235.92 20.26 236.04 ;
      RECT 19.34 235.92 19.54 236.04 ;
      RECT 18.62 235.92 18.82 236.04 ;
      RECT 17.9 235.92 18.1 236.04 ;
      RECT 17.18 235.92 17.38 236.04 ;
      RECT 20.42 235.29 20.62 235.41 ;
      RECT 18.98 235.29 19.18 235.41 ;
      RECT 17.54 235.29 17.74 235.41 ;
      RECT 17.18 267.42 17.38 267.54 ;
      RECT 20.42 266.79 20.62 266.91 ;
      RECT 18.98 266.79 19.18 266.91 ;
      RECT 17.54 266.79 17.74 266.91 ;
      RECT 20.06 266.16 20.26 266.28 ;
      RECT 19.34 266.16 19.54 266.28 ;
      RECT 18.62 266.16 18.82 266.28 ;
      RECT 17.9 266.16 18.1 266.28 ;
      RECT 17.18 266.16 17.38 266.28 ;
      RECT 20.42 265.53 20.62 265.65 ;
      RECT 18.98 265.53 19.18 265.65 ;
      RECT 17.54 265.53 17.74 265.65 ;
      RECT 20.06 264.9 20.26 265.02 ;
      RECT 19.34 264.9 19.54 265.02 ;
      RECT 18.62 264.9 18.82 265.02 ;
      RECT 17.9 264.9 18.1 265.02 ;
      RECT 17.18 264.9 17.38 265.02 ;
      RECT 20.42 264.27 20.62 264.39 ;
      RECT 18.98 264.27 19.18 264.39 ;
      RECT 17.54 264.27 17.74 264.39 ;
      RECT 20.06 263.64 20.26 263.76 ;
      RECT 19.34 263.64 19.54 263.76 ;
      RECT 18.62 263.64 18.82 263.76 ;
      RECT 17.9 263.64 18.1 263.76 ;
      RECT 17.18 263.64 17.38 263.76 ;
      RECT 20.42 263.01 20.62 263.13 ;
      RECT 18.98 263.01 19.18 263.13 ;
      RECT 17.54 263.01 17.74 263.13 ;
      RECT 20.06 262.38 20.26 262.5 ;
      RECT 19.34 262.38 19.54 262.5 ;
      RECT 18.62 262.38 18.82 262.5 ;
      RECT 17.9 262.38 18.1 262.5 ;
      RECT 17.18 262.38 17.38 262.5 ;
      RECT 20.42 261.75 20.62 261.87 ;
      RECT 18.98 261.75 19.18 261.87 ;
      RECT 17.54 261.75 17.74 261.87 ;
      RECT 17.9 261.12 18.1 261.24 ;
      RECT 20.06 261.12 20.26 261.24 ;
      RECT 18.62 261.12 18.82 261.24 ;
      RECT 19.34 261.12 19.54 261.24 ;
      RECT 17.18 261.12 17.38 261.24 ;
      RECT 20.42 260.49 20.62 260.61 ;
      RECT 18.98 260.49 19.18 260.61 ;
      RECT 17.54 260.49 17.74 260.61 ;
      RECT 20.06 259.86 20.26 259.98 ;
      RECT 19.34 259.86 19.54 259.98 ;
      RECT 18.62 259.86 18.82 259.98 ;
      RECT 17.9 259.86 18.1 259.98 ;
      RECT 17.18 259.86 17.38 259.98 ;
      RECT 20.42 259.23 20.62 259.35 ;
      RECT 18.98 259.23 19.18 259.35 ;
      RECT 17.54 259.23 17.74 259.35 ;
      RECT 20.06 258.6 20.26 258.72 ;
      RECT 19.34 258.6 19.54 258.72 ;
      RECT 18.62 258.6 18.82 258.72 ;
      RECT 17.9 258.6 18.1 258.72 ;
      RECT 17.18 258.6 17.38 258.72 ;
      RECT 20.42 257.97 20.62 258.09 ;
      RECT 18.98 257.97 19.18 258.09 ;
      RECT 17.54 257.97 17.74 258.09 ;
      RECT 20.06 257.34 20.26 257.46 ;
      RECT 19.34 257.34 19.54 257.46 ;
      RECT 18.62 257.34 18.82 257.46 ;
      RECT 17.9 257.34 18.1 257.46 ;
      RECT 17.18 257.34 17.38 257.46 ;
      RECT 20.42 256.71 20.62 256.83 ;
      RECT 18.98 256.71 19.18 256.83 ;
      RECT 17.54 256.71 17.74 256.83 ;
      RECT 20.06 256.08 20.26 256.2 ;
      RECT 19.34 256.08 19.54 256.2 ;
      RECT 18.62 256.08 18.82 256.2 ;
      RECT 17.9 256.08 18.1 256.2 ;
      RECT 17.18 256.08 17.38 256.2 ;
      RECT 20.42 255.45 20.62 255.57 ;
      RECT 18.98 255.45 19.18 255.57 ;
      RECT 17.54 255.45 17.74 255.57 ;
      RECT 20.06 254.82 20.26 254.94 ;
      RECT 19.34 254.82 19.54 254.94 ;
      RECT 18.62 254.82 18.82 254.94 ;
      RECT 17.9 254.82 18.1 254.94 ;
      RECT 17.18 254.82 17.38 254.94 ;
      RECT 20.42 254.19 20.62 254.31 ;
      RECT 18.98 254.19 19.18 254.31 ;
      RECT 17.54 254.19 17.74 254.31 ;
      RECT 20.06 253.56 20.26 253.68 ;
      RECT 19.34 253.56 19.54 253.68 ;
      RECT 18.62 253.56 18.82 253.68 ;
      RECT 17.9 253.56 18.1 253.68 ;
      RECT 17.18 253.56 17.38 253.68 ;
      RECT 20.42 252.93 20.62 253.05 ;
      RECT 18.98 252.93 19.18 253.05 ;
      RECT 17.54 252.93 17.74 253.05 ;
      RECT 20.06 252.3 20.26 252.42 ;
      RECT 19.34 252.3 19.54 252.42 ;
      RECT 18.62 252.3 18.82 252.42 ;
      RECT 17.9 252.3 18.1 252.42 ;
      RECT 17.18 252.3 17.38 252.42 ;
      RECT 20.42 251.67 20.62 251.79 ;
      RECT 18.98 251.67 19.18 251.79 ;
      RECT 17.54 251.67 17.74 251.79 ;
      RECT 20.06 251.04 20.26 251.16 ;
      RECT 19.34 251.04 19.54 251.16 ;
      RECT 20.78 118.978 20.98 119.098 ;
      RECT 24.38 118.5 24.58 118.62 ;
      RECT 22.94 118.5 23.14 118.62 ;
      RECT 23.66 118.26 23.86 118.38 ;
      RECT 20.78 118.26 20.98 118.38 ;
      RECT 19.7 348.339 19.9 348.459 ;
      RECT 18.26 348.339 18.46 348.459 ;
      RECT 20.06 325.9425 20.26 326.0625 ;
      RECT 19.34 325.9425 19.54 326.0625 ;
      RECT 18.62 325.9425 18.82 326.0625 ;
      RECT 17.9 325.9425 18.1 326.0625 ;
      RECT 17.18 325.9425 17.38 326.0625 ;
      RECT 19.7 323.3835 19.9 323.5035 ;
      RECT 18.26 323.3835 18.46 323.5035 ;
      RECT 17.18 305.967 17.38 306.087 ;
      RECT 20.06 305.967 20.26 306.087 ;
      RECT 17.9 305.967 18.1 306.087 ;
      RECT 18.62 305.967 18.82 306.087 ;
      RECT 19.34 305.967 19.54 306.087 ;
      RECT 19.7 305.498 19.9 305.618 ;
      RECT 18.26 305.498 18.46 305.618 ;
      RECT 20.06 283.087 20.26 283.207 ;
      RECT 19.34 283.087 19.54 283.207 ;
      RECT 18.62 283.087 18.82 283.207 ;
      RECT 17.9 283.087 18.1 283.207 ;
      RECT 17.18 283.087 17.38 283.207 ;
      RECT 17.9 278.76 18.1 278.88 ;
      RECT 18.62 278.76 18.82 278.88 ;
      RECT 17.18 278.76 17.38 278.88 ;
      RECT 20.06 278.76 20.26 278.88 ;
      RECT 19.34 278.76 19.54 278.88 ;
      RECT 20.42 278.13 20.62 278.25 ;
      RECT 18.98 278.13 19.18 278.25 ;
      RECT 17.54 278.13 17.74 278.25 ;
      RECT 20.06 277.5 20.26 277.62 ;
      RECT 19.34 277.5 19.54 277.62 ;
      RECT 18.62 277.5 18.82 277.62 ;
      RECT 17.9 277.5 18.1 277.62 ;
      RECT 17.18 277.5 17.38 277.62 ;
      RECT 20.42 276.87 20.62 276.99 ;
      RECT 18.98 276.87 19.18 276.99 ;
      RECT 17.54 276.87 17.74 276.99 ;
      RECT 20.06 276.24 20.26 276.36 ;
      RECT 19.34 276.24 19.54 276.36 ;
      RECT 18.62 276.24 18.82 276.36 ;
      RECT 17.9 276.24 18.1 276.36 ;
      RECT 17.18 276.24 17.38 276.36 ;
      RECT 20.42 275.61 20.62 275.73 ;
      RECT 18.98 275.61 19.18 275.73 ;
      RECT 17.54 275.61 17.74 275.73 ;
      RECT 20.06 274.98 20.26 275.1 ;
      RECT 19.34 274.98 19.54 275.1 ;
      RECT 18.62 274.98 18.82 275.1 ;
      RECT 17.9 274.98 18.1 275.1 ;
      RECT 17.18 274.98 17.38 275.1 ;
      RECT 20.42 274.35 20.62 274.47 ;
      RECT 18.98 274.35 19.18 274.47 ;
      RECT 17.54 274.35 17.74 274.47 ;
      RECT 20.06 273.72 20.26 273.84 ;
      RECT 19.34 273.72 19.54 273.84 ;
      RECT 18.62 273.72 18.82 273.84 ;
      RECT 17.9 273.72 18.1 273.84 ;
      RECT 17.18 273.72 17.38 273.84 ;
      RECT 20.42 273.09 20.62 273.21 ;
      RECT 18.98 273.09 19.18 273.21 ;
      RECT 17.54 273.09 17.74 273.21 ;
      RECT 20.06 272.46 20.26 272.58 ;
      RECT 19.34 272.46 19.54 272.58 ;
      RECT 18.62 272.46 18.82 272.58 ;
      RECT 17.9 272.46 18.1 272.58 ;
      RECT 17.18 272.46 17.38 272.58 ;
      RECT 20.42 271.83 20.62 271.95 ;
      RECT 18.98 271.83 19.18 271.95 ;
      RECT 17.54 271.83 17.74 271.95 ;
      RECT 20.06 271.2 20.26 271.32 ;
      RECT 19.34 271.2 19.54 271.32 ;
      RECT 18.62 271.2 18.82 271.32 ;
      RECT 17.9 271.2 18.1 271.32 ;
      RECT 17.18 271.2 17.38 271.32 ;
      RECT 20.42 270.57 20.62 270.69 ;
      RECT 18.98 270.57 19.18 270.69 ;
      RECT 17.54 270.57 17.74 270.69 ;
      RECT 20.06 269.94 20.26 270.06 ;
      RECT 19.34 269.94 19.54 270.06 ;
      RECT 18.62 269.94 18.82 270.06 ;
      RECT 17.9 269.94 18.1 270.06 ;
      RECT 17.18 269.94 17.38 270.06 ;
      RECT 20.42 269.31 20.62 269.43 ;
      RECT 18.98 269.31 19.18 269.43 ;
      RECT 17.54 269.31 17.74 269.43 ;
      RECT 17.18 268.68 17.38 268.8 ;
      RECT 17.9 268.68 18.1 268.8 ;
      RECT 20.06 268.68 20.26 268.8 ;
      RECT 19.34 268.68 19.54 268.8 ;
      RECT 18.62 268.68 18.82 268.8 ;
      RECT 20.42 268.05 20.62 268.17 ;
      RECT 18.98 268.05 19.18 268.17 ;
      RECT 17.54 268.05 17.74 268.17 ;
      RECT 20.06 267.42 20.26 267.54 ;
      RECT 19.34 267.42 19.54 267.54 ;
      RECT 18.62 267.42 18.82 267.54 ;
      RECT 17.9 267.42 18.1 267.54 ;
      RECT 22.94 156.3 23.14 156.42 ;
      RECT 23.3 156.842 23.5 156.962 ;
      RECT 24.02 155.04 24.22 155.16 ;
      RECT 20.78 153.54 20.98 153.66 ;
      RECT 24.38 153.78 24.58 153.9 ;
      RECT 23.66 153.78 23.86 153.9 ;
      RECT 22.94 153.78 23.14 153.9 ;
      RECT 24.02 152.28 24.22 152.4 ;
      RECT 20.78 148.74 20.98 148.86 ;
      RECT 22.94 148.5 23.14 148.62 ;
      RECT 24.38 148.5 24.58 148.62 ;
      RECT 23.66 148.74 23.86 148.86 ;
      RECT 20.78 145.98 20.98 146.1 ;
      RECT 24.02 144.96 24.22 145.08 ;
      RECT 24.38 145.98 24.58 146.1 ;
      RECT 23.66 145.98 23.86 146.1 ;
      RECT 22.94 145.98 23.14 146.1 ;
      RECT 24.38 143.46 24.58 143.58 ;
      RECT 22.94 143.46 23.14 143.58 ;
      RECT 20.78 143.7 20.98 143.82 ;
      RECT 23.66 143.7 23.86 143.82 ;
      RECT 24.02 142.44 24.22 142.56 ;
      RECT 23.66 141.18 23.86 141.3 ;
      RECT 22.94 140.94 23.14 141.06 ;
      RECT 24.38 140.94 24.58 141.06 ;
      RECT 20.78 141.18 20.98 141.3 ;
      RECT 24.02 139.68 24.22 139.8 ;
      RECT 22.94 139.138 23.14 139.258 ;
      RECT 23.66 139.138 23.86 139.258 ;
      RECT 24.38 139.138 24.58 139.258 ;
      RECT 22.94 138.66 23.14 138.78 ;
      RECT 24.38 138.66 24.58 138.78 ;
      RECT 23.66 138.42 23.86 138.54 ;
      RECT 20.78 139.138 20.98 139.258 ;
      RECT 20.78 138.42 20.98 138.54 ;
      RECT 24.02 137.16 24.22 137.28 ;
      RECT 22.94 136.618 23.14 136.738 ;
      RECT 23.66 136.618 23.86 136.738 ;
      RECT 24.38 136.618 24.58 136.738 ;
      RECT 20.78 136.618 20.98 136.738 ;
      RECT 24.38 136.14 24.58 136.26 ;
      RECT 23.66 136.14 23.86 136.26 ;
      RECT 22.94 135.9 23.14 136.02 ;
      RECT 20.78 136.14 20.98 136.26 ;
      RECT 24.02 134.88 24.22 135 ;
      RECT 22.94 134.098 23.14 134.218 ;
      RECT 23.66 134.098 23.86 134.218 ;
      RECT 24.38 134.098 24.58 134.218 ;
      RECT 20.78 134.098 20.98 134.218 ;
      RECT 22.94 133.62 23.14 133.74 ;
      RECT 24.38 133.62 24.58 133.74 ;
      RECT 23.66 133.38 23.86 133.5 ;
      RECT 20.78 133.62 20.98 133.74 ;
      RECT 24.02 132.36 24.22 132.48 ;
      RECT 22.94 131.578 23.14 131.698 ;
      RECT 23.66 131.578 23.86 131.698 ;
      RECT 24.38 131.578 24.58 131.698 ;
      RECT 23.66 131.1 23.86 131.22 ;
      RECT 20.78 131.578 20.98 131.698 ;
      RECT 20.78 131.1 20.98 131.22 ;
      RECT 22.94 130.86 23.14 130.98 ;
      RECT 24.38 130.86 24.58 130.98 ;
      RECT 24.02 129.84 24.22 129.96 ;
      RECT 22.94 129.058 23.14 129.178 ;
      RECT 23.66 129.058 23.86 129.178 ;
      RECT 24.38 129.058 24.58 129.178 ;
      RECT 23.66 128.58 23.86 128.7 ;
      RECT 24.38 128.34 24.58 128.46 ;
      RECT 22.94 128.34 23.14 128.46 ;
      RECT 20.78 129.058 20.98 129.178 ;
      RECT 20.78 128.58 20.98 128.7 ;
      RECT 24.02 127.32 24.22 127.44 ;
      RECT 22.94 126.538 23.14 126.658 ;
      RECT 23.66 126.538 23.86 126.658 ;
      RECT 24.38 126.538 24.58 126.658 ;
      RECT 23.66 126.06 23.86 126.18 ;
      RECT 24.38 126.06 24.58 126.18 ;
      RECT 22.94 125.82 23.14 125.94 ;
      RECT 20.78 126.538 20.98 126.658 ;
      RECT 20.78 126.06 20.98 126.18 ;
      RECT 24.02 124.8 24.22 124.92 ;
      RECT 22.94 124.018 23.14 124.138 ;
      RECT 23.66 124.018 23.86 124.138 ;
      RECT 24.38 124.018 24.58 124.138 ;
      RECT 22.94 123.54 23.14 123.66 ;
      RECT 23.66 123.54 23.86 123.66 ;
      RECT 24.38 123.54 24.58 123.66 ;
      RECT 20.78 124.018 20.98 124.138 ;
      RECT 20.78 123.3 20.98 123.42 ;
      RECT 24.02 122.28 24.22 122.4 ;
      RECT 22.94 121.498 23.14 121.618 ;
      RECT 23.66 121.498 23.86 121.618 ;
      RECT 24.38 121.498 24.58 121.618 ;
      RECT 20.78 121.498 20.98 121.618 ;
      RECT 23.66 121.02 23.86 121.14 ;
      RECT 22.94 120.78 23.14 120.9 ;
      RECT 24.38 120.78 24.58 120.9 ;
      RECT 20.78 121.02 20.98 121.14 ;
      RECT 24.02 119.76 24.22 119.88 ;
      RECT 22.94 118.978 23.14 119.098 ;
      RECT 23.66 118.978 23.86 119.098 ;
      RECT 24.38 118.978 24.58 119.098 ;
      RECT 24.38 204.18 24.58 204.3 ;
      RECT 22.94 204.18 23.14 204.3 ;
      RECT 24.02 202.68 24.22 202.8 ;
      RECT 23.3 203.222 23.5 203.342 ;
      RECT 20.78 201.42 20.98 201.54 ;
      RECT 23.3 200.702 23.5 200.822 ;
      RECT 23.66 201.42 23.86 201.54 ;
      RECT 22.94 201.66 23.14 201.78 ;
      RECT 24.38 201.66 24.58 201.78 ;
      RECT 24.02 200.16 24.22 200.28 ;
      RECT 20.78 199.14 20.98 199.26 ;
      RECT 23.3 198.182 23.5 198.302 ;
      RECT 22.94 198.9 23.14 199.02 ;
      RECT 24.38 199.14 24.58 199.26 ;
      RECT 23.66 199.14 23.86 199.26 ;
      RECT 20.78 196.62 20.98 196.74 ;
      RECT 22.94 196.62 23.14 196.74 ;
      RECT 24.38 196.62 24.58 196.74 ;
      RECT 24.02 197.64 24.22 197.76 ;
      RECT 23.3 195.662 23.5 195.782 ;
      RECT 23.66 196.38 23.86 196.5 ;
      RECT 20.78 194.1 20.98 194.22 ;
      RECT 24.38 193.86 24.58 193.98 ;
      RECT 22.94 194.1 23.14 194.22 ;
      RECT 23.66 194.1 23.86 194.22 ;
      RECT 23.3 194.642 23.5 194.762 ;
      RECT 24.02 195.12 24.22 195.24 ;
      RECT 24.02 192.84 24.22 192.96 ;
      RECT 23.3 193.382 23.5 193.502 ;
      RECT 20.78 191.34 20.98 191.46 ;
      RECT 22.94 191.34 23.14 191.46 ;
      RECT 23.66 191.58 23.86 191.7 ;
      RECT 24.38 191.58 24.58 191.7 ;
      RECT 23.3 192.122 23.5 192.242 ;
      RECT 24.02 190.32 24.22 190.44 ;
      RECT 23.3 190.862 23.5 190.982 ;
      RECT 20.78 188.82 20.98 188.94 ;
      RECT 24.38 188.82 24.58 188.94 ;
      RECT 23.66 189.06 23.86 189.18 ;
      RECT 22.94 189.06 23.14 189.18 ;
      RECT 24.02 187.8 24.22 187.92 ;
      RECT 20.78 186.54 20.98 186.66 ;
      RECT 24.38 186.3 24.58 186.42 ;
      RECT 22.94 186.3 23.14 186.42 ;
      RECT 23.66 186.54 23.86 186.66 ;
      RECT 24.02 185.28 24.22 185.4 ;
      RECT 20.78 183.78 20.98 183.9 ;
      RECT 23.66 183.78 23.86 183.9 ;
      RECT 22.94 184.02 23.14 184.14 ;
      RECT 24.38 184.02 24.58 184.14 ;
      RECT 24.02 182.76 24.22 182.88 ;
      RECT 20.78 181.26 20.98 181.38 ;
      RECT 23.66 181.26 23.86 181.38 ;
      RECT 24.38 181.5 24.58 181.62 ;
      RECT 22.94 181.5 23.14 181.62 ;
      RECT 24.38 178.98 24.58 179.1 ;
      RECT 22.94 178.98 23.14 179.1 ;
      RECT 24.02 180 24.22 180.12 ;
      RECT 20.78 178.74 20.98 178.86 ;
      RECT 24.02 177.72 24.22 177.84 ;
      RECT 23.66 178.74 23.86 178.86 ;
      RECT 20.78 176.46 20.98 176.58 ;
      RECT 22.94 176.22 23.14 176.34 ;
      RECT 23.66 176.46 23.86 176.58 ;
      RECT 24.38 176.46 24.58 176.58 ;
      RECT 24.02 175.2 24.22 175.32 ;
      RECT 20.78 173.94 20.98 174.06 ;
      RECT 22.94 173.7 23.14 173.82 ;
      RECT 24.38 173.7 24.58 173.82 ;
      RECT 23.66 173.94 23.86 174.06 ;
      RECT 24.02 172.68 24.22 172.8 ;
      RECT 20.78 171.42 20.98 171.54 ;
      RECT 23.66 171.18 23.86 171.3 ;
      RECT 22.94 171.42 23.14 171.54 ;
      RECT 24.38 171.42 24.58 171.54 ;
      RECT 24.02 170.16 24.22 170.28 ;
      RECT 20.78 168.9 20.98 169.02 ;
      RECT 22.94 168.66 23.14 168.78 ;
      RECT 23.66 168.9 23.86 169.02 ;
      RECT 24.38 168.9 24.58 169.02 ;
      RECT 24.02 167.4 24.22 167.52 ;
      RECT 20.78 166.38 20.98 166.5 ;
      RECT 24.38 166.14 24.58 166.26 ;
      RECT 22.94 166.38 23.14 166.5 ;
      RECT 23.66 166.38 23.86 166.5 ;
      RECT 20.78 163.86 20.98 163.98 ;
      RECT 23.66 163.86 23.86 163.98 ;
      RECT 24.38 163.86 24.58 163.98 ;
      RECT 24.02 165.12 24.22 165.24 ;
      RECT 24.02 162.6 24.22 162.72 ;
      RECT 22.94 163.62 23.14 163.74 ;
      RECT 24.38 161.1 24.58 161.22 ;
      RECT 24.02 160.08 24.22 160.2 ;
      RECT 20.78 158.82 20.98 158.94 ;
      RECT 22.94 158.58 23.14 158.7 ;
      RECT 24.38 158.58 24.58 158.7 ;
      RECT 23.66 158.82 23.86 158.94 ;
      RECT 24.02 157.32 24.22 157.44 ;
      RECT 23.3 158.038 23.5 158.158 ;
      RECT 20.78 156.06 20.98 156.18 ;
      RECT 23.66 156.06 23.86 156.18 ;
      RECT 24.38 156.3 24.58 156.42 ;
      RECT 23.66 233.4 23.86 233.52 ;
      RECT 22.94 233.4 23.14 233.52 ;
      RECT 20.78 230.88 20.98 231 ;
      RECT 22.94 230.88 23.14 231 ;
      RECT 23.66 230.88 23.86 231 ;
      RECT 24.38 230.88 24.58 231 ;
      RECT 23.3 231.51 23.5 231.63 ;
      RECT 20.78 229.62 20.98 229.74 ;
      RECT 24.38 229.62 24.58 229.74 ;
      RECT 23.66 229.62 23.86 229.74 ;
      RECT 22.94 229.62 23.14 229.74 ;
      RECT 23.3 230.25 23.5 230.37 ;
      RECT 20.78 228.36 20.98 228.48 ;
      RECT 24.38 228.36 24.58 228.48 ;
      RECT 23.66 228.36 23.86 228.48 ;
      RECT 22.94 228.36 23.14 228.48 ;
      RECT 23.3 228.99 23.5 229.11 ;
      RECT 20.78 227.1 20.98 227.22 ;
      RECT 24.38 227.1 24.58 227.22 ;
      RECT 23.66 227.1 23.86 227.22 ;
      RECT 22.94 227.1 23.14 227.22 ;
      RECT 23.3 227.73 23.5 227.85 ;
      RECT 20.78 225.84 20.98 225.96 ;
      RECT 24.38 225.84 24.58 225.96 ;
      RECT 23.66 225.84 23.86 225.96 ;
      RECT 22.94 225.84 23.14 225.96 ;
      RECT 23.3 226.47 23.5 226.59 ;
      RECT 20.78 224.58 20.98 224.7 ;
      RECT 23.3 223.95 23.5 224.07 ;
      RECT 24.38 224.58 24.58 224.7 ;
      RECT 23.66 224.58 23.86 224.7 ;
      RECT 22.94 224.58 23.14 224.7 ;
      RECT 23.3 225.21 23.5 225.33 ;
      RECT 20.78 223.32 20.98 223.44 ;
      RECT 23.3 222.69 23.5 222.81 ;
      RECT 24.38 223.32 24.58 223.44 ;
      RECT 23.66 223.32 23.86 223.44 ;
      RECT 22.94 223.32 23.14 223.44 ;
      RECT 20.78 222.06 20.98 222.18 ;
      RECT 23.3 221.43 23.5 221.55 ;
      RECT 24.38 222.06 24.58 222.18 ;
      RECT 23.66 222.06 23.86 222.18 ;
      RECT 22.94 222.06 23.14 222.18 ;
      RECT 20.78 220.8 20.98 220.92 ;
      RECT 24.38 220.8 24.58 220.92 ;
      RECT 23.66 220.8 23.86 220.92 ;
      RECT 22.94 220.8 23.14 220.92 ;
      RECT 23.3 220.17 23.5 220.29 ;
      RECT 20.78 219.54 20.98 219.66 ;
      RECT 23.3 218.91 23.5 219.03 ;
      RECT 22.94 219.54 23.14 219.66 ;
      RECT 23.66 219.54 23.86 219.66 ;
      RECT 24.38 219.54 24.58 219.66 ;
      RECT 20.78 218.28 20.98 218.4 ;
      RECT 23.3 217.65 23.5 217.77 ;
      RECT 22.94 218.28 23.14 218.4 ;
      RECT 23.66 218.28 23.86 218.4 ;
      RECT 24.38 218.28 24.58 218.4 ;
      RECT 20.78 217.02 20.98 217.14 ;
      RECT 20.78 215.76 20.98 215.88 ;
      RECT 24.38 215.76 24.58 215.88 ;
      RECT 23.66 215.76 23.86 215.88 ;
      RECT 22.94 215.76 23.14 215.88 ;
      RECT 23.3 216.39 23.5 216.51 ;
      RECT 24.38 217.02 24.58 217.14 ;
      RECT 23.66 217.02 23.86 217.14 ;
      RECT 22.94 217.02 23.14 217.14 ;
      RECT 20.78 214.5 20.98 214.62 ;
      RECT 22.94 214.5 23.14 214.62 ;
      RECT 23.66 214.5 23.86 214.62 ;
      RECT 24.38 214.5 24.58 214.62 ;
      RECT 23.3 215.13 23.5 215.25 ;
      RECT 20.78 213.24 20.98 213.36 ;
      RECT 24.38 213.24 24.58 213.36 ;
      RECT 23.66 213.24 23.86 213.36 ;
      RECT 22.94 213.24 23.14 213.36 ;
      RECT 23.3 213.87 23.5 213.99 ;
      RECT 20.78 211.98 20.98 212.1 ;
      RECT 22.94 211.98 23.14 212.1 ;
      RECT 23.66 211.98 23.86 212.1 ;
      RECT 24.38 211.98 24.58 212.1 ;
      RECT 23.3 212.61 23.5 212.73 ;
      RECT 20.78 210.72 20.98 210.84 ;
      RECT 24.38 210.72 24.58 210.84 ;
      RECT 23.66 210.72 23.86 210.84 ;
      RECT 22.94 210.72 23.14 210.84 ;
      RECT 23.3 211.35 23.5 211.47 ;
      RECT 20.78 209.46 20.98 209.58 ;
      RECT 22.94 209.46 23.14 209.58 ;
      RECT 23.66 209.46 23.86 209.58 ;
      RECT 24.38 209.46 24.58 209.58 ;
      RECT 23.3 210.09 23.5 210.21 ;
      RECT 24.02 207.72 24.22 207.84 ;
      RECT 23.3 208.262 23.5 208.382 ;
      RECT 20.78 206.46 20.98 206.58 ;
      RECT 23.66 206.46 23.86 206.58 ;
      RECT 22.94 206.7 23.14 206.82 ;
      RECT 24.38 206.7 24.58 206.82 ;
      RECT 24.02 205.2 24.22 205.32 ;
      RECT 23.3 205.742 23.5 205.862 ;
      RECT 20.78 204.18 20.98 204.3 ;
      RECT 23.66 203.94 23.86 204.06 ;
      RECT 23.3 256.71 23.5 256.83 ;
      RECT 22.94 257.34 23.14 257.46 ;
      RECT 23.66 257.34 23.86 257.46 ;
      RECT 24.38 257.34 24.58 257.46 ;
      RECT 23.3 257.97 23.5 258.09 ;
      RECT 20.78 256.08 20.98 256.2 ;
      RECT 23.3 255.45 23.5 255.57 ;
      RECT 22.94 256.08 23.14 256.2 ;
      RECT 23.66 256.08 23.86 256.2 ;
      RECT 24.38 256.08 24.58 256.2 ;
      RECT 20.78 254.82 20.98 254.94 ;
      RECT 23.3 254.19 23.5 254.31 ;
      RECT 22.94 254.82 23.14 254.94 ;
      RECT 23.66 254.82 23.86 254.94 ;
      RECT 24.38 254.82 24.58 254.94 ;
      RECT 20.78 253.56 20.98 253.68 ;
      RECT 23.3 252.93 23.5 253.05 ;
      RECT 22.94 253.56 23.14 253.68 ;
      RECT 23.66 253.56 23.86 253.68 ;
      RECT 24.38 253.56 24.58 253.68 ;
      RECT 20.78 252.3 20.98 252.42 ;
      RECT 23.3 251.67 23.5 251.79 ;
      RECT 22.94 252.3 23.14 252.42 ;
      RECT 23.66 252.3 23.86 252.42 ;
      RECT 24.38 252.3 24.58 252.42 ;
      RECT 22.94 251.04 23.14 251.16 ;
      RECT 23.3 250.41 23.5 250.53 ;
      RECT 20.78 251.04 20.98 251.16 ;
      RECT 23.66 251.04 23.86 251.16 ;
      RECT 24.38 251.04 24.58 251.16 ;
      RECT 24.38 249.78 24.58 249.9 ;
      RECT 23.66 249.78 23.86 249.9 ;
      RECT 22.94 249.78 23.14 249.9 ;
      RECT 23.3 249.15 23.5 249.27 ;
      RECT 24.38 248.52 24.58 248.64 ;
      RECT 23.66 248.52 23.86 248.64 ;
      RECT 22.94 248.52 23.14 248.64 ;
      RECT 20.78 249.78 20.98 249.9 ;
      RECT 20.78 248.52 20.98 248.64 ;
      RECT 23.3 247.89 23.5 248.01 ;
      RECT 24.38 247.26 24.58 247.38 ;
      RECT 23.66 247.26 23.86 247.38 ;
      RECT 22.94 247.26 23.14 247.38 ;
      RECT 20.78 247.26 20.98 247.38 ;
      RECT 23.3 246.63 23.5 246.75 ;
      RECT 20.78 246 20.98 246.12 ;
      RECT 24.38 246 24.58 246.12 ;
      RECT 23.66 246 23.86 246.12 ;
      RECT 22.94 246 23.14 246.12 ;
      RECT 20.78 244.74 20.98 244.86 ;
      RECT 24.38 244.74 24.58 244.86 ;
      RECT 22.94 244.74 23.14 244.86 ;
      RECT 23.66 244.74 23.86 244.86 ;
      RECT 23.3 245.37 23.5 245.49 ;
      RECT 20.78 243.48 20.98 243.6 ;
      RECT 22.94 243.48 23.14 243.6 ;
      RECT 23.66 243.48 23.86 243.6 ;
      RECT 24.38 243.48 24.58 243.6 ;
      RECT 23.3 244.11 23.5 244.23 ;
      RECT 20.78 242.22 20.98 242.34 ;
      RECT 22.94 242.22 23.14 242.34 ;
      RECT 23.66 242.22 23.86 242.34 ;
      RECT 24.38 242.22 24.58 242.34 ;
      RECT 23.3 242.85 23.5 242.97 ;
      RECT 20.78 240.96 20.98 241.08 ;
      RECT 23.3 240.33 23.5 240.45 ;
      RECT 22.94 240.96 23.14 241.08 ;
      RECT 23.66 240.96 23.86 241.08 ;
      RECT 24.38 240.96 24.58 241.08 ;
      RECT 23.3 241.59 23.5 241.71 ;
      RECT 20.78 239.7 20.98 239.82 ;
      RECT 23.3 239.07 23.5 239.19 ;
      RECT 22.94 239.7 23.14 239.82 ;
      RECT 23.66 239.7 23.86 239.82 ;
      RECT 24.38 239.7 24.58 239.82 ;
      RECT 20.78 238.44 20.98 238.56 ;
      RECT 23.3 237.81 23.5 237.93 ;
      RECT 24.38 238.44 24.58 238.56 ;
      RECT 23.66 238.44 23.86 238.56 ;
      RECT 22.94 238.44 23.14 238.56 ;
      RECT 20.78 237.18 20.98 237.3 ;
      RECT 23.3 236.55 23.5 236.67 ;
      RECT 24.38 237.18 24.58 237.3 ;
      RECT 23.66 237.18 23.86 237.3 ;
      RECT 22.94 237.18 23.14 237.3 ;
      RECT 20.78 235.92 20.98 236.04 ;
      RECT 23.3 235.29 23.5 235.41 ;
      RECT 22.94 235.92 23.14 236.04 ;
      RECT 23.66 235.92 23.86 236.04 ;
      RECT 24.38 235.92 24.58 236.04 ;
      RECT 20.78 234.66 20.98 234.78 ;
      RECT 23.3 234.03 23.5 234.15 ;
      RECT 22.94 234.66 23.14 234.78 ;
      RECT 23.66 234.66 23.86 234.78 ;
      RECT 24.38 234.66 24.58 234.78 ;
      RECT 20.78 233.4 20.98 233.52 ;
      RECT 20.78 232.14 20.98 232.26 ;
      RECT 22.94 232.14 23.14 232.26 ;
      RECT 23.66 232.14 23.86 232.26 ;
      RECT 24.38 232.14 24.58 232.26 ;
      RECT 23.3 232.77 23.5 232.89 ;
      RECT 24.38 233.4 24.58 233.52 ;
      RECT 26.54 118.26 26.74 118.38 ;
      RECT 25.1 118.26 25.3 118.38 ;
      RECT 24.02 348.339 24.22 348.459 ;
      RECT 20.78 325.9425 20.98 326.0625 ;
      RECT 24.38 325.9425 24.58 326.0625 ;
      RECT 23.66 325.9425 23.86 326.0625 ;
      RECT 22.94 325.9425 23.14 326.0625 ;
      RECT 24.02 323.3835 24.22 323.5035 ;
      RECT 20.78 305.967 20.98 306.087 ;
      RECT 24.38 305.967 24.58 306.087 ;
      RECT 23.66 305.967 23.86 306.087 ;
      RECT 22.94 305.967 23.14 306.087 ;
      RECT 24.02 305.498 24.22 305.618 ;
      RECT 24.38 283.087 24.58 283.207 ;
      RECT 23.66 283.087 23.86 283.207 ;
      RECT 22.94 283.087 23.14 283.207 ;
      RECT 20.78 283.087 20.98 283.207 ;
      RECT 24.38 278.76 24.58 278.88 ;
      RECT 23.66 278.76 23.86 278.88 ;
      RECT 22.94 278.76 23.14 278.88 ;
      RECT 20.78 278.76 20.98 278.88 ;
      RECT 23.3 278.13 23.5 278.25 ;
      RECT 24.38 277.5 24.58 277.62 ;
      RECT 23.66 277.5 23.86 277.62 ;
      RECT 22.94 277.5 23.14 277.62 ;
      RECT 20.78 277.5 20.98 277.62 ;
      RECT 23.3 276.87 23.5 276.99 ;
      RECT 24.38 276.24 24.58 276.36 ;
      RECT 23.66 276.24 23.86 276.36 ;
      RECT 22.94 276.24 23.14 276.36 ;
      RECT 20.78 276.24 20.98 276.36 ;
      RECT 23.3 275.61 23.5 275.73 ;
      RECT 24.38 274.98 24.58 275.1 ;
      RECT 23.66 274.98 23.86 275.1 ;
      RECT 22.94 274.98 23.14 275.1 ;
      RECT 20.78 274.98 20.98 275.1 ;
      RECT 23.3 274.35 23.5 274.47 ;
      RECT 24.38 273.72 24.58 273.84 ;
      RECT 23.66 273.72 23.86 273.84 ;
      RECT 22.94 273.72 23.14 273.84 ;
      RECT 23.3 273.09 23.5 273.21 ;
      RECT 20.78 273.72 20.98 273.84 ;
      RECT 24.38 272.46 24.58 272.58 ;
      RECT 23.66 272.46 23.86 272.58 ;
      RECT 22.94 272.46 23.14 272.58 ;
      RECT 23.3 271.83 23.5 271.95 ;
      RECT 20.78 272.46 20.98 272.58 ;
      RECT 20.78 271.2 20.98 271.32 ;
      RECT 23.3 270.57 23.5 270.69 ;
      RECT 22.94 271.2 23.14 271.32 ;
      RECT 23.66 271.2 23.86 271.32 ;
      RECT 24.38 271.2 24.58 271.32 ;
      RECT 20.78 269.94 20.98 270.06 ;
      RECT 23.3 269.31 23.5 269.43 ;
      RECT 22.94 269.94 23.14 270.06 ;
      RECT 23.66 269.94 23.86 270.06 ;
      RECT 24.38 269.94 24.58 270.06 ;
      RECT 20.78 268.68 20.98 268.8 ;
      RECT 23.3 268.05 23.5 268.17 ;
      RECT 22.94 268.68 23.14 268.8 ;
      RECT 23.66 268.68 23.86 268.8 ;
      RECT 24.38 268.68 24.58 268.8 ;
      RECT 20.78 267.42 20.98 267.54 ;
      RECT 23.3 266.79 23.5 266.91 ;
      RECT 22.94 267.42 23.14 267.54 ;
      RECT 23.66 267.42 23.86 267.54 ;
      RECT 24.38 267.42 24.58 267.54 ;
      RECT 20.78 266.16 20.98 266.28 ;
      RECT 20.78 264.9 20.98 265.02 ;
      RECT 22.94 264.9 23.14 265.02 ;
      RECT 23.66 264.9 23.86 265.02 ;
      RECT 24.38 264.9 24.58 265.02 ;
      RECT 23.3 265.53 23.5 265.65 ;
      RECT 22.94 266.16 23.14 266.28 ;
      RECT 23.66 266.16 23.86 266.28 ;
      RECT 24.38 266.16 24.58 266.28 ;
      RECT 20.78 263.64 20.98 263.76 ;
      RECT 22.94 263.64 23.14 263.76 ;
      RECT 23.66 263.64 23.86 263.76 ;
      RECT 24.38 263.64 24.58 263.76 ;
      RECT 23.3 264.27 23.5 264.39 ;
      RECT 20.78 262.38 20.98 262.5 ;
      RECT 22.94 262.38 23.14 262.5 ;
      RECT 23.66 262.38 23.86 262.5 ;
      RECT 24.38 262.38 24.58 262.5 ;
      RECT 23.3 263.01 23.5 263.13 ;
      RECT 20.78 261.12 20.98 261.24 ;
      RECT 22.94 261.12 23.14 261.24 ;
      RECT 23.66 261.12 23.86 261.24 ;
      RECT 24.38 261.12 24.58 261.24 ;
      RECT 23.3 261.75 23.5 261.87 ;
      RECT 20.78 259.86 20.98 259.98 ;
      RECT 22.94 259.86 23.14 259.98 ;
      RECT 23.66 259.86 23.86 259.98 ;
      RECT 24.38 259.86 24.58 259.98 ;
      RECT 23.3 260.49 23.5 260.61 ;
      RECT 20.78 258.6 20.98 258.72 ;
      RECT 22.94 258.6 23.14 258.72 ;
      RECT 23.66 258.6 23.86 258.72 ;
      RECT 24.38 258.6 24.58 258.72 ;
      RECT 23.3 259.23 23.5 259.35 ;
      RECT 20.78 257.34 20.98 257.46 ;
      RECT 25.46 162.6 25.66 162.72 ;
      RECT 25.82 163.62 26.02 163.74 ;
      RECT 25.1 163.62 25.3 163.74 ;
      RECT 26.54 161.1 26.74 161.22 ;
      RECT 25.82 161.1 26.02 161.22 ;
      RECT 25.1 161.1 25.3 161.22 ;
      RECT 25.46 160.08 25.66 160.2 ;
      RECT 25.82 158.58 26.02 158.7 ;
      RECT 26.54 158.82 26.74 158.94 ;
      RECT 25.1 158.82 25.3 158.94 ;
      RECT 25.46 157.56 25.66 157.68 ;
      RECT 26.18 158.038 26.38 158.158 ;
      RECT 24.74 158.278 24.94 158.398 ;
      RECT 25.82 156.06 26.02 156.18 ;
      RECT 26.54 156.3 26.74 156.42 ;
      RECT 25.1 156.3 25.3 156.42 ;
      RECT 24.74 156.842 24.94 156.962 ;
      RECT 26.18 156.842 26.38 156.962 ;
      RECT 25.46 154.8 25.66 154.92 ;
      RECT 25.1 153.54 25.3 153.66 ;
      RECT 26.54 153.78 26.74 153.9 ;
      RECT 25.82 153.78 26.02 153.9 ;
      RECT 25.46 152.52 25.66 152.64 ;
      RECT 25.1 151.26 25.3 151.38 ;
      RECT 25.82 151.26 26.02 151.38 ;
      RECT 26.54 151.26 26.74 151.38 ;
      RECT 25.46 150 25.66 150.12 ;
      RECT 26.54 148.5 26.74 148.62 ;
      RECT 25.82 148.74 26.02 148.86 ;
      RECT 25.1 148.74 25.3 148.86 ;
      RECT 25.46 144.72 25.66 144.84 ;
      RECT 26.54 145.98 26.74 146.1 ;
      RECT 25.82 145.98 26.02 146.1 ;
      RECT 25.1 145.98 25.3 146.1 ;
      RECT 25.82 143.46 26.02 143.58 ;
      RECT 25.1 143.7 25.3 143.82 ;
      RECT 26.54 143.7 26.74 143.82 ;
      RECT 25.46 142.2 25.66 142.32 ;
      RECT 25.82 140.94 26.02 141.06 ;
      RECT 25.1 141.18 25.3 141.3 ;
      RECT 26.54 141.18 26.74 141.3 ;
      RECT 25.46 139.92 25.66 140.04 ;
      RECT 25.1 138.42 25.3 138.54 ;
      RECT 26.54 138.42 26.74 138.54 ;
      RECT 25.82 138.66 26.02 138.78 ;
      RECT 26.54 139.138 26.74 139.258 ;
      RECT 25.82 139.138 26.02 139.258 ;
      RECT 25.1 139.138 25.3 139.258 ;
      RECT 26.54 136.618 26.74 136.738 ;
      RECT 25.82 136.618 26.02 136.738 ;
      RECT 25.1 136.618 25.3 136.738 ;
      RECT 25.46 137.4 25.66 137.52 ;
      RECT 25.1 135.9 25.3 136.02 ;
      RECT 26.54 135.9 26.74 136.02 ;
      RECT 25.82 136.14 26.02 136.26 ;
      RECT 26.54 134.098 26.74 134.218 ;
      RECT 25.82 134.098 26.02 134.218 ;
      RECT 25.1 134.098 25.3 134.218 ;
      RECT 25.46 134.64 25.66 134.76 ;
      RECT 26.54 133.38 26.74 133.5 ;
      RECT 25.82 133.62 26.02 133.74 ;
      RECT 25.1 133.62 25.3 133.74 ;
      RECT 25.1 131.1 25.3 131.22 ;
      RECT 25.82 131.1 26.02 131.22 ;
      RECT 26.54 131.578 26.74 131.698 ;
      RECT 25.82 131.578 26.02 131.698 ;
      RECT 25.1 131.578 25.3 131.698 ;
      RECT 25.46 132.36 25.66 132.48 ;
      RECT 26.54 130.86 26.74 130.98 ;
      RECT 25.1 129.058 25.3 129.178 ;
      RECT 25.82 129.058 26.02 129.178 ;
      RECT 26.54 129.058 26.74 129.178 ;
      RECT 26.54 128.58 26.74 128.7 ;
      RECT 25.1 128.58 25.3 128.7 ;
      RECT 25.82 128.34 26.02 128.46 ;
      RECT 25.46 129.6 25.66 129.72 ;
      RECT 25.46 127.08 25.66 127.2 ;
      RECT 25.1 126.538 25.3 126.658 ;
      RECT 25.82 126.538 26.02 126.658 ;
      RECT 26.54 126.538 26.74 126.658 ;
      RECT 25.82 126.06 26.02 126.18 ;
      RECT 25.1 125.82 25.3 125.94 ;
      RECT 26.54 125.82 26.74 125.94 ;
      RECT 25.46 124.56 25.66 124.68 ;
      RECT 25.1 124.018 25.3 124.138 ;
      RECT 25.82 124.018 26.02 124.138 ;
      RECT 26.54 124.018 26.74 124.138 ;
      RECT 25.82 123.54 26.02 123.66 ;
      RECT 26.54 123.54 26.74 123.66 ;
      RECT 25.1 123.3 25.3 123.42 ;
      RECT 25.46 122.04 25.66 122.16 ;
      RECT 25.1 121.498 25.3 121.618 ;
      RECT 25.82 121.498 26.02 121.618 ;
      RECT 26.54 121.498 26.74 121.618 ;
      RECT 25.1 121.02 25.3 121.14 ;
      RECT 26.54 121.02 26.74 121.14 ;
      RECT 25.82 120.78 26.02 120.9 ;
      RECT 25.46 119.52 25.66 119.64 ;
      RECT 25.1 118.978 25.3 119.098 ;
      RECT 25.82 118.978 26.02 119.098 ;
      RECT 26.54 118.978 26.74 119.098 ;
      RECT 25.82 118.5 26.02 118.62 ;
      RECT 26.18 212.61 26.38 212.73 ;
      RECT 24.74 212.61 24.94 212.73 ;
      RECT 26.54 210.72 26.74 210.84 ;
      RECT 25.82 210.72 26.02 210.84 ;
      RECT 25.1 210.72 25.3 210.84 ;
      RECT 26.18 211.35 26.38 211.47 ;
      RECT 24.74 211.35 24.94 211.47 ;
      RECT 25.1 209.46 25.3 209.58 ;
      RECT 25.82 209.46 26.02 209.58 ;
      RECT 26.54 209.46 26.74 209.58 ;
      RECT 24.74 210.09 24.94 210.21 ;
      RECT 26.18 210.09 26.38 210.21 ;
      RECT 25.46 207.96 25.66 208.08 ;
      RECT 26.18 208.262 26.38 208.382 ;
      RECT 24.74 208.502 24.94 208.622 ;
      RECT 26.54 206.46 26.74 206.58 ;
      RECT 25.1 206.7 25.3 206.82 ;
      RECT 25.82 206.7 26.02 206.82 ;
      RECT 25.46 205.44 25.66 205.56 ;
      RECT 26.18 205.742 26.38 205.862 ;
      RECT 24.74 205.982 24.94 206.102 ;
      RECT 24.74 203.462 24.94 203.582 ;
      RECT 25.82 203.94 26.02 204.06 ;
      RECT 26.54 204.18 26.74 204.3 ;
      RECT 25.1 204.18 25.3 204.3 ;
      RECT 25.46 202.92 25.66 203.04 ;
      RECT 26.18 203.222 26.38 203.342 ;
      RECT 26.18 200.702 26.38 200.822 ;
      RECT 24.74 200.942 24.94 201.062 ;
      RECT 25.1 201.42 25.3 201.54 ;
      RECT 25.82 201.66 26.02 201.78 ;
      RECT 26.54 201.66 26.74 201.78 ;
      RECT 25.46 200.4 25.66 200.52 ;
      RECT 26.18 198.182 26.38 198.302 ;
      RECT 24.74 198.422 24.94 198.542 ;
      RECT 26.54 198.9 26.74 199.02 ;
      RECT 25.82 199.14 26.02 199.26 ;
      RECT 25.1 199.14 25.3 199.26 ;
      RECT 25.1 196.62 25.3 196.74 ;
      RECT 25.82 196.62 26.02 196.74 ;
      RECT 25.46 197.88 25.66 198 ;
      RECT 25.46 195.36 25.66 195.48 ;
      RECT 24.74 195.902 24.94 196.022 ;
      RECT 26.18 195.902 26.38 196.022 ;
      RECT 26.54 196.38 26.74 196.5 ;
      RECT 25.82 193.86 26.02 193.98 ;
      RECT 25.1 194.1 25.3 194.22 ;
      RECT 26.54 194.1 26.74 194.22 ;
      RECT 26.18 194.402 26.38 194.522 ;
      RECT 24.74 194.642 24.94 194.762 ;
      RECT 25.46 192.6 25.66 192.72 ;
      RECT 24.74 193.142 24.94 193.262 ;
      RECT 26.18 193.382 26.38 193.502 ;
      RECT 26.54 191.34 26.74 191.46 ;
      RECT 25.1 191.58 25.3 191.7 ;
      RECT 25.82 191.58 26.02 191.7 ;
      RECT 24.74 191.882 24.94 192.002 ;
      RECT 26.18 192.122 26.38 192.242 ;
      RECT 25.46 190.08 25.66 190.2 ;
      RECT 24.74 190.622 24.94 190.742 ;
      RECT 26.18 190.862 26.38 190.982 ;
      RECT 26.54 189.06 26.74 189.18 ;
      RECT 25.82 189.06 26.02 189.18 ;
      RECT 25.1 189.06 25.3 189.18 ;
      RECT 25.46 187.56 25.66 187.68 ;
      RECT 26.54 186.54 26.74 186.66 ;
      RECT 25.82 186.54 26.02 186.66 ;
      RECT 25.1 186.54 25.3 186.66 ;
      RECT 25.46 185.04 25.66 185.16 ;
      RECT 26.54 183.78 26.74 183.9 ;
      RECT 25.1 184.02 25.3 184.14 ;
      RECT 25.82 184.02 26.02 184.14 ;
      RECT 25.46 182.76 25.66 182.88 ;
      RECT 25.46 180.24 25.66 180.36 ;
      RECT 25.82 181.26 26.02 181.38 ;
      RECT 26.54 181.5 26.74 181.62 ;
      RECT 25.1 181.5 25.3 181.62 ;
      RECT 26.54 178.98 26.74 179.1 ;
      RECT 25.1 178.98 25.3 179.1 ;
      RECT 25.46 177.48 25.66 177.6 ;
      RECT 25.82 178.74 26.02 178.86 ;
      RECT 25.82 176.22 26.02 176.34 ;
      RECT 25.1 176.46 25.3 176.58 ;
      RECT 26.54 176.46 26.74 176.58 ;
      RECT 25.46 174.96 25.66 175.08 ;
      RECT 26.54 173.7 26.74 173.82 ;
      RECT 25.1 173.94 25.3 174.06 ;
      RECT 25.82 173.94 26.02 174.06 ;
      RECT 25.46 172.44 25.66 172.56 ;
      RECT 25.82 171.18 26.02 171.3 ;
      RECT 25.1 171.42 25.3 171.54 ;
      RECT 26.54 171.42 26.74 171.54 ;
      RECT 25.46 170.16 25.66 170.28 ;
      RECT 26.54 168.66 26.74 168.78 ;
      RECT 25.1 168.66 25.3 168.78 ;
      RECT 25.82 168.9 26.02 169.02 ;
      RECT 25.46 167.64 25.66 167.76 ;
      RECT 26.54 166.14 26.74 166.26 ;
      RECT 25.1 166.38 25.3 166.5 ;
      RECT 25.82 166.38 26.02 166.5 ;
      RECT 26.54 163.86 26.74 163.98 ;
      RECT 25.46 164.88 25.66 165 ;
      RECT 25.1 238.44 25.3 238.56 ;
      RECT 24.74 236.55 24.94 236.67 ;
      RECT 26.18 236.55 26.38 236.67 ;
      RECT 26.54 237.18 26.74 237.3 ;
      RECT 25.82 237.18 26.02 237.3 ;
      RECT 25.1 237.18 25.3 237.3 ;
      RECT 24.74 235.29 24.94 235.41 ;
      RECT 26.18 235.29 26.38 235.41 ;
      RECT 25.1 235.92 25.3 236.04 ;
      RECT 25.82 235.92 26.02 236.04 ;
      RECT 26.54 235.92 26.74 236.04 ;
      RECT 26.18 234.03 26.38 234.15 ;
      RECT 24.74 234.03 24.94 234.15 ;
      RECT 25.1 234.66 25.3 234.78 ;
      RECT 25.82 234.66 26.02 234.78 ;
      RECT 26.54 234.66 26.74 234.78 ;
      RECT 25.1 232.14 25.3 232.26 ;
      RECT 25.82 232.14 26.02 232.26 ;
      RECT 26.54 232.14 26.74 232.26 ;
      RECT 24.74 232.77 24.94 232.89 ;
      RECT 26.18 232.77 26.38 232.89 ;
      RECT 26.54 233.4 26.74 233.52 ;
      RECT 25.82 233.4 26.02 233.52 ;
      RECT 25.1 233.4 25.3 233.52 ;
      RECT 25.1 230.88 25.3 231 ;
      RECT 25.82 230.88 26.02 231 ;
      RECT 26.54 230.88 26.74 231 ;
      RECT 24.74 231.51 24.94 231.63 ;
      RECT 26.18 231.51 26.38 231.63 ;
      RECT 26.54 229.62 26.74 229.74 ;
      RECT 25.82 229.62 26.02 229.74 ;
      RECT 25.1 229.62 25.3 229.74 ;
      RECT 24.74 230.25 24.94 230.37 ;
      RECT 26.18 230.25 26.38 230.37 ;
      RECT 26.54 228.36 26.74 228.48 ;
      RECT 25.82 228.36 26.02 228.48 ;
      RECT 25.1 228.36 25.3 228.48 ;
      RECT 26.18 228.99 26.38 229.11 ;
      RECT 24.74 228.99 24.94 229.11 ;
      RECT 26.54 227.1 26.74 227.22 ;
      RECT 25.82 227.1 26.02 227.22 ;
      RECT 25.1 227.1 25.3 227.22 ;
      RECT 26.18 227.73 26.38 227.85 ;
      RECT 24.74 227.73 24.94 227.85 ;
      RECT 26.54 225.84 26.74 225.96 ;
      RECT 25.82 225.84 26.02 225.96 ;
      RECT 25.1 225.84 25.3 225.96 ;
      RECT 26.18 226.47 26.38 226.59 ;
      RECT 24.74 226.47 24.94 226.59 ;
      RECT 26.18 223.95 26.38 224.07 ;
      RECT 24.74 223.95 24.94 224.07 ;
      RECT 26.54 224.58 26.74 224.7 ;
      RECT 25.82 224.58 26.02 224.7 ;
      RECT 25.1 224.58 25.3 224.7 ;
      RECT 26.18 225.21 26.38 225.33 ;
      RECT 24.74 225.21 24.94 225.33 ;
      RECT 26.18 222.69 26.38 222.81 ;
      RECT 24.74 222.69 24.94 222.81 ;
      RECT 26.54 223.32 26.74 223.44 ;
      RECT 25.82 223.32 26.02 223.44 ;
      RECT 25.1 223.32 25.3 223.44 ;
      RECT 26.18 221.43 26.38 221.55 ;
      RECT 24.74 221.43 24.94 221.55 ;
      RECT 26.54 222.06 26.74 222.18 ;
      RECT 25.82 222.06 26.02 222.18 ;
      RECT 25.1 222.06 25.3 222.18 ;
      RECT 26.54 220.8 26.74 220.92 ;
      RECT 25.82 220.8 26.02 220.92 ;
      RECT 25.1 220.8 25.3 220.92 ;
      RECT 24.74 220.17 24.94 220.29 ;
      RECT 26.18 220.17 26.38 220.29 ;
      RECT 26.18 218.91 26.38 219.03 ;
      RECT 24.74 218.91 24.94 219.03 ;
      RECT 25.1 219.54 25.3 219.66 ;
      RECT 25.82 219.54 26.02 219.66 ;
      RECT 26.54 219.54 26.74 219.66 ;
      RECT 26.18 217.65 26.38 217.77 ;
      RECT 24.74 217.65 24.94 217.77 ;
      RECT 25.82 218.28 26.02 218.4 ;
      RECT 26.54 218.28 26.74 218.4 ;
      RECT 25.1 218.28 25.3 218.4 ;
      RECT 26.54 215.76 26.74 215.88 ;
      RECT 25.82 215.76 26.02 215.88 ;
      RECT 25.1 215.76 25.3 215.88 ;
      RECT 24.74 216.39 24.94 216.51 ;
      RECT 26.18 216.39 26.38 216.51 ;
      RECT 26.54 217.02 26.74 217.14 ;
      RECT 25.82 217.02 26.02 217.14 ;
      RECT 25.1 217.02 25.3 217.14 ;
      RECT 25.1 214.5 25.3 214.62 ;
      RECT 25.82 214.5 26.02 214.62 ;
      RECT 26.54 214.5 26.74 214.62 ;
      RECT 26.18 215.13 26.38 215.25 ;
      RECT 24.74 215.13 24.94 215.25 ;
      RECT 25.1 213.24 25.3 213.36 ;
      RECT 25.82 213.24 26.02 213.36 ;
      RECT 26.54 213.24 26.74 213.36 ;
      RECT 26.18 213.87 26.38 213.99 ;
      RECT 24.74 213.87 24.94 213.99 ;
      RECT 25.1 211.98 25.3 212.1 ;
      RECT 25.82 211.98 26.02 212.1 ;
      RECT 26.54 211.98 26.74 212.1 ;
      RECT 26.18 264.27 26.38 264.39 ;
      RECT 25.1 262.38 25.3 262.5 ;
      RECT 25.82 262.38 26.02 262.5 ;
      RECT 26.54 262.38 26.74 262.5 ;
      RECT 24.74 263.01 24.94 263.13 ;
      RECT 26.18 263.01 26.38 263.13 ;
      RECT 25.1 261.12 25.3 261.24 ;
      RECT 25.82 261.12 26.02 261.24 ;
      RECT 26.54 261.12 26.74 261.24 ;
      RECT 24.74 261.75 24.94 261.87 ;
      RECT 26.18 261.75 26.38 261.87 ;
      RECT 25.1 259.86 25.3 259.98 ;
      RECT 25.82 259.86 26.02 259.98 ;
      RECT 26.54 259.86 26.74 259.98 ;
      RECT 26.18 260.49 26.38 260.61 ;
      RECT 24.74 260.49 24.94 260.61 ;
      RECT 25.1 258.6 25.3 258.72 ;
      RECT 25.82 258.6 26.02 258.72 ;
      RECT 26.54 258.6 26.74 258.72 ;
      RECT 24.74 259.23 24.94 259.35 ;
      RECT 26.18 259.23 26.38 259.35 ;
      RECT 24.74 256.71 24.94 256.83 ;
      RECT 26.18 256.71 26.38 256.83 ;
      RECT 25.1 257.34 25.3 257.46 ;
      RECT 25.82 257.34 26.02 257.46 ;
      RECT 26.54 257.34 26.74 257.46 ;
      RECT 24.74 257.97 24.94 258.09 ;
      RECT 26.18 257.97 26.38 258.09 ;
      RECT 24.74 255.45 24.94 255.57 ;
      RECT 26.18 255.45 26.38 255.57 ;
      RECT 25.1 256.08 25.3 256.2 ;
      RECT 25.82 256.08 26.02 256.2 ;
      RECT 26.54 256.08 26.74 256.2 ;
      RECT 24.74 254.19 24.94 254.31 ;
      RECT 26.18 254.19 26.38 254.31 ;
      RECT 25.1 254.82 25.3 254.94 ;
      RECT 25.82 254.82 26.02 254.94 ;
      RECT 26.54 254.82 26.74 254.94 ;
      RECT 24.74 252.93 24.94 253.05 ;
      RECT 26.18 252.93 26.38 253.05 ;
      RECT 25.1 253.56 25.3 253.68 ;
      RECT 25.82 253.56 26.02 253.68 ;
      RECT 26.54 253.56 26.74 253.68 ;
      RECT 24.74 251.67 24.94 251.79 ;
      RECT 26.18 251.67 26.38 251.79 ;
      RECT 25.1 252.3 25.3 252.42 ;
      RECT 25.82 252.3 26.02 252.42 ;
      RECT 26.54 252.3 26.74 252.42 ;
      RECT 24.74 250.41 24.94 250.53 ;
      RECT 26.18 250.41 26.38 250.53 ;
      RECT 25.1 251.04 25.3 251.16 ;
      RECT 25.82 251.04 26.02 251.16 ;
      RECT 26.54 251.04 26.74 251.16 ;
      RECT 25.1 248.52 25.3 248.64 ;
      RECT 25.82 248.52 26.02 248.64 ;
      RECT 26.54 248.52 26.74 248.64 ;
      RECT 24.74 249.15 24.94 249.27 ;
      RECT 26.18 249.15 26.38 249.27 ;
      RECT 25.1 249.78 25.3 249.9 ;
      RECT 25.82 249.78 26.02 249.9 ;
      RECT 26.54 249.78 26.74 249.9 ;
      RECT 25.1 247.26 25.3 247.38 ;
      RECT 25.82 247.26 26.02 247.38 ;
      RECT 26.54 247.26 26.74 247.38 ;
      RECT 24.74 247.89 24.94 248.01 ;
      RECT 26.18 247.89 26.38 248.01 ;
      RECT 24.74 246.63 24.94 246.75 ;
      RECT 26.18 246.63 26.38 246.75 ;
      RECT 26.54 246 26.74 246.12 ;
      RECT 25.82 246 26.02 246.12 ;
      RECT 25.1 246 25.3 246.12 ;
      RECT 26.54 244.74 26.74 244.86 ;
      RECT 25.82 244.74 26.02 244.86 ;
      RECT 25.1 244.74 25.3 244.86 ;
      RECT 26.18 245.37 26.38 245.49 ;
      RECT 24.74 245.37 24.94 245.49 ;
      RECT 25.1 243.48 25.3 243.6 ;
      RECT 25.82 243.48 26.02 243.6 ;
      RECT 26.54 243.48 26.74 243.6 ;
      RECT 24.74 244.11 24.94 244.23 ;
      RECT 26.18 244.11 26.38 244.23 ;
      RECT 25.1 242.22 25.3 242.34 ;
      RECT 25.82 242.22 26.02 242.34 ;
      RECT 26.54 242.22 26.74 242.34 ;
      RECT 24.74 242.85 24.94 242.97 ;
      RECT 26.18 242.85 26.38 242.97 ;
      RECT 24.74 240.33 24.94 240.45 ;
      RECT 26.18 240.33 26.38 240.45 ;
      RECT 26.54 240.96 26.74 241.08 ;
      RECT 25.82 240.96 26.02 241.08 ;
      RECT 25.1 240.96 25.3 241.08 ;
      RECT 26.18 241.59 26.38 241.71 ;
      RECT 24.74 241.59 24.94 241.71 ;
      RECT 24.74 239.07 24.94 239.19 ;
      RECT 26.18 239.07 26.38 239.19 ;
      RECT 25.1 239.7 25.3 239.82 ;
      RECT 25.82 239.7 26.02 239.82 ;
      RECT 26.54 239.7 26.74 239.82 ;
      RECT 26.18 237.81 26.38 237.93 ;
      RECT 24.74 237.81 24.94 237.93 ;
      RECT 25.82 238.44 26.02 238.56 ;
      RECT 26.54 238.44 26.74 238.56 ;
      RECT 29.78 122.28 29.98 122.4 ;
      RECT 31.22 122.04 31.42 122.16 ;
      RECT 28.7 121.498 28.9 121.618 ;
      RECT 29.42 121.498 29.62 121.618 ;
      RECT 30.14 121.498 30.34 121.618 ;
      RECT 30.86 121.498 31.06 121.618 ;
      RECT 31.58 121.498 31.78 121.618 ;
      RECT 32.3 121.498 32.5 121.618 ;
      RECT 29.42 121.02 29.62 121.14 ;
      RECT 30.86 121.02 31.06 121.14 ;
      RECT 32.3 121.02 32.5 121.14 ;
      RECT 28.7 120.78 28.9 120.9 ;
      RECT 30.14 120.78 30.34 120.9 ;
      RECT 31.58 120.78 31.78 120.9 ;
      RECT 29.78 119.76 29.98 119.88 ;
      RECT 31.22 119.52 31.42 119.64 ;
      RECT 28.7 118.978 28.9 119.098 ;
      RECT 29.42 118.978 29.62 119.098 ;
      RECT 30.14 118.978 30.34 119.098 ;
      RECT 30.86 118.978 31.06 119.098 ;
      RECT 31.58 118.978 31.78 119.098 ;
      RECT 32.3 118.978 32.5 119.098 ;
      RECT 32.3 118.5 32.5 118.62 ;
      RECT 31.58 118.5 31.78 118.62 ;
      RECT 30.14 118.5 30.34 118.62 ;
      RECT 29.42 118.5 29.62 118.62 ;
      RECT 28.7 118.5 28.9 118.62 ;
      RECT 30.86 118.26 31.06 118.38 ;
      RECT 25.46 348.339 25.66 348.459 ;
      RECT 26.54 325.9425 26.74 326.0625 ;
      RECT 25.82 325.9425 26.02 326.0625 ;
      RECT 25.1 325.9425 25.3 326.0625 ;
      RECT 25.46 323.3835 25.66 323.5035 ;
      RECT 26.54 305.967 26.74 306.087 ;
      RECT 25.82 305.967 26.02 306.087 ;
      RECT 25.1 305.967 25.3 306.087 ;
      RECT 25.46 305.498 25.66 305.618 ;
      RECT 26.54 283.087 26.74 283.207 ;
      RECT 25.82 283.087 26.02 283.207 ;
      RECT 25.1 283.087 25.3 283.207 ;
      RECT 26.54 278.76 26.74 278.88 ;
      RECT 25.82 278.76 26.02 278.88 ;
      RECT 25.1 278.76 25.3 278.88 ;
      RECT 26.18 278.13 26.38 278.25 ;
      RECT 24.74 278.13 24.94 278.25 ;
      RECT 26.54 277.5 26.74 277.62 ;
      RECT 25.82 277.5 26.02 277.62 ;
      RECT 25.1 277.5 25.3 277.62 ;
      RECT 26.18 276.87 26.38 276.99 ;
      RECT 24.74 276.87 24.94 276.99 ;
      RECT 26.54 276.24 26.74 276.36 ;
      RECT 25.82 276.24 26.02 276.36 ;
      RECT 25.1 276.24 25.3 276.36 ;
      RECT 26.18 275.61 26.38 275.73 ;
      RECT 24.74 275.61 24.94 275.73 ;
      RECT 26.54 274.98 26.74 275.1 ;
      RECT 25.82 274.98 26.02 275.1 ;
      RECT 25.1 274.98 25.3 275.1 ;
      RECT 26.18 274.35 26.38 274.47 ;
      RECT 24.74 274.35 24.94 274.47 ;
      RECT 26.54 273.72 26.74 273.84 ;
      RECT 25.82 273.72 26.02 273.84 ;
      RECT 25.1 273.72 25.3 273.84 ;
      RECT 26.18 273.09 26.38 273.21 ;
      RECT 24.74 273.09 24.94 273.21 ;
      RECT 26.54 272.46 26.74 272.58 ;
      RECT 25.82 272.46 26.02 272.58 ;
      RECT 25.1 272.46 25.3 272.58 ;
      RECT 26.18 271.83 26.38 271.95 ;
      RECT 24.74 271.83 24.94 271.95 ;
      RECT 24.74 270.57 24.94 270.69 ;
      RECT 26.18 270.57 26.38 270.69 ;
      RECT 25.1 271.2 25.3 271.32 ;
      RECT 25.82 271.2 26.02 271.32 ;
      RECT 26.54 271.2 26.74 271.32 ;
      RECT 24.74 269.31 24.94 269.43 ;
      RECT 26.18 269.31 26.38 269.43 ;
      RECT 25.1 269.94 25.3 270.06 ;
      RECT 25.82 269.94 26.02 270.06 ;
      RECT 26.54 269.94 26.74 270.06 ;
      RECT 24.74 268.05 24.94 268.17 ;
      RECT 26.18 268.05 26.38 268.17 ;
      RECT 25.1 268.68 25.3 268.8 ;
      RECT 25.82 268.68 26.02 268.8 ;
      RECT 26.54 268.68 26.74 268.8 ;
      RECT 24.74 266.79 24.94 266.91 ;
      RECT 26.18 266.79 26.38 266.91 ;
      RECT 25.1 267.42 25.3 267.54 ;
      RECT 25.82 267.42 26.02 267.54 ;
      RECT 26.54 267.42 26.74 267.54 ;
      RECT 25.1 264.9 25.3 265.02 ;
      RECT 25.82 264.9 26.02 265.02 ;
      RECT 26.54 264.9 26.74 265.02 ;
      RECT 24.74 265.53 24.94 265.65 ;
      RECT 26.18 265.53 26.38 265.65 ;
      RECT 25.1 266.16 25.3 266.28 ;
      RECT 25.82 266.16 26.02 266.28 ;
      RECT 26.54 266.16 26.74 266.28 ;
      RECT 25.1 263.64 25.3 263.76 ;
      RECT 25.82 263.64 26.02 263.76 ;
      RECT 26.54 263.64 26.74 263.76 ;
      RECT 24.74 264.27 24.94 264.39 ;
      RECT 28.7 140.94 28.9 141.06 ;
      RECT 29.42 141.18 29.62 141.3 ;
      RECT 30.86 141.18 31.06 141.3 ;
      RECT 31.58 141.18 31.78 141.3 ;
      RECT 29.78 139.68 29.98 139.8 ;
      RECT 31.22 139.92 31.42 140.04 ;
      RECT 29.42 138.42 29.62 138.54 ;
      RECT 31.58 138.42 31.78 138.54 ;
      RECT 32.3 138.66 32.5 138.78 ;
      RECT 30.86 138.66 31.06 138.78 ;
      RECT 30.14 138.66 30.34 138.78 ;
      RECT 28.7 138.66 28.9 138.78 ;
      RECT 32.3 139.138 32.5 139.258 ;
      RECT 31.58 139.138 31.78 139.258 ;
      RECT 30.86 139.138 31.06 139.258 ;
      RECT 30.14 139.138 30.34 139.258 ;
      RECT 29.42 139.138 29.62 139.258 ;
      RECT 28.7 139.138 28.9 139.258 ;
      RECT 32.3 136.618 32.5 136.738 ;
      RECT 31.58 136.618 31.78 136.738 ;
      RECT 30.86 136.618 31.06 136.738 ;
      RECT 30.14 136.618 30.34 136.738 ;
      RECT 29.42 136.618 29.62 136.738 ;
      RECT 28.7 136.618 28.9 136.738 ;
      RECT 29.78 137.16 29.98 137.28 ;
      RECT 31.22 137.4 31.42 137.52 ;
      RECT 29.42 135.9 29.62 136.02 ;
      RECT 30.86 135.9 31.06 136.02 ;
      RECT 32.3 135.9 32.5 136.02 ;
      RECT 28.7 136.14 28.9 136.26 ;
      RECT 30.14 136.14 30.34 136.26 ;
      RECT 31.58 136.14 31.78 136.26 ;
      RECT 32.3 134.098 32.5 134.218 ;
      RECT 31.58 134.098 31.78 134.218 ;
      RECT 30.86 134.098 31.06 134.218 ;
      RECT 30.14 134.098 30.34 134.218 ;
      RECT 29.42 134.098 29.62 134.218 ;
      RECT 28.7 134.098 28.9 134.218 ;
      RECT 29.78 134.88 29.98 135 ;
      RECT 31.22 134.88 31.42 135 ;
      RECT 29.42 133.38 29.62 133.5 ;
      RECT 30.86 133.38 31.06 133.5 ;
      RECT 32.3 133.62 32.5 133.74 ;
      RECT 31.58 133.62 31.78 133.74 ;
      RECT 30.14 133.62 30.34 133.74 ;
      RECT 28.7 133.62 28.9 133.74 ;
      RECT 28.7 131.1 28.9 131.22 ;
      RECT 30.14 131.1 30.34 131.22 ;
      RECT 30.86 131.1 31.06 131.22 ;
      RECT 31.58 131.1 31.78 131.22 ;
      RECT 32.3 131.578 32.5 131.698 ;
      RECT 31.58 131.578 31.78 131.698 ;
      RECT 30.86 131.578 31.06 131.698 ;
      RECT 30.14 131.578 30.34 131.698 ;
      RECT 29.42 131.578 29.62 131.698 ;
      RECT 28.7 131.578 28.9 131.698 ;
      RECT 29.78 132.12 29.98 132.24 ;
      RECT 31.22 132.36 31.42 132.48 ;
      RECT 29.78 129.84 29.98 129.96 ;
      RECT 32.3 130.86 32.5 130.98 ;
      RECT 29.42 130.86 29.62 130.98 ;
      RECT 28.7 129.058 28.9 129.178 ;
      RECT 29.42 129.058 29.62 129.178 ;
      RECT 30.14 129.058 30.34 129.178 ;
      RECT 30.86 129.058 31.06 129.178 ;
      RECT 31.58 129.058 31.78 129.178 ;
      RECT 32.3 129.058 32.5 129.178 ;
      RECT 32.3 128.58 32.5 128.7 ;
      RECT 30.86 128.58 31.06 128.7 ;
      RECT 29.42 128.58 29.62 128.7 ;
      RECT 31.58 128.34 31.78 128.46 ;
      RECT 30.14 128.34 30.34 128.46 ;
      RECT 28.7 128.34 28.9 128.46 ;
      RECT 31.22 129.6 31.42 129.72 ;
      RECT 29.78 127.32 29.98 127.44 ;
      RECT 31.22 127.08 31.42 127.2 ;
      RECT 28.7 126.538 28.9 126.658 ;
      RECT 29.42 126.538 29.62 126.658 ;
      RECT 30.14 126.538 30.34 126.658 ;
      RECT 30.86 126.538 31.06 126.658 ;
      RECT 31.58 126.538 31.78 126.658 ;
      RECT 32.3 126.538 32.5 126.658 ;
      RECT 28.7 126.06 28.9 126.18 ;
      RECT 30.14 126.06 30.34 126.18 ;
      RECT 31.58 126.06 31.78 126.18 ;
      RECT 32.3 126.06 32.5 126.18 ;
      RECT 29.42 125.82 29.62 125.94 ;
      RECT 30.86 125.82 31.06 125.94 ;
      RECT 29.78 124.8 29.98 124.92 ;
      RECT 31.22 124.56 31.42 124.68 ;
      RECT 28.7 124.018 28.9 124.138 ;
      RECT 29.42 124.018 29.62 124.138 ;
      RECT 30.14 124.018 30.34 124.138 ;
      RECT 30.86 124.018 31.06 124.138 ;
      RECT 31.58 124.018 31.78 124.138 ;
      RECT 32.3 124.018 32.5 124.138 ;
      RECT 28.7 123.54 28.9 123.66 ;
      RECT 30.14 123.54 30.34 123.66 ;
      RECT 31.58 123.54 31.78 123.66 ;
      RECT 32.3 123.54 32.5 123.66 ;
      RECT 29.42 123.3 29.62 123.42 ;
      RECT 30.86 123.3 31.06 123.42 ;
      RECT 30.86 171.18 31.06 171.3 ;
      RECT 28.7 171.18 28.9 171.3 ;
      RECT 29.42 171.42 29.62 171.54 ;
      RECT 30.14 171.42 30.34 171.54 ;
      RECT 31.58 171.42 31.78 171.54 ;
      RECT 32.3 171.42 32.5 171.54 ;
      RECT 29.78 170.16 29.98 170.28 ;
      RECT 31.22 170.16 31.42 170.28 ;
      RECT 32.3 168.66 32.5 168.78 ;
      RECT 31.58 168.66 31.78 168.78 ;
      RECT 30.14 168.66 30.34 168.78 ;
      RECT 28.7 168.9 28.9 169.02 ;
      RECT 29.42 168.9 29.62 169.02 ;
      RECT 30.86 168.9 31.06 169.02 ;
      RECT 31.22 167.4 31.42 167.52 ;
      RECT 29.78 167.64 29.98 167.76 ;
      RECT 30.14 166.14 30.34 166.26 ;
      RECT 30.86 166.14 31.06 166.26 ;
      RECT 32.3 166.14 32.5 166.26 ;
      RECT 28.7 166.38 28.9 166.5 ;
      RECT 29.42 166.38 29.62 166.5 ;
      RECT 31.58 166.38 31.78 166.5 ;
      RECT 29.42 163.86 29.62 163.98 ;
      RECT 30.86 163.86 31.06 163.98 ;
      RECT 31.58 163.86 31.78 163.98 ;
      RECT 29.78 165.12 29.98 165.24 ;
      RECT 31.22 165.12 31.42 165.24 ;
      RECT 29.78 162.6 29.98 162.72 ;
      RECT 31.22 162.6 31.42 162.72 ;
      RECT 32.3 163.62 32.5 163.74 ;
      RECT 30.14 163.62 30.34 163.74 ;
      RECT 28.7 163.62 28.9 163.74 ;
      RECT 32.3 161.1 32.5 161.22 ;
      RECT 31.58 161.1 31.78 161.22 ;
      RECT 30.86 161.1 31.06 161.22 ;
      RECT 30.14 161.1 30.34 161.22 ;
      RECT 29.42 161.1 29.62 161.22 ;
      RECT 28.7 161.1 28.9 161.22 ;
      RECT 29.78 159.84 29.98 159.96 ;
      RECT 31.22 160.08 31.42 160.2 ;
      RECT 32.3 158.58 32.5 158.7 ;
      RECT 30.86 158.58 31.06 158.7 ;
      RECT 29.42 158.58 29.62 158.7 ;
      RECT 31.58 158.82 31.78 158.94 ;
      RECT 30.14 158.82 30.34 158.94 ;
      RECT 28.7 158.82 28.9 158.94 ;
      RECT 31.22 157.32 31.42 157.44 ;
      RECT 29.78 157.56 29.98 157.68 ;
      RECT 30.5 158.038 30.7 158.158 ;
      RECT 29.06 158.278 29.26 158.398 ;
      RECT 31.94 158.278 32.14 158.398 ;
      RECT 28.7 156.06 28.9 156.18 ;
      RECT 30.14 156.06 30.34 156.18 ;
      RECT 31.58 156.06 31.78 156.18 ;
      RECT 32.3 156.3 32.5 156.42 ;
      RECT 30.86 156.3 31.06 156.42 ;
      RECT 29.42 156.3 29.62 156.42 ;
      RECT 29.06 156.602 29.26 156.722 ;
      RECT 31.94 156.602 32.14 156.722 ;
      RECT 30.5 156.842 30.7 156.962 ;
      RECT 31.22 154.8 31.42 154.92 ;
      RECT 29.78 155.04 29.98 155.16 ;
      RECT 28.7 153.54 28.9 153.66 ;
      RECT 32.3 153.54 32.5 153.66 ;
      RECT 30.14 153.78 30.34 153.9 ;
      RECT 30.86 153.78 31.06 153.9 ;
      RECT 31.58 153.78 31.78 153.9 ;
      RECT 29.42 153.78 29.62 153.9 ;
      RECT 29.78 152.28 29.98 152.4 ;
      RECT 31.22 152.52 31.42 152.64 ;
      RECT 28.7 151.02 28.9 151.14 ;
      RECT 31.58 151.02 31.78 151.14 ;
      RECT 29.42 151.26 29.62 151.38 ;
      RECT 30.14 151.26 30.34 151.38 ;
      RECT 30.86 151.26 31.06 151.38 ;
      RECT 32.3 151.26 32.5 151.38 ;
      RECT 29.78 149.76 29.98 149.88 ;
      RECT 31.22 150 31.42 150.12 ;
      RECT 30.86 148.5 31.06 148.62 ;
      RECT 32.3 148.5 32.5 148.62 ;
      RECT 31.58 148.74 31.78 148.86 ;
      RECT 30.14 148.74 30.34 148.86 ;
      RECT 29.42 148.74 29.62 148.86 ;
      RECT 28.7 148.74 28.9 148.86 ;
      RECT 31.22 144.72 31.42 144.84 ;
      RECT 29.78 144.96 29.98 145.08 ;
      RECT 32.3 145.98 32.5 146.1 ;
      RECT 31.58 145.98 31.78 146.1 ;
      RECT 30.86 145.98 31.06 146.1 ;
      RECT 30.14 145.98 30.34 146.1 ;
      RECT 29.42 145.98 29.62 146.1 ;
      RECT 28.7 145.98 28.9 146.1 ;
      RECT 28.7 143.46 28.9 143.58 ;
      RECT 30.14 143.46 30.34 143.58 ;
      RECT 31.58 143.46 31.78 143.58 ;
      RECT 29.42 143.7 29.62 143.82 ;
      RECT 30.86 143.7 31.06 143.82 ;
      RECT 32.3 143.7 32.5 143.82 ;
      RECT 31.22 142.2 31.42 142.32 ;
      RECT 29.78 142.44 29.98 142.56 ;
      RECT 32.3 140.94 32.5 141.06 ;
      RECT 30.14 140.94 30.34 141.06 ;
      RECT 30.5 190.862 30.7 190.982 ;
      RECT 29.42 188.82 29.62 188.94 ;
      RECT 30.86 188.82 31.06 188.94 ;
      RECT 32.3 188.82 32.5 188.94 ;
      RECT 31.58 189.06 31.78 189.18 ;
      RECT 30.14 189.06 30.34 189.18 ;
      RECT 28.7 189.06 28.9 189.18 ;
      RECT 31.22 187.56 31.42 187.68 ;
      RECT 29.78 187.8 29.98 187.92 ;
      RECT 31.58 186.3 31.78 186.42 ;
      RECT 30.14 186.3 30.34 186.42 ;
      RECT 29.42 186.3 29.62 186.42 ;
      RECT 32.3 186.54 32.5 186.66 ;
      RECT 30.86 186.54 31.06 186.66 ;
      RECT 28.7 186.54 28.9 186.66 ;
      RECT 31.22 185.04 31.42 185.16 ;
      RECT 29.78 185.28 29.98 185.4 ;
      RECT 28.7 183.78 28.9 183.9 ;
      RECT 30.14 183.78 30.34 183.9 ;
      RECT 29.42 184.02 29.62 184.14 ;
      RECT 30.86 184.02 31.06 184.14 ;
      RECT 31.58 184.02 31.78 184.14 ;
      RECT 32.3 184.02 32.5 184.14 ;
      RECT 29.78 182.52 29.98 182.64 ;
      RECT 31.22 182.76 31.42 182.88 ;
      RECT 29.78 180.24 29.98 180.36 ;
      RECT 30.14 181.26 30.34 181.38 ;
      RECT 32.3 181.26 32.5 181.38 ;
      RECT 31.58 181.5 31.78 181.62 ;
      RECT 30.86 181.5 31.06 181.62 ;
      RECT 29.42 181.5 29.62 181.62 ;
      RECT 28.7 181.5 28.9 181.62 ;
      RECT 31.58 178.98 31.78 179.1 ;
      RECT 30.86 178.98 31.06 179.1 ;
      RECT 29.42 178.98 29.62 179.1 ;
      RECT 28.7 178.98 28.9 179.1 ;
      RECT 31.22 180 31.42 180.12 ;
      RECT 31.22 177.48 31.42 177.6 ;
      RECT 29.78 177.72 29.98 177.84 ;
      RECT 30.14 178.74 30.34 178.86 ;
      RECT 32.3 178.74 32.5 178.86 ;
      RECT 32.3 176.22 32.5 176.34 ;
      RECT 28.7 176.46 28.9 176.58 ;
      RECT 29.42 176.46 29.62 176.58 ;
      RECT 30.14 176.46 30.34 176.58 ;
      RECT 30.86 176.46 31.06 176.58 ;
      RECT 31.58 176.46 31.78 176.58 ;
      RECT 31.22 175.2 31.42 175.32 ;
      RECT 29.78 175.2 29.98 175.32 ;
      RECT 31.58 173.7 31.78 173.82 ;
      RECT 32.3 173.7 32.5 173.82 ;
      RECT 28.7 173.94 28.9 174.06 ;
      RECT 29.42 173.94 29.62 174.06 ;
      RECT 30.14 173.94 30.34 174.06 ;
      RECT 30.86 173.94 31.06 174.06 ;
      RECT 31.22 172.44 31.42 172.56 ;
      RECT 29.78 172.68 29.98 172.8 ;
      RECT 29.78 190.32 29.98 190.44 ;
      RECT 31.94 190.622 32.14 190.742 ;
      RECT 29.06 190.622 29.26 190.742 ;
      RECT 32.3 204.18 32.5 204.3 ;
      RECT 30.86 204.18 31.06 204.3 ;
      RECT 29.42 204.18 29.62 204.3 ;
      RECT 29.78 202.68 29.98 202.8 ;
      RECT 31.22 202.92 31.42 203.04 ;
      RECT 30.5 203.222 30.7 203.342 ;
      RECT 30.5 200.702 30.7 200.822 ;
      RECT 29.06 200.942 29.26 201.062 ;
      RECT 31.94 200.942 32.14 201.062 ;
      RECT 30.14 201.42 30.34 201.54 ;
      RECT 30.86 201.66 31.06 201.78 ;
      RECT 31.58 201.66 31.78 201.78 ;
      RECT 32.3 201.66 32.5 201.78 ;
      RECT 28.7 201.66 28.9 201.78 ;
      RECT 29.42 201.66 29.62 201.78 ;
      RECT 29.78 200.16 29.98 200.28 ;
      RECT 31.22 200.4 31.42 200.52 ;
      RECT 30.5 198.182 30.7 198.302 ;
      RECT 31.94 198.422 32.14 198.542 ;
      RECT 29.06 198.422 29.26 198.542 ;
      RECT 30.14 198.9 30.34 199.02 ;
      RECT 32.3 199.14 32.5 199.26 ;
      RECT 31.58 199.14 31.78 199.26 ;
      RECT 30.86 199.14 31.06 199.26 ;
      RECT 29.42 199.14 29.62 199.26 ;
      RECT 28.7 199.14 28.9 199.26 ;
      RECT 28.7 196.62 28.9 196.74 ;
      RECT 29.42 196.62 29.62 196.74 ;
      RECT 30.14 196.62 30.34 196.74 ;
      RECT 30.86 196.62 31.06 196.74 ;
      RECT 32.3 196.62 32.5 196.74 ;
      RECT 31.22 197.64 31.42 197.76 ;
      RECT 29.78 197.88 29.98 198 ;
      RECT 29.78 195.36 29.98 195.48 ;
      RECT 31.94 195.662 32.14 195.782 ;
      RECT 30.5 195.902 30.7 196.022 ;
      RECT 29.06 195.902 29.26 196.022 ;
      RECT 31.58 196.38 31.78 196.5 ;
      RECT 31.58 193.86 31.78 193.98 ;
      RECT 29.42 193.86 29.62 193.98 ;
      RECT 28.7 194.1 28.9 194.22 ;
      RECT 30.14 194.1 30.34 194.22 ;
      RECT 30.86 194.1 31.06 194.22 ;
      RECT 32.3 194.1 32.5 194.22 ;
      RECT 31.94 194.402 32.14 194.522 ;
      RECT 30.5 194.642 30.7 194.762 ;
      RECT 29.06 194.642 29.26 194.762 ;
      RECT 31.22 195.12 31.42 195.24 ;
      RECT 29.78 192.84 29.98 192.96 ;
      RECT 31.22 192.84 31.42 192.96 ;
      RECT 31.94 193.142 32.14 193.262 ;
      RECT 29.06 193.142 29.26 193.262 ;
      RECT 30.5 193.382 30.7 193.502 ;
      RECT 30.86 191.34 31.06 191.46 ;
      RECT 29.42 191.34 29.62 191.46 ;
      RECT 30.14 191.58 30.34 191.7 ;
      RECT 31.58 191.58 31.78 191.7 ;
      RECT 32.3 191.58 32.5 191.7 ;
      RECT 28.7 191.58 28.9 191.7 ;
      RECT 31.94 191.882 32.14 192.002 ;
      RECT 29.06 191.882 29.26 192.002 ;
      RECT 30.5 192.122 30.7 192.242 ;
      RECT 31.22 190.08 31.42 190.2 ;
      RECT 29.06 220.17 29.26 220.29 ;
      RECT 30.5 220.17 30.7 220.29 ;
      RECT 31.94 220.17 32.14 220.29 ;
      RECT 31.94 218.91 32.14 219.03 ;
      RECT 30.5 218.91 30.7 219.03 ;
      RECT 29.06 218.91 29.26 219.03 ;
      RECT 28.7 219.54 28.9 219.66 ;
      RECT 29.42 219.54 29.62 219.66 ;
      RECT 30.14 219.54 30.34 219.66 ;
      RECT 30.86 219.54 31.06 219.66 ;
      RECT 31.58 219.54 31.78 219.66 ;
      RECT 32.3 219.54 32.5 219.66 ;
      RECT 31.94 217.65 32.14 217.77 ;
      RECT 30.5 217.65 30.7 217.77 ;
      RECT 29.06 217.65 29.26 217.77 ;
      RECT 28.7 218.28 28.9 218.4 ;
      RECT 29.42 218.28 29.62 218.4 ;
      RECT 30.14 218.28 30.34 218.4 ;
      RECT 30.86 218.28 31.06 218.4 ;
      RECT 31.58 218.28 31.78 218.4 ;
      RECT 32.3 218.28 32.5 218.4 ;
      RECT 32.3 215.76 32.5 215.88 ;
      RECT 31.58 215.76 31.78 215.88 ;
      RECT 30.86 215.76 31.06 215.88 ;
      RECT 30.14 215.76 30.34 215.88 ;
      RECT 29.42 215.76 29.62 215.88 ;
      RECT 28.7 215.76 28.9 215.88 ;
      RECT 29.06 216.39 29.26 216.51 ;
      RECT 30.5 216.39 30.7 216.51 ;
      RECT 31.94 216.39 32.14 216.51 ;
      RECT 32.3 217.02 32.5 217.14 ;
      RECT 31.58 217.02 31.78 217.14 ;
      RECT 30.86 217.02 31.06 217.14 ;
      RECT 30.14 217.02 30.34 217.14 ;
      RECT 29.42 217.02 29.62 217.14 ;
      RECT 28.7 217.02 28.9 217.14 ;
      RECT 28.7 214.5 28.9 214.62 ;
      RECT 29.42 214.5 29.62 214.62 ;
      RECT 30.14 214.5 30.34 214.62 ;
      RECT 30.86 214.5 31.06 214.62 ;
      RECT 31.58 214.5 31.78 214.62 ;
      RECT 32.3 214.5 32.5 214.62 ;
      RECT 31.94 215.13 32.14 215.25 ;
      RECT 30.5 215.13 30.7 215.25 ;
      RECT 29.06 215.13 29.26 215.25 ;
      RECT 32.3 213.24 32.5 213.36 ;
      RECT 31.58 213.24 31.78 213.36 ;
      RECT 30.86 213.24 31.06 213.36 ;
      RECT 30.14 213.24 30.34 213.36 ;
      RECT 29.42 213.24 29.62 213.36 ;
      RECT 28.7 213.24 28.9 213.36 ;
      RECT 31.94 213.87 32.14 213.99 ;
      RECT 30.5 213.87 30.7 213.99 ;
      RECT 29.06 213.87 29.26 213.99 ;
      RECT 28.7 211.98 28.9 212.1 ;
      RECT 29.42 211.98 29.62 212.1 ;
      RECT 30.14 211.98 30.34 212.1 ;
      RECT 30.86 211.98 31.06 212.1 ;
      RECT 31.58 211.98 31.78 212.1 ;
      RECT 32.3 211.98 32.5 212.1 ;
      RECT 31.94 212.61 32.14 212.73 ;
      RECT 30.5 212.61 30.7 212.73 ;
      RECT 29.06 212.61 29.26 212.73 ;
      RECT 32.3 210.72 32.5 210.84 ;
      RECT 31.58 210.72 31.78 210.84 ;
      RECT 30.86 210.72 31.06 210.84 ;
      RECT 30.14 210.72 30.34 210.84 ;
      RECT 29.42 210.72 29.62 210.84 ;
      RECT 28.7 210.72 28.9 210.84 ;
      RECT 31.94 211.35 32.14 211.47 ;
      RECT 30.5 211.35 30.7 211.47 ;
      RECT 29.06 211.35 29.26 211.47 ;
      RECT 28.7 209.46 28.9 209.58 ;
      RECT 29.42 209.46 29.62 209.58 ;
      RECT 30.14 209.46 30.34 209.58 ;
      RECT 30.86 209.46 31.06 209.58 ;
      RECT 31.58 209.46 31.78 209.58 ;
      RECT 32.3 209.46 32.5 209.58 ;
      RECT 29.06 210.09 29.26 210.21 ;
      RECT 30.5 210.09 30.7 210.21 ;
      RECT 31.94 210.09 32.14 210.21 ;
      RECT 31.22 207.72 31.42 207.84 ;
      RECT 29.78 207.96 29.98 208.08 ;
      RECT 30.5 208.262 30.7 208.382 ;
      RECT 31.94 208.502 32.14 208.622 ;
      RECT 29.06 208.502 29.26 208.622 ;
      RECT 30.14 206.46 30.34 206.58 ;
      RECT 32.3 206.46 32.5 206.58 ;
      RECT 28.7 206.7 28.9 206.82 ;
      RECT 29.42 206.7 29.62 206.82 ;
      RECT 30.86 206.7 31.06 206.82 ;
      RECT 31.58 206.7 31.78 206.82 ;
      RECT 29.78 205.2 29.98 205.32 ;
      RECT 31.22 205.44 31.42 205.56 ;
      RECT 30.5 205.742 30.7 205.862 ;
      RECT 31.94 205.982 32.14 206.102 ;
      RECT 29.06 205.982 29.26 206.102 ;
      RECT 29.06 203.462 29.26 203.582 ;
      RECT 31.94 203.462 32.14 203.582 ;
      RECT 28.7 203.94 28.9 204.06 ;
      RECT 30.14 203.94 30.34 204.06 ;
      RECT 31.58 203.94 31.78 204.06 ;
      RECT 28.7 234.66 28.9 234.78 ;
      RECT 29.42 234.66 29.62 234.78 ;
      RECT 30.14 234.66 30.34 234.78 ;
      RECT 30.86 234.66 31.06 234.78 ;
      RECT 31.58 234.66 31.78 234.78 ;
      RECT 32.3 234.66 32.5 234.78 ;
      RECT 28.7 232.14 28.9 232.26 ;
      RECT 29.42 232.14 29.62 232.26 ;
      RECT 30.14 232.14 30.34 232.26 ;
      RECT 30.86 232.14 31.06 232.26 ;
      RECT 31.58 232.14 31.78 232.26 ;
      RECT 32.3 232.14 32.5 232.26 ;
      RECT 29.06 232.77 29.26 232.89 ;
      RECT 30.5 232.77 30.7 232.89 ;
      RECT 31.94 232.77 32.14 232.89 ;
      RECT 32.3 233.4 32.5 233.52 ;
      RECT 31.58 233.4 31.78 233.52 ;
      RECT 30.86 233.4 31.06 233.52 ;
      RECT 30.14 233.4 30.34 233.52 ;
      RECT 29.42 233.4 29.62 233.52 ;
      RECT 28.7 233.4 28.9 233.52 ;
      RECT 28.7 230.88 28.9 231 ;
      RECT 29.42 230.88 29.62 231 ;
      RECT 30.14 230.88 30.34 231 ;
      RECT 30.86 230.88 31.06 231 ;
      RECT 31.58 230.88 31.78 231 ;
      RECT 32.3 230.88 32.5 231 ;
      RECT 29.06 231.51 29.26 231.63 ;
      RECT 30.5 231.51 30.7 231.63 ;
      RECT 31.94 231.51 32.14 231.63 ;
      RECT 32.3 229.62 32.5 229.74 ;
      RECT 31.58 229.62 31.78 229.74 ;
      RECT 30.86 229.62 31.06 229.74 ;
      RECT 30.14 229.62 30.34 229.74 ;
      RECT 29.42 229.62 29.62 229.74 ;
      RECT 28.7 229.62 28.9 229.74 ;
      RECT 29.06 230.25 29.26 230.37 ;
      RECT 30.5 230.25 30.7 230.37 ;
      RECT 31.94 230.25 32.14 230.37 ;
      RECT 32.3 228.36 32.5 228.48 ;
      RECT 31.58 228.36 31.78 228.48 ;
      RECT 30.86 228.36 31.06 228.48 ;
      RECT 30.14 228.36 30.34 228.48 ;
      RECT 29.42 228.36 29.62 228.48 ;
      RECT 28.7 228.36 28.9 228.48 ;
      RECT 31.94 228.99 32.14 229.11 ;
      RECT 30.5 228.99 30.7 229.11 ;
      RECT 29.06 228.99 29.26 229.11 ;
      RECT 32.3 227.1 32.5 227.22 ;
      RECT 31.58 227.1 31.78 227.22 ;
      RECT 30.86 227.1 31.06 227.22 ;
      RECT 30.14 227.1 30.34 227.22 ;
      RECT 29.42 227.1 29.62 227.22 ;
      RECT 28.7 227.1 28.9 227.22 ;
      RECT 31.94 227.73 32.14 227.85 ;
      RECT 30.5 227.73 30.7 227.85 ;
      RECT 29.06 227.73 29.26 227.85 ;
      RECT 32.3 225.84 32.5 225.96 ;
      RECT 31.58 225.84 31.78 225.96 ;
      RECT 30.86 225.84 31.06 225.96 ;
      RECT 30.14 225.84 30.34 225.96 ;
      RECT 29.42 225.84 29.62 225.96 ;
      RECT 28.7 225.84 28.9 225.96 ;
      RECT 31.94 226.47 32.14 226.59 ;
      RECT 30.5 226.47 30.7 226.59 ;
      RECT 29.06 226.47 29.26 226.59 ;
      RECT 31.94 223.95 32.14 224.07 ;
      RECT 30.5 223.95 30.7 224.07 ;
      RECT 29.06 223.95 29.26 224.07 ;
      RECT 32.3 224.58 32.5 224.7 ;
      RECT 31.58 224.58 31.78 224.7 ;
      RECT 30.86 224.58 31.06 224.7 ;
      RECT 30.14 224.58 30.34 224.7 ;
      RECT 29.42 224.58 29.62 224.7 ;
      RECT 28.7 224.58 28.9 224.7 ;
      RECT 31.94 225.21 32.14 225.33 ;
      RECT 30.5 225.21 30.7 225.33 ;
      RECT 29.06 225.21 29.26 225.33 ;
      RECT 31.94 222.69 32.14 222.81 ;
      RECT 30.5 222.69 30.7 222.81 ;
      RECT 29.06 222.69 29.26 222.81 ;
      RECT 32.3 223.32 32.5 223.44 ;
      RECT 31.58 223.32 31.78 223.44 ;
      RECT 30.86 223.32 31.06 223.44 ;
      RECT 30.14 223.32 30.34 223.44 ;
      RECT 29.42 223.32 29.62 223.44 ;
      RECT 28.7 223.32 28.9 223.44 ;
      RECT 29.06 221.43 29.26 221.55 ;
      RECT 30.5 221.43 30.7 221.55 ;
      RECT 31.94 221.43 32.14 221.55 ;
      RECT 32.3 222.06 32.5 222.18 ;
      RECT 31.58 222.06 31.78 222.18 ;
      RECT 30.86 222.06 31.06 222.18 ;
      RECT 30.14 222.06 30.34 222.18 ;
      RECT 29.42 222.06 29.62 222.18 ;
      RECT 28.7 222.06 28.9 222.18 ;
      RECT 32.3 220.8 32.5 220.92 ;
      RECT 31.58 220.8 31.78 220.92 ;
      RECT 30.86 220.8 31.06 220.92 ;
      RECT 30.14 220.8 30.34 220.92 ;
      RECT 29.42 220.8 29.62 220.92 ;
      RECT 28.7 220.8 28.9 220.92 ;
      RECT 28.7 249.78 28.9 249.9 ;
      RECT 29.42 249.78 29.62 249.9 ;
      RECT 30.14 249.78 30.34 249.9 ;
      RECT 30.86 249.78 31.06 249.9 ;
      RECT 31.58 249.78 31.78 249.9 ;
      RECT 32.3 249.78 32.5 249.9 ;
      RECT 28.7 247.26 28.9 247.38 ;
      RECT 29.42 247.26 29.62 247.38 ;
      RECT 30.14 247.26 30.34 247.38 ;
      RECT 30.86 247.26 31.06 247.38 ;
      RECT 31.58 247.26 31.78 247.38 ;
      RECT 32.3 247.26 32.5 247.38 ;
      RECT 29.06 247.89 29.26 248.01 ;
      RECT 30.5 247.89 30.7 248.01 ;
      RECT 31.94 247.89 32.14 248.01 ;
      RECT 29.06 246.63 29.26 246.75 ;
      RECT 30.5 246.63 30.7 246.75 ;
      RECT 31.94 246.63 32.14 246.75 ;
      RECT 32.3 246 32.5 246.12 ;
      RECT 31.58 246 31.78 246.12 ;
      RECT 30.86 246 31.06 246.12 ;
      RECT 30.14 246 30.34 246.12 ;
      RECT 29.42 246 29.62 246.12 ;
      RECT 28.7 246 28.9 246.12 ;
      RECT 32.3 244.74 32.5 244.86 ;
      RECT 31.58 244.74 31.78 244.86 ;
      RECT 30.86 244.74 31.06 244.86 ;
      RECT 30.14 244.74 30.34 244.86 ;
      RECT 29.42 244.74 29.62 244.86 ;
      RECT 28.7 244.74 28.9 244.86 ;
      RECT 31.94 245.37 32.14 245.49 ;
      RECT 30.5 245.37 30.7 245.49 ;
      RECT 29.06 245.37 29.26 245.49 ;
      RECT 28.7 243.48 28.9 243.6 ;
      RECT 29.42 243.48 29.62 243.6 ;
      RECT 30.14 243.48 30.34 243.6 ;
      RECT 30.86 243.48 31.06 243.6 ;
      RECT 31.58 243.48 31.78 243.6 ;
      RECT 32.3 243.48 32.5 243.6 ;
      RECT 29.06 244.11 29.26 244.23 ;
      RECT 30.5 244.11 30.7 244.23 ;
      RECT 31.94 244.11 32.14 244.23 ;
      RECT 28.7 242.22 28.9 242.34 ;
      RECT 29.42 242.22 29.62 242.34 ;
      RECT 30.14 242.22 30.34 242.34 ;
      RECT 30.86 242.22 31.06 242.34 ;
      RECT 31.58 242.22 31.78 242.34 ;
      RECT 32.3 242.22 32.5 242.34 ;
      RECT 29.06 242.85 29.26 242.97 ;
      RECT 30.5 242.85 30.7 242.97 ;
      RECT 31.94 242.85 32.14 242.97 ;
      RECT 29.06 240.33 29.26 240.45 ;
      RECT 30.5 240.33 30.7 240.45 ;
      RECT 31.94 240.33 32.14 240.45 ;
      RECT 32.3 240.96 32.5 241.08 ;
      RECT 31.58 240.96 31.78 241.08 ;
      RECT 30.86 240.96 31.06 241.08 ;
      RECT 30.14 240.96 30.34 241.08 ;
      RECT 29.42 240.96 29.62 241.08 ;
      RECT 28.7 240.96 28.9 241.08 ;
      RECT 31.94 241.59 32.14 241.71 ;
      RECT 30.5 241.59 30.7 241.71 ;
      RECT 29.06 241.59 29.26 241.71 ;
      RECT 29.06 239.07 29.26 239.19 ;
      RECT 30.5 239.07 30.7 239.19 ;
      RECT 31.94 239.07 32.14 239.19 ;
      RECT 28.7 239.7 28.9 239.82 ;
      RECT 29.42 239.7 29.62 239.82 ;
      RECT 30.14 239.7 30.34 239.82 ;
      RECT 30.86 239.7 31.06 239.82 ;
      RECT 31.58 239.7 31.78 239.82 ;
      RECT 32.3 239.7 32.5 239.82 ;
      RECT 31.94 237.81 32.14 237.93 ;
      RECT 30.5 237.81 30.7 237.93 ;
      RECT 29.06 237.81 29.26 237.93 ;
      RECT 28.7 238.44 28.9 238.56 ;
      RECT 29.42 238.44 29.62 238.56 ;
      RECT 30.14 238.44 30.34 238.56 ;
      RECT 30.86 238.44 31.06 238.56 ;
      RECT 31.58 238.44 31.78 238.56 ;
      RECT 32.3 238.44 32.5 238.56 ;
      RECT 29.06 236.55 29.26 236.67 ;
      RECT 30.5 236.55 30.7 236.67 ;
      RECT 31.94 236.55 32.14 236.67 ;
      RECT 31.58 237.18 31.78 237.3 ;
      RECT 30.86 237.18 31.06 237.3 ;
      RECT 30.14 237.18 30.34 237.3 ;
      RECT 29.42 237.18 29.62 237.3 ;
      RECT 28.7 237.18 28.9 237.3 ;
      RECT 32.3 237.18 32.5 237.3 ;
      RECT 29.06 235.29 29.26 235.41 ;
      RECT 30.5 235.29 30.7 235.41 ;
      RECT 31.94 235.29 32.14 235.41 ;
      RECT 28.7 235.92 28.9 236.04 ;
      RECT 29.42 235.92 29.62 236.04 ;
      RECT 30.14 235.92 30.34 236.04 ;
      RECT 30.86 235.92 31.06 236.04 ;
      RECT 31.58 235.92 31.78 236.04 ;
      RECT 32.3 235.92 32.5 236.04 ;
      RECT 31.94 234.03 32.14 234.15 ;
      RECT 30.5 234.03 30.7 234.15 ;
      RECT 29.06 234.03 29.26 234.15 ;
      RECT 28.7 262.38 28.9 262.5 ;
      RECT 29.42 262.38 29.62 262.5 ;
      RECT 30.14 262.38 30.34 262.5 ;
      RECT 30.86 262.38 31.06 262.5 ;
      RECT 31.58 262.38 31.78 262.5 ;
      RECT 32.3 262.38 32.5 262.5 ;
      RECT 31.94 263.01 32.14 263.13 ;
      RECT 30.5 263.01 30.7 263.13 ;
      RECT 29.06 263.01 29.26 263.13 ;
      RECT 32.3 261.12 32.5 261.24 ;
      RECT 30.86 261.12 31.06 261.24 ;
      RECT 31.58 261.12 31.78 261.24 ;
      RECT 28.7 261.12 28.9 261.24 ;
      RECT 29.42 261.12 29.62 261.24 ;
      RECT 30.14 261.12 30.34 261.24 ;
      RECT 29.06 261.75 29.26 261.87 ;
      RECT 30.5 261.75 30.7 261.87 ;
      RECT 31.94 261.75 32.14 261.87 ;
      RECT 28.7 259.86 28.9 259.98 ;
      RECT 29.42 259.86 29.62 259.98 ;
      RECT 30.14 259.86 30.34 259.98 ;
      RECT 30.86 259.86 31.06 259.98 ;
      RECT 31.58 259.86 31.78 259.98 ;
      RECT 32.3 259.86 32.5 259.98 ;
      RECT 30.5 260.49 30.7 260.61 ;
      RECT 31.94 260.49 32.14 260.61 ;
      RECT 29.06 260.49 29.26 260.61 ;
      RECT 28.7 258.6 28.9 258.72 ;
      RECT 29.42 258.6 29.62 258.72 ;
      RECT 30.14 258.6 30.34 258.72 ;
      RECT 30.86 258.6 31.06 258.72 ;
      RECT 31.58 258.6 31.78 258.72 ;
      RECT 32.3 258.6 32.5 258.72 ;
      RECT 29.06 259.23 29.26 259.35 ;
      RECT 30.5 259.23 30.7 259.35 ;
      RECT 31.94 259.23 32.14 259.35 ;
      RECT 29.06 256.71 29.26 256.83 ;
      RECT 30.5 256.71 30.7 256.83 ;
      RECT 31.94 256.71 32.14 256.83 ;
      RECT 28.7 257.34 28.9 257.46 ;
      RECT 29.42 257.34 29.62 257.46 ;
      RECT 30.14 257.34 30.34 257.46 ;
      RECT 30.86 257.34 31.06 257.46 ;
      RECT 31.58 257.34 31.78 257.46 ;
      RECT 32.3 257.34 32.5 257.46 ;
      RECT 29.06 257.97 29.26 258.09 ;
      RECT 30.5 257.97 30.7 258.09 ;
      RECT 31.94 257.97 32.14 258.09 ;
      RECT 29.06 255.45 29.26 255.57 ;
      RECT 31.94 255.45 32.14 255.57 ;
      RECT 30.5 255.45 30.7 255.57 ;
      RECT 28.7 256.08 28.9 256.2 ;
      RECT 29.42 256.08 29.62 256.2 ;
      RECT 30.14 256.08 30.34 256.2 ;
      RECT 30.86 256.08 31.06 256.2 ;
      RECT 31.58 256.08 31.78 256.2 ;
      RECT 32.3 256.08 32.5 256.2 ;
      RECT 29.06 254.19 29.26 254.31 ;
      RECT 30.5 254.19 30.7 254.31 ;
      RECT 31.94 254.19 32.14 254.31 ;
      RECT 28.7 254.82 28.9 254.94 ;
      RECT 29.42 254.82 29.62 254.94 ;
      RECT 30.14 254.82 30.34 254.94 ;
      RECT 30.86 254.82 31.06 254.94 ;
      RECT 31.58 254.82 31.78 254.94 ;
      RECT 32.3 254.82 32.5 254.94 ;
      RECT 30.5 252.93 30.7 253.05 ;
      RECT 31.94 252.93 32.14 253.05 ;
      RECT 29.06 252.93 29.26 253.05 ;
      RECT 28.7 253.56 28.9 253.68 ;
      RECT 29.42 253.56 29.62 253.68 ;
      RECT 30.14 253.56 30.34 253.68 ;
      RECT 30.86 253.56 31.06 253.68 ;
      RECT 31.58 253.56 31.78 253.68 ;
      RECT 32.3 253.56 32.5 253.68 ;
      RECT 29.06 251.67 29.26 251.79 ;
      RECT 30.5 251.67 30.7 251.79 ;
      RECT 31.94 251.67 32.14 251.79 ;
      RECT 28.7 252.3 28.9 252.42 ;
      RECT 29.42 252.3 29.62 252.42 ;
      RECT 30.14 252.3 30.34 252.42 ;
      RECT 30.86 252.3 31.06 252.42 ;
      RECT 31.58 252.3 31.78 252.42 ;
      RECT 32.3 252.3 32.5 252.42 ;
      RECT 29.06 250.41 29.26 250.53 ;
      RECT 30.5 250.41 30.7 250.53 ;
      RECT 31.94 250.41 32.14 250.53 ;
      RECT 28.7 251.04 28.9 251.16 ;
      RECT 29.42 251.04 29.62 251.16 ;
      RECT 30.14 251.04 30.34 251.16 ;
      RECT 30.86 251.04 31.06 251.16 ;
      RECT 31.58 251.04 31.78 251.16 ;
      RECT 32.3 251.04 32.5 251.16 ;
      RECT 28.7 248.52 28.9 248.64 ;
      RECT 29.42 248.52 29.62 248.64 ;
      RECT 30.14 248.52 30.34 248.64 ;
      RECT 30.86 248.52 31.06 248.64 ;
      RECT 31.58 248.52 31.78 248.64 ;
      RECT 32.3 248.52 32.5 248.64 ;
      RECT 29.06 249.15 29.26 249.27 ;
      RECT 30.5 249.15 30.7 249.27 ;
      RECT 31.94 249.15 32.14 249.27 ;
      RECT 30.86 268.68 31.06 268.8 ;
      RECT 31.58 268.68 31.78 268.8 ;
      RECT 32.3 268.68 32.5 268.8 ;
      RECT 29.06 266.79 29.26 266.91 ;
      RECT 30.5 266.79 30.7 266.91 ;
      RECT 31.94 266.79 32.14 266.91 ;
      RECT 28.7 267.42 28.9 267.54 ;
      RECT 29.42 267.42 29.62 267.54 ;
      RECT 30.14 267.42 30.34 267.54 ;
      RECT 30.86 267.42 31.06 267.54 ;
      RECT 31.58 267.42 31.78 267.54 ;
      RECT 32.3 267.42 32.5 267.54 ;
      RECT 28.7 264.9 28.9 265.02 ;
      RECT 29.42 264.9 29.62 265.02 ;
      RECT 30.14 264.9 30.34 265.02 ;
      RECT 30.86 264.9 31.06 265.02 ;
      RECT 31.58 264.9 31.78 265.02 ;
      RECT 32.3 264.9 32.5 265.02 ;
      RECT 29.06 265.53 29.26 265.65 ;
      RECT 30.5 265.53 30.7 265.65 ;
      RECT 31.94 265.53 32.14 265.65 ;
      RECT 28.7 266.16 28.9 266.28 ;
      RECT 29.42 266.16 29.62 266.28 ;
      RECT 30.14 266.16 30.34 266.28 ;
      RECT 30.86 266.16 31.06 266.28 ;
      RECT 31.58 266.16 31.78 266.28 ;
      RECT 32.3 266.16 32.5 266.28 ;
      RECT 30.86 263.64 31.06 263.76 ;
      RECT 31.58 263.64 31.78 263.76 ;
      RECT 32.3 263.64 32.5 263.76 ;
      RECT 28.7 263.64 28.9 263.76 ;
      RECT 29.42 263.64 29.62 263.76 ;
      RECT 30.14 263.64 30.34 263.76 ;
      RECT 29.06 264.27 29.26 264.39 ;
      RECT 30.5 264.27 30.7 264.39 ;
      RECT 31.94 264.27 32.14 264.39 ;
      RECT 30.86 273.72 31.06 273.84 ;
      RECT 30.14 273.72 30.34 273.84 ;
      RECT 29.42 273.72 29.62 273.84 ;
      RECT 28.7 273.72 28.9 273.84 ;
      RECT 31.94 273.09 32.14 273.21 ;
      RECT 30.5 273.09 30.7 273.21 ;
      RECT 29.06 273.09 29.26 273.21 ;
      RECT 32.3 272.46 32.5 272.58 ;
      RECT 31.58 272.46 31.78 272.58 ;
      RECT 30.86 272.46 31.06 272.58 ;
      RECT 30.14 272.46 30.34 272.58 ;
      RECT 29.42 272.46 29.62 272.58 ;
      RECT 28.7 272.46 28.9 272.58 ;
      RECT 31.94 271.83 32.14 271.95 ;
      RECT 30.5 271.83 30.7 271.95 ;
      RECT 29.06 271.83 29.26 271.95 ;
      RECT 29.06 270.57 29.26 270.69 ;
      RECT 30.5 270.57 30.7 270.69 ;
      RECT 31.94 270.57 32.14 270.69 ;
      RECT 32.3 271.2 32.5 271.32 ;
      RECT 28.7 271.2 28.9 271.32 ;
      RECT 29.42 271.2 29.62 271.32 ;
      RECT 30.14 271.2 30.34 271.32 ;
      RECT 30.86 271.2 31.06 271.32 ;
      RECT 31.58 271.2 31.78 271.32 ;
      RECT 29.06 269.31 29.26 269.43 ;
      RECT 30.5 269.31 30.7 269.43 ;
      RECT 31.94 269.31 32.14 269.43 ;
      RECT 28.7 269.94 28.9 270.06 ;
      RECT 29.42 269.94 29.62 270.06 ;
      RECT 30.14 269.94 30.34 270.06 ;
      RECT 30.86 269.94 31.06 270.06 ;
      RECT 31.58 269.94 31.78 270.06 ;
      RECT 32.3 269.94 32.5 270.06 ;
      RECT 29.06 268.05 29.26 268.17 ;
      RECT 30.5 268.05 30.7 268.17 ;
      RECT 31.94 268.05 32.14 268.17 ;
      RECT 28.7 268.68 28.9 268.8 ;
      RECT 29.42 268.68 29.62 268.8 ;
      RECT 30.14 268.68 30.34 268.8 ;
      RECT 30.14 305.967 30.34 306.087 ;
      RECT 29.42 305.967 29.62 306.087 ;
      RECT 28.7 305.967 28.9 306.087 ;
      RECT 31.22 305.498 31.42 305.618 ;
      RECT 29.78 305.498 29.98 305.618 ;
      RECT 32.3 283.087 32.5 283.207 ;
      RECT 31.58 283.087 31.78 283.207 ;
      RECT 30.86 283.087 31.06 283.207 ;
      RECT 30.14 283.087 30.34 283.207 ;
      RECT 29.42 283.087 29.62 283.207 ;
      RECT 28.7 283.087 28.9 283.207 ;
      RECT 32.3 278.76 32.5 278.88 ;
      RECT 31.58 278.76 31.78 278.88 ;
      RECT 30.86 278.76 31.06 278.88 ;
      RECT 30.14 278.76 30.34 278.88 ;
      RECT 29.42 278.76 29.62 278.88 ;
      RECT 28.7 278.76 28.9 278.88 ;
      RECT 31.94 278.13 32.14 278.25 ;
      RECT 30.5 278.13 30.7 278.25 ;
      RECT 29.06 278.13 29.26 278.25 ;
      RECT 31.58 277.5 31.78 277.62 ;
      RECT 30.86 277.5 31.06 277.62 ;
      RECT 30.14 277.5 30.34 277.62 ;
      RECT 29.42 277.5 29.62 277.62 ;
      RECT 28.7 277.5 28.9 277.62 ;
      RECT 32.3 277.5 32.5 277.62 ;
      RECT 31.94 276.87 32.14 276.99 ;
      RECT 30.5 276.87 30.7 276.99 ;
      RECT 29.06 276.87 29.26 276.99 ;
      RECT 32.3 276.24 32.5 276.36 ;
      RECT 31.58 276.24 31.78 276.36 ;
      RECT 30.86 276.24 31.06 276.36 ;
      RECT 30.14 276.24 30.34 276.36 ;
      RECT 29.42 276.24 29.62 276.36 ;
      RECT 28.7 276.24 28.9 276.36 ;
      RECT 31.94 275.61 32.14 275.73 ;
      RECT 30.5 275.61 30.7 275.73 ;
      RECT 29.06 275.61 29.26 275.73 ;
      RECT 32.3 274.98 32.5 275.1 ;
      RECT 31.58 274.98 31.78 275.1 ;
      RECT 30.86 274.98 31.06 275.1 ;
      RECT 30.14 274.98 30.34 275.1 ;
      RECT 29.42 274.98 29.62 275.1 ;
      RECT 28.7 274.98 28.9 275.1 ;
      RECT 31.94 274.35 32.14 274.47 ;
      RECT 30.5 274.35 30.7 274.47 ;
      RECT 29.06 274.35 29.26 274.47 ;
      RECT 32.3 273.72 32.5 273.84 ;
      RECT 31.58 273.72 31.78 273.84 ;
      RECT 36.62 123.3 36.82 123.42 ;
      RECT 35.54 122.28 35.74 122.4 ;
      RECT 34.46 121.498 34.66 121.618 ;
      RECT 35.18 121.498 35.38 121.618 ;
      RECT 35.9 121.498 36.1 121.618 ;
      RECT 36.62 121.498 36.82 121.618 ;
      RECT 34.46 121.02 34.66 121.14 ;
      RECT 35.9 121.02 36.1 121.14 ;
      RECT 36.62 120.78 36.82 120.9 ;
      RECT 35.18 120.78 35.38 120.9 ;
      RECT 35.54 119.76 35.74 119.88 ;
      RECT 34.46 118.978 34.66 119.098 ;
      RECT 35.18 118.978 35.38 119.098 ;
      RECT 35.9 118.978 36.1 119.098 ;
      RECT 36.62 118.978 36.82 119.098 ;
      RECT 36.62 118.5 36.82 118.62 ;
      RECT 34.46 118.5 34.66 118.62 ;
      RECT 35.9 118.26 36.1 118.38 ;
      RECT 35.18 118.26 35.38 118.38 ;
      RECT 31.22 348.339 31.42 348.459 ;
      RECT 29.78 348.339 29.98 348.459 ;
      RECT 32.3 325.9425 32.5 326.0625 ;
      RECT 31.58 325.9425 31.78 326.0625 ;
      RECT 30.86 325.9425 31.06 326.0625 ;
      RECT 30.14 325.9425 30.34 326.0625 ;
      RECT 29.42 325.9425 29.62 326.0625 ;
      RECT 28.7 325.9425 28.9 326.0625 ;
      RECT 31.22 323.3835 31.42 323.5035 ;
      RECT 29.78 323.3835 29.98 323.5035 ;
      RECT 32.3 305.967 32.5 306.087 ;
      RECT 31.58 305.967 31.78 306.087 ;
      RECT 30.86 305.967 31.06 306.087 ;
      RECT 36.62 140.94 36.82 141.06 ;
      RECT 35.54 139.68 35.74 139.8 ;
      RECT 34.46 139.138 34.66 139.258 ;
      RECT 35.18 139.138 35.38 139.258 ;
      RECT 35.9 139.138 36.1 139.258 ;
      RECT 36.62 139.138 36.82 139.258 ;
      RECT 36.62 138.66 36.82 138.78 ;
      RECT 35.18 138.66 35.38 138.78 ;
      RECT 35.9 138.42 36.1 138.54 ;
      RECT 34.46 138.42 34.66 138.54 ;
      RECT 35.54 137.4 35.74 137.52 ;
      RECT 34.46 136.618 34.66 136.738 ;
      RECT 35.18 136.618 35.38 136.738 ;
      RECT 35.9 136.618 36.1 136.738 ;
      RECT 36.62 136.618 36.82 136.738 ;
      RECT 34.46 136.14 34.66 136.26 ;
      RECT 35.18 136.14 35.38 136.26 ;
      RECT 36.62 136.14 36.82 136.26 ;
      RECT 35.9 135.9 36.1 136.02 ;
      RECT 35.54 134.64 35.74 134.76 ;
      RECT 34.46 134.098 34.66 134.218 ;
      RECT 35.18 134.098 35.38 134.218 ;
      RECT 35.9 134.098 36.1 134.218 ;
      RECT 36.62 134.098 36.82 134.218 ;
      RECT 35.9 133.62 36.1 133.74 ;
      RECT 36.62 133.38 36.82 133.5 ;
      RECT 35.18 133.38 35.38 133.5 ;
      RECT 34.46 133.38 34.66 133.5 ;
      RECT 35.54 132.36 35.74 132.48 ;
      RECT 34.46 131.578 34.66 131.698 ;
      RECT 35.18 131.578 35.38 131.698 ;
      RECT 35.9 131.578 36.1 131.698 ;
      RECT 36.62 131.578 36.82 131.698 ;
      RECT 36.62 131.1 36.82 131.22 ;
      RECT 35.18 131.1 35.38 131.22 ;
      RECT 34.46 130.86 34.66 130.98 ;
      RECT 35.9 130.86 36.1 130.98 ;
      RECT 35.54 129.84 35.74 129.96 ;
      RECT 34.46 129.058 34.66 129.178 ;
      RECT 35.18 129.058 35.38 129.178 ;
      RECT 35.9 129.058 36.1 129.178 ;
      RECT 36.62 129.058 36.82 129.178 ;
      RECT 36.62 128.58 36.82 128.7 ;
      RECT 35.18 128.58 35.38 128.7 ;
      RECT 35.9 128.34 36.1 128.46 ;
      RECT 34.46 128.34 34.66 128.46 ;
      RECT 35.54 127.32 35.74 127.44 ;
      RECT 34.46 126.538 34.66 126.658 ;
      RECT 35.18 126.538 35.38 126.658 ;
      RECT 35.9 126.538 36.1 126.658 ;
      RECT 36.62 126.538 36.82 126.658 ;
      RECT 35.18 126.06 35.38 126.18 ;
      RECT 35.9 126.06 36.1 126.18 ;
      RECT 36.62 126.06 36.82 126.18 ;
      RECT 34.46 125.82 34.66 125.94 ;
      RECT 35.54 124.8 35.74 124.92 ;
      RECT 34.46 124.018 34.66 124.138 ;
      RECT 35.18 124.018 35.38 124.138 ;
      RECT 35.9 124.018 36.1 124.138 ;
      RECT 36.62 124.018 36.82 124.138 ;
      RECT 35.18 123.54 35.38 123.66 ;
      RECT 35.9 123.54 36.1 123.66 ;
      RECT 34.46 123.3 34.66 123.42 ;
      RECT 35.9 140.94 36.1 141.06 ;
      RECT 34.46 141.18 34.66 141.3 ;
      RECT 35.9 158.82 36.1 158.94 ;
      RECT 35.18 158.82 35.38 158.94 ;
      RECT 34.46 158.82 34.66 158.94 ;
      RECT 35.54 157.56 35.74 157.68 ;
      RECT 34.82 158.038 35.02 158.158 ;
      RECT 36.26 158.278 36.46 158.398 ;
      RECT 35.9 156.06 36.1 156.18 ;
      RECT 36.62 156.06 36.82 156.18 ;
      RECT 35.18 156.3 35.38 156.42 ;
      RECT 34.46 156.3 34.66 156.42 ;
      RECT 34.82 156.842 35.02 156.962 ;
      RECT 36.26 156.842 36.46 156.962 ;
      RECT 35.54 155.04 35.74 155.16 ;
      RECT 35.18 153.54 35.38 153.66 ;
      RECT 36.62 153.54 36.82 153.66 ;
      RECT 34.46 153.78 34.66 153.9 ;
      RECT 35.9 153.78 36.1 153.9 ;
      RECT 35.54 152.28 35.74 152.4 ;
      RECT 34.46 151.02 34.66 151.14 ;
      RECT 35.9 151.02 36.1 151.14 ;
      RECT 35.18 151.26 35.38 151.38 ;
      RECT 36.62 151.26 36.82 151.38 ;
      RECT 35.54 150 35.74 150.12 ;
      RECT 35.18 148.5 35.38 148.62 ;
      RECT 35.9 148.5 36.1 148.62 ;
      RECT 36.62 148.74 36.82 148.86 ;
      RECT 34.46 148.74 34.66 148.86 ;
      RECT 35.54 144.96 35.74 145.08 ;
      RECT 36.62 145.98 36.82 146.1 ;
      RECT 35.9 145.98 36.1 146.1 ;
      RECT 35.18 145.98 35.38 146.1 ;
      RECT 34.46 145.98 34.66 146.1 ;
      RECT 35.9 143.46 36.1 143.58 ;
      RECT 34.46 143.46 34.66 143.58 ;
      RECT 35.18 143.7 35.38 143.82 ;
      RECT 36.62 143.7 36.82 143.82 ;
      RECT 35.54 142.44 35.74 142.56 ;
      RECT 35.18 141.18 35.38 141.3 ;
      RECT 35.54 177.72 35.74 177.84 ;
      RECT 35.18 178.74 35.38 178.86 ;
      RECT 34.46 176.46 34.66 176.58 ;
      RECT 35.18 176.46 35.38 176.58 ;
      RECT 35.9 176.46 36.1 176.58 ;
      RECT 36.62 176.46 36.82 176.58 ;
      RECT 35.54 175.2 35.74 175.32 ;
      RECT 35.9 173.7 36.1 173.82 ;
      RECT 36.62 173.7 36.82 173.82 ;
      RECT 34.46 173.94 34.66 174.06 ;
      RECT 35.18 173.94 35.38 174.06 ;
      RECT 35.54 172.68 35.74 172.8 ;
      RECT 36.62 171.18 36.82 171.3 ;
      RECT 35.18 171.18 35.38 171.3 ;
      RECT 34.46 171.18 34.66 171.3 ;
      RECT 35.9 171.42 36.1 171.54 ;
      RECT 35.54 169.92 35.74 170.04 ;
      RECT 36.62 168.66 36.82 168.78 ;
      RECT 35.9 168.66 36.1 168.78 ;
      RECT 34.46 168.9 34.66 169.02 ;
      RECT 35.18 168.9 35.38 169.02 ;
      RECT 35.54 167.64 35.74 167.76 ;
      RECT 36.62 166.14 36.82 166.26 ;
      RECT 34.46 166.38 34.66 166.5 ;
      RECT 35.18 166.38 35.38 166.5 ;
      RECT 35.9 166.38 36.1 166.5 ;
      RECT 34.46 163.86 34.66 163.98 ;
      RECT 35.9 163.86 36.1 163.98 ;
      RECT 36.62 163.86 36.82 163.98 ;
      RECT 35.54 165.12 35.74 165.24 ;
      RECT 35.54 162.6 35.74 162.72 ;
      RECT 35.18 163.62 35.38 163.74 ;
      RECT 36.62 161.1 36.82 161.22 ;
      RECT 35.9 161.1 36.1 161.22 ;
      RECT 35.18 161.1 35.38 161.22 ;
      RECT 34.46 161.1 34.66 161.22 ;
      RECT 35.54 160.08 35.74 160.2 ;
      RECT 36.62 158.82 36.82 158.94 ;
      RECT 36.62 186.3 36.82 186.42 ;
      RECT 35.18 186.3 35.38 186.42 ;
      RECT 35.9 186.54 36.1 186.66 ;
      RECT 34.46 186.54 34.66 186.66 ;
      RECT 35.54 185.28 35.74 185.4 ;
      RECT 34.46 183.78 34.66 183.9 ;
      RECT 36.62 183.78 36.82 183.9 ;
      RECT 35.18 184.02 35.38 184.14 ;
      RECT 35.9 184.02 36.1 184.14 ;
      RECT 35.54 182.76 35.74 182.88 ;
      RECT 35.54 180.24 35.74 180.36 ;
      RECT 35.18 181.26 35.38 181.38 ;
      RECT 35.9 181.26 36.1 181.38 ;
      RECT 36.62 181.5 36.82 181.62 ;
      RECT 34.46 181.5 34.66 181.62 ;
      RECT 36.62 178.98 36.82 179.1 ;
      RECT 35.9 178.98 36.1 179.1 ;
      RECT 34.46 178.98 34.66 179.1 ;
      RECT 35.54 187.8 35.74 187.92 ;
      RECT 34.46 196.38 34.66 196.5 ;
      RECT 35.9 193.86 36.1 193.98 ;
      RECT 34.46 193.86 34.66 193.98 ;
      RECT 35.18 194.1 35.38 194.22 ;
      RECT 36.62 194.1 36.82 194.22 ;
      RECT 36.26 194.402 36.46 194.522 ;
      RECT 34.82 194.642 35.02 194.762 ;
      RECT 35.54 192.6 35.74 192.72 ;
      RECT 36.26 193.142 36.46 193.262 ;
      RECT 34.82 193.382 35.02 193.502 ;
      RECT 36.62 191.34 36.82 191.46 ;
      RECT 35.18 191.34 35.38 191.46 ;
      RECT 34.46 191.34 34.66 191.46 ;
      RECT 35.9 191.58 36.1 191.7 ;
      RECT 36.26 191.882 36.46 192.002 ;
      RECT 34.82 192.122 35.02 192.242 ;
      RECT 35.54 190.32 35.74 190.44 ;
      RECT 36.26 190.622 36.46 190.742 ;
      RECT 34.82 190.862 35.02 190.982 ;
      RECT 35.9 188.82 36.1 188.94 ;
      RECT 36.62 189.06 36.82 189.18 ;
      RECT 35.18 189.06 35.38 189.18 ;
      RECT 34.46 189.06 34.66 189.18 ;
      RECT 201.14 323.3835 201.34 323.5035 ;
      RECT 200.78 306.041 200.98 306.161 ;
      RECT 200.06 306.041 200.26 306.161 ;
      RECT 199.34 306.041 199.54 306.161 ;
      RECT 198.62 306.041 198.82 306.161 ;
      RECT 201.14 348.339 201.34 348.459 ;
      RECT 188.9 282.3 189.1 282.42 ;
      RECT 192.14 285.8245 192.34 285.9445 ;
      RECT 191.42 285.8245 191.62 285.9445 ;
      RECT 190.7 285.8245 190.9 285.9445 ;
      RECT 189.98 285.8245 190.18 285.9445 ;
      RECT 189.26 285.8245 189.46 285.9445 ;
      RECT 188.54 285.8245 188.74 285.9445 ;
      RECT 192.5 305.625 192.7 305.745 ;
      RECT 189.62 305.625 189.82 305.745 ;
      RECT 191.42 306.041 191.62 306.161 ;
      RECT 192.14 306.041 192.34 306.161 ;
      RECT 190.7 306.041 190.9 306.161 ;
      RECT 189.98 306.041 190.18 306.161 ;
      RECT 189.26 306.041 189.46 306.161 ;
      RECT 188.54 306.041 188.74 306.161 ;
      RECT 192.5 323.3835 192.7 323.5035 ;
      RECT 189.62 323.3835 189.82 323.5035 ;
      RECT 192.14 325.9425 192.34 326.0625 ;
      RECT 191.42 325.9425 191.62 326.0625 ;
      RECT 190.7 325.9425 190.9 326.0625 ;
      RECT 189.98 325.9425 190.18 326.0625 ;
      RECT 189.26 325.9425 189.46 326.0625 ;
      RECT 188.54 325.9425 188.74 326.0625 ;
      RECT 192.5 348.339 192.7 348.459 ;
      RECT 189.62 348.339 189.82 348.459 ;
      RECT 194.3 118.324 194.5 118.444 ;
      RECT 195.02 118.084 195.22 118.204 ;
      RECT 193.58 118.084 193.78 118.204 ;
      RECT 192.86 118.084 193.06 118.204 ;
      RECT 193.58 223.558 193.78 223.678 ;
      RECT 192.86 222.885 193.06 223.005 ;
      RECT 193.58 222.885 193.78 223.005 ;
      RECT 194.3 222.885 194.5 223.005 ;
      RECT 195.02 222.885 195.22 223.005 ;
      RECT 195.02 223.558 195.22 223.678 ;
      RECT 194.3 223.798 194.5 223.918 ;
      RECT 192.86 223.798 193.06 223.918 ;
      RECT 194.66 275.1295 194.86 275.2495 ;
      RECT 193.94 275.1295 194.14 275.2495 ;
      RECT 193.22 275.1295 193.42 275.2495 ;
      RECT 195.02 274.74 195.22 274.86 ;
      RECT 194.3 274.5 194.5 274.62 ;
      RECT 193.58 274.5 193.78 274.62 ;
      RECT 192.86 274.5 193.06 274.62 ;
      RECT 194.66 277.618 194.86 277.738 ;
      RECT 193.94 277.618 194.14 277.738 ;
      RECT 193.22 277.618 193.42 277.738 ;
      RECT 194.66 279.54 194.86 279.66 ;
      RECT 193.94 279.54 194.14 279.66 ;
      RECT 193.22 279.54 193.42 279.66 ;
      RECT 194.66 282.06 194.86 282.18 ;
      RECT 193.94 282.06 194.14 282.18 ;
      RECT 193.22 282.06 193.42 282.18 ;
      RECT 195.02 285.8245 195.22 285.9445 ;
      RECT 194.3 285.8245 194.5 285.9445 ;
      RECT 193.58 285.8245 193.78 285.9445 ;
      RECT 192.86 285.8245 193.06 285.9445 ;
      RECT 195.02 306.041 195.22 306.161 ;
      RECT 194.3 306.041 194.5 306.161 ;
      RECT 192.86 306.041 193.06 306.161 ;
      RECT 193.58 306.041 193.78 306.161 ;
      RECT 192.86 325.9425 193.06 326.0625 ;
      RECT 194.3 325.9425 194.5 326.0625 ;
      RECT 195.02 325.9425 195.22 326.0625 ;
      RECT 193.58 325.9425 193.78 326.0625 ;
      RECT 199.34 118.324 199.54 118.444 ;
      RECT 198.62 118.324 198.82 118.444 ;
      RECT 200.78 118.084 200.98 118.204 ;
      RECT 200.06 118.084 200.26 118.204 ;
      RECT 201.14 170.505 201.34 170.625 ;
      RECT 199.34 223.798 199.54 223.918 ;
      RECT 199.34 222.885 199.54 223.005 ;
      RECT 200.78 222.885 200.98 223.005 ;
      RECT 200.06 222.885 200.26 223.005 ;
      RECT 198.62 222.885 198.82 223.005 ;
      RECT 200.78 223.558 200.98 223.678 ;
      RECT 200.06 223.558 200.26 223.678 ;
      RECT 198.62 223.558 198.82 223.678 ;
      RECT 200.42 282.06 200.62 282.18 ;
      RECT 199.7 282.06 199.9 282.18 ;
      RECT 198.98 282.06 199.18 282.18 ;
      RECT 199.7 279.54 199.9 279.66 ;
      RECT 198.98 279.54 199.18 279.66 ;
      RECT 200.42 279.54 200.62 279.66 ;
      RECT 200.42 277.618 200.62 277.738 ;
      RECT 199.7 277.618 199.9 277.738 ;
      RECT 198.98 277.618 199.18 277.738 ;
      RECT 200.42 275.1295 200.62 275.2495 ;
      RECT 199.7 275.1295 199.9 275.2495 ;
      RECT 198.98 275.1295 199.18 275.2495 ;
      RECT 199.34 274.74 199.54 274.86 ;
      RECT 200.06 274.5 200.26 274.62 ;
      RECT 198.62 274.5 198.82 274.62 ;
      RECT 200.78 285.8245 200.98 285.9445 ;
      RECT 200.06 285.8245 200.26 285.9445 ;
      RECT 199.34 285.8245 199.54 285.9445 ;
      RECT 198.62 285.8245 198.82 285.9445 ;
      RECT 201.14 305.625 201.34 305.745 ;
      RECT 200.78 325.9425 200.98 326.0625 ;
      RECT 200.06 325.9425 200.26 326.0625 ;
      RECT 199.34 325.9425 199.54 326.0625 ;
      RECT 198.62 325.9425 198.82 326.0625 ;
      RECT 187.82 274.74 188.02 274.86 ;
      RECT 182.06 274.74 182.26 274.86 ;
      RECT 180.62 274.74 180.82 274.86 ;
      RECT 187.1 274.5 187.3 274.62 ;
      RECT 183.5 274.5 183.7 274.62 ;
      RECT 182.78 274.5 182.98 274.62 ;
      RECT 181.34 274.5 181.54 274.62 ;
      RECT 188.18 277.858 188.38 277.978 ;
      RECT 187.46 277.858 187.66 277.978 ;
      RECT 183.14 277.618 183.34 277.738 ;
      RECT 182.42 277.618 182.62 277.738 ;
      RECT 181.7 277.618 181.9 277.738 ;
      RECT 180.26 277.618 180.46 277.738 ;
      RECT 187.82 277.26 188.02 277.38 ;
      RECT 183.5 277.26 183.7 277.38 ;
      RECT 182.06 277.26 182.26 277.38 ;
      RECT 180.62 277.26 180.82 277.38 ;
      RECT 187.1 277.02 187.3 277.14 ;
      RECT 182.78 277.02 182.98 277.14 ;
      RECT 181.34 277.02 181.54 277.14 ;
      RECT 188.18 279.78 188.38 279.9 ;
      RECT 180.26 279.54 180.46 279.66 ;
      RECT 187.46 279.54 187.66 279.66 ;
      RECT 183.14 279.54 183.34 279.66 ;
      RECT 182.42 279.54 182.62 279.66 ;
      RECT 181.7 279.54 181.9 279.66 ;
      RECT 188.18 282.3 188.38 282.42 ;
      RECT 187.46 282.06 187.66 282.18 ;
      RECT 183.14 282.06 183.34 282.18 ;
      RECT 182.42 282.06 182.62 282.18 ;
      RECT 181.7 282.06 181.9 282.18 ;
      RECT 180.26 282.06 180.46 282.18 ;
      RECT 187.82 285.8245 188.02 285.9445 ;
      RECT 187.1 285.8245 187.3 285.9445 ;
      RECT 183.5 285.8245 183.7 285.9445 ;
      RECT 182.78 285.8245 182.98 285.9445 ;
      RECT 182.06 285.8245 182.26 285.9445 ;
      RECT 181.34 285.8245 181.54 285.9445 ;
      RECT 180.62 285.8245 180.82 285.9445 ;
      RECT 180.98 305.625 181.18 305.745 ;
      RECT 187.82 306.041 188.02 306.161 ;
      RECT 187.1 306.041 187.3 306.161 ;
      RECT 183.5 306.041 183.7 306.161 ;
      RECT 182.78 306.041 182.98 306.161 ;
      RECT 182.06 306.041 182.26 306.161 ;
      RECT 181.34 306.041 181.54 306.161 ;
      RECT 180.62 306.041 180.82 306.161 ;
      RECT 180.98 323.3835 181.18 323.5035 ;
      RECT 187.82 325.9425 188.02 326.0625 ;
      RECT 187.1 325.9425 187.3 326.0625 ;
      RECT 183.5 325.9425 183.7 326.0625 ;
      RECT 182.78 325.9425 182.98 326.0625 ;
      RECT 182.06 325.9425 182.26 326.0625 ;
      RECT 181.34 325.9425 181.54 326.0625 ;
      RECT 180.62 325.9425 180.82 326.0625 ;
      RECT 180.98 348.339 181.18 348.459 ;
      RECT 192.14 118.324 192.34 118.444 ;
      RECT 189.26 118.324 189.46 118.444 ;
      RECT 188.54 118.324 188.74 118.444 ;
      RECT 191.42 118.084 191.62 118.204 ;
      RECT 190.7 118.084 190.9 118.204 ;
      RECT 189.98 118.084 190.18 118.204 ;
      RECT 192.5 170.505 192.7 170.625 ;
      RECT 189.62 170.505 189.82 170.625 ;
      RECT 188.54 223.798 188.74 223.918 ;
      RECT 190.7 223.798 190.9 223.918 ;
      RECT 191.42 223.798 191.62 223.918 ;
      RECT 189.26 223.558 189.46 223.678 ;
      RECT 189.98 223.558 190.18 223.678 ;
      RECT 192.14 223.558 192.34 223.678 ;
      RECT 190.7 222.885 190.9 223.005 ;
      RECT 192.14 222.885 192.34 223.005 ;
      RECT 189.98 222.885 190.18 223.005 ;
      RECT 189.26 222.885 189.46 223.005 ;
      RECT 188.54 222.885 188.74 223.005 ;
      RECT 191.06 275.3695 191.26 275.4895 ;
      RECT 190.34 275.3695 190.54 275.4895 ;
      RECT 188.9 275.3695 189.1 275.4895 ;
      RECT 191.78 275.1295 191.98 275.2495 ;
      RECT 189.26 274.74 189.46 274.86 ;
      RECT 191.42 274.74 191.62 274.86 ;
      RECT 190.7 274.74 190.9 274.86 ;
      RECT 192.14 274.5 192.34 274.62 ;
      RECT 189.98 274.5 190.18 274.62 ;
      RECT 188.54 274.5 188.74 274.62 ;
      RECT 192.14 277.02 192.34 277.14 ;
      RECT 191.42 277.02 191.62 277.14 ;
      RECT 189.98 277.02 190.18 277.14 ;
      RECT 188.54 277.02 188.74 277.14 ;
      RECT 191.78 277.858 191.98 277.978 ;
      RECT 191.06 277.858 191.26 277.978 ;
      RECT 190.34 277.858 190.54 277.978 ;
      RECT 188.9 277.858 189.1 277.978 ;
      RECT 190.7 277.26 190.9 277.38 ;
      RECT 189.26 277.26 189.46 277.38 ;
      RECT 191.78 279.78 191.98 279.9 ;
      RECT 191.06 279.78 191.26 279.9 ;
      RECT 190.34 279.78 190.54 279.9 ;
      RECT 188.9 279.78 189.1 279.9 ;
      RECT 191.78 282.3 191.98 282.42 ;
      RECT 191.06 282.3 191.26 282.42 ;
      RECT 190.34 282.3 190.54 282.42 ;
      RECT 179.18 118.324 179.38 118.444 ;
      RECT 179.9 118.084 180.1 118.204 ;
      RECT 178.1 170.505 178.3 170.625 ;
      RECT 175.58 223.798 175.78 223.918 ;
      RECT 177.02 223.798 177.22 223.918 ;
      RECT 177.74 223.798 177.94 223.918 ;
      RECT 179.18 222.885 179.38 223.005 ;
      RECT 179.9 222.885 180.1 223.005 ;
      RECT 179.18 223.558 179.38 223.678 ;
      RECT 179.9 223.798 180.1 223.918 ;
      RECT 177.74 222.885 177.94 223.005 ;
      RECT 177.02 222.885 177.22 223.005 ;
      RECT 176.3 222.885 176.5 223.005 ;
      RECT 175.58 222.885 175.78 223.005 ;
      RECT 178.46 223.558 178.66 223.678 ;
      RECT 176.3 223.558 176.5 223.678 ;
      RECT 179.54 275.1295 179.74 275.2495 ;
      RECT 179.9 274.74 180.1 274.86 ;
      RECT 179.18 274.74 179.38 274.86 ;
      RECT 178.82 275.3695 179.02 275.4895 ;
      RECT 177.38 275.3695 177.58 275.4895 ;
      RECT 176.66 275.3695 176.86 275.4895 ;
      RECT 175.94 275.3695 176.14 275.4895 ;
      RECT 178.46 274.74 178.66 274.86 ;
      RECT 177.02 274.74 177.22 274.86 ;
      RECT 175.58 274.74 175.78 274.86 ;
      RECT 177.74 274.5 177.94 274.62 ;
      RECT 176.3 274.5 176.5 274.62 ;
      RECT 179.54 277.618 179.74 277.738 ;
      RECT 179.9 277.02 180.1 277.14 ;
      RECT 179.18 277.02 179.38 277.14 ;
      RECT 178.82 277.858 179.02 277.978 ;
      RECT 177.38 277.858 177.58 277.978 ;
      RECT 176.66 277.858 176.86 277.978 ;
      RECT 175.94 277.858 176.14 277.978 ;
      RECT 178.46 277.26 178.66 277.38 ;
      RECT 177.74 277.26 177.94 277.38 ;
      RECT 177.02 277.26 177.22 277.38 ;
      RECT 175.58 277.26 175.78 277.38 ;
      RECT 176.3 277.02 176.5 277.14 ;
      RECT 179.54 279.78 179.74 279.9 ;
      RECT 178.82 279.78 179.02 279.9 ;
      RECT 177.38 279.78 177.58 279.9 ;
      RECT 176.66 279.78 176.86 279.9 ;
      RECT 175.94 279.78 176.14 279.9 ;
      RECT 179.54 282.3 179.74 282.42 ;
      RECT 178.82 282.3 179.02 282.42 ;
      RECT 177.38 282.3 177.58 282.42 ;
      RECT 176.66 282.3 176.86 282.42 ;
      RECT 175.94 282.3 176.14 282.42 ;
      RECT 179.9 285.8245 180.1 285.9445 ;
      RECT 179.18 285.8245 179.38 285.9445 ;
      RECT 178.46 285.8245 178.66 285.9445 ;
      RECT 177.74 285.8245 177.94 285.9445 ;
      RECT 177.02 285.8245 177.22 285.9445 ;
      RECT 176.3 285.8245 176.5 285.9445 ;
      RECT 175.58 285.8245 175.78 285.9445 ;
      RECT 178.1 305.625 178.3 305.745 ;
      RECT 178.46 306.041 178.66 306.161 ;
      RECT 177.74 306.041 177.94 306.161 ;
      RECT 177.02 306.041 177.22 306.161 ;
      RECT 176.3 306.041 176.5 306.161 ;
      RECT 175.58 306.041 175.78 306.161 ;
      RECT 179.9 306.041 180.1 306.161 ;
      RECT 179.18 306.041 179.38 306.161 ;
      RECT 178.1 323.3835 178.3 323.5035 ;
      RECT 178.46 325.9425 178.66 326.0625 ;
      RECT 177.74 325.9425 177.94 326.0625 ;
      RECT 177.02 325.9425 177.22 326.0625 ;
      RECT 176.3 325.9425 176.5 326.0625 ;
      RECT 175.58 325.9425 175.78 326.0625 ;
      RECT 179.9 325.9425 180.1 326.0625 ;
      RECT 179.18 325.9425 179.38 326.0625 ;
      RECT 178.1 348.339 178.3 348.459 ;
      RECT 187.82 118.324 188.02 118.444 ;
      RECT 182.78 118.324 182.98 118.444 ;
      RECT 182.06 118.324 182.26 118.444 ;
      RECT 180.62 118.084 180.82 118.204 ;
      RECT 181.34 118.084 181.54 118.204 ;
      RECT 183.5 118.084 183.7 118.204 ;
      RECT 187.1 118.084 187.3 118.204 ;
      RECT 180.98 170.505 181.18 170.625 ;
      RECT 182.06 223.798 182.26 223.918 ;
      RECT 182.78 223.798 182.98 223.918 ;
      RECT 187.1 223.798 187.3 223.918 ;
      RECT 180.62 223.558 180.82 223.678 ;
      RECT 180.62 222.885 180.82 223.005 ;
      RECT 181.34 222.885 181.54 223.005 ;
      RECT 182.06 222.885 182.26 223.005 ;
      RECT 182.78 222.885 182.98 223.005 ;
      RECT 183.5 222.885 183.7 223.005 ;
      RECT 187.1 222.885 187.3 223.005 ;
      RECT 187.82 222.885 188.02 223.005 ;
      RECT 187.82 223.558 188.02 223.678 ;
      RECT 183.5 223.558 183.7 223.678 ;
      RECT 181.34 223.558 181.54 223.678 ;
      RECT 188.18 275.3695 188.38 275.4895 ;
      RECT 187.46 275.3695 187.66 275.4895 ;
      RECT 183.14 275.1295 183.34 275.2495 ;
      RECT 182.42 275.1295 182.62 275.2495 ;
      RECT 181.7 275.1295 181.9 275.2495 ;
      RECT 180.26 275.1295 180.46 275.2495 ;
      RECT 170.9 275.1295 171.1 275.2495 ;
      RECT 170.18 275.1295 170.38 275.2495 ;
      RECT 168.74 275.1295 168.94 275.2495 ;
      RECT 168.02 275.1295 168.22 275.2495 ;
      RECT 168.38 274.74 168.58 274.86 ;
      RECT 166.94 274.74 167.14 274.86 ;
      RECT 166.22 274.74 166.42 274.86 ;
      RECT 164.78 274.74 164.98 274.86 ;
      RECT 170.54 274.5 170.74 274.62 ;
      RECT 169.82 274.5 170.02 274.62 ;
      RECT 171.26 274.5 171.46 274.62 ;
      RECT 169.1 274.5 169.3 274.62 ;
      RECT 167.66 274.5 167.86 274.62 ;
      RECT 165.5 274.5 165.7 274.62 ;
      RECT 164.06 274.5 164.26 274.62 ;
      RECT 171.98 274.5 172.18 274.62 ;
      RECT 167.3 277.858 167.5 277.978 ;
      RECT 165.86 277.858 166.06 277.978 ;
      RECT 165.14 277.858 165.34 277.978 ;
      RECT 164.42 277.858 164.62 277.978 ;
      RECT 171.62 277.618 171.82 277.738 ;
      RECT 170.9 277.618 171.1 277.738 ;
      RECT 170.18 277.618 170.38 277.738 ;
      RECT 168.74 277.618 168.94 277.738 ;
      RECT 168.02 277.618 168.22 277.738 ;
      RECT 168.38 277.26 168.58 277.38 ;
      RECT 166.94 277.26 167.14 277.38 ;
      RECT 164.78 277.26 164.98 277.38 ;
      RECT 164.06 277.26 164.26 277.38 ;
      RECT 171.98 277.02 172.18 277.14 ;
      RECT 171.26 277.02 171.46 277.14 ;
      RECT 170.54 277.02 170.74 277.14 ;
      RECT 169.82 277.02 170.02 277.14 ;
      RECT 169.1 277.02 169.3 277.14 ;
      RECT 167.66 277.02 167.86 277.14 ;
      RECT 166.22 277.02 166.42 277.14 ;
      RECT 165.5 277.02 165.7 277.14 ;
      RECT 167.3 279.78 167.5 279.9 ;
      RECT 165.86 279.78 166.06 279.9 ;
      RECT 165.14 279.78 165.34 279.9 ;
      RECT 164.42 279.78 164.62 279.9 ;
      RECT 171.62 279.54 171.82 279.66 ;
      RECT 170.9 279.54 171.1 279.66 ;
      RECT 170.18 279.54 170.38 279.66 ;
      RECT 168.74 279.54 168.94 279.66 ;
      RECT 168.02 279.54 168.22 279.66 ;
      RECT 167.3 282.3 167.5 282.42 ;
      RECT 165.86 282.3 166.06 282.42 ;
      RECT 165.14 282.3 165.34 282.42 ;
      RECT 164.42 282.3 164.62 282.42 ;
      RECT 171.62 282.06 171.82 282.18 ;
      RECT 170.9 282.06 171.1 282.18 ;
      RECT 170.18 282.06 170.38 282.18 ;
      RECT 168.74 282.06 168.94 282.18 ;
      RECT 168.02 282.06 168.22 282.18 ;
      RECT 171.98 285.8245 172.18 285.9445 ;
      RECT 171.26 285.8245 171.46 285.9445 ;
      RECT 170.54 285.8245 170.74 285.9445 ;
      RECT 169.82 285.8245 170.02 285.9445 ;
      RECT 169.1 285.8245 169.3 285.9445 ;
      RECT 168.38 285.8245 168.58 285.9445 ;
      RECT 167.66 285.8245 167.86 285.9445 ;
      RECT 166.94 285.8245 167.14 285.9445 ;
      RECT 166.22 285.8245 166.42 285.9445 ;
      RECT 165.5 285.8245 165.7 285.9445 ;
      RECT 164.78 285.8245 164.98 285.9445 ;
      RECT 164.06 285.8245 164.26 285.9445 ;
      RECT 169.46 305.625 169.66 305.745 ;
      RECT 166.58 305.625 166.78 305.745 ;
      RECT 171.98 306.041 172.18 306.161 ;
      RECT 171.26 306.041 171.46 306.161 ;
      RECT 170.54 306.041 170.74 306.161 ;
      RECT 169.82 306.041 170.02 306.161 ;
      RECT 169.1 306.041 169.3 306.161 ;
      RECT 168.38 306.041 168.58 306.161 ;
      RECT 167.66 306.041 167.86 306.161 ;
      RECT 166.94 306.041 167.14 306.161 ;
      RECT 166.22 306.041 166.42 306.161 ;
      RECT 165.5 306.041 165.7 306.161 ;
      RECT 164.78 306.041 164.98 306.161 ;
      RECT 164.06 306.041 164.26 306.161 ;
      RECT 169.46 323.3835 169.66 323.5035 ;
      RECT 166.58 323.3835 166.78 323.5035 ;
      RECT 164.06 325.9425 164.26 326.0625 ;
      RECT 171.98 325.9425 172.18 326.0625 ;
      RECT 171.26 325.9425 171.46 326.0625 ;
      RECT 170.54 325.9425 170.74 326.0625 ;
      RECT 169.82 325.9425 170.02 326.0625 ;
      RECT 169.1 325.9425 169.3 326.0625 ;
      RECT 168.38 325.9425 168.58 326.0625 ;
      RECT 167.66 325.9425 167.86 326.0625 ;
      RECT 166.94 325.9425 167.14 326.0625 ;
      RECT 166.22 325.9425 166.42 326.0625 ;
      RECT 165.5 325.9425 165.7 326.0625 ;
      RECT 164.78 325.9425 164.98 326.0625 ;
      RECT 169.46 348.339 169.66 348.459 ;
      RECT 166.58 348.339 166.78 348.459 ;
      RECT 177.74 118.324 177.94 118.444 ;
      RECT 176.3 118.324 176.5 118.444 ;
      RECT 175.58 118.084 175.78 118.204 ;
      RECT 177.02 118.084 177.22 118.204 ;
      RECT 178.46 118.084 178.66 118.204 ;
      RECT 165.5 219.06 165.7 219.18 ;
      RECT 164.06 219.06 164.26 219.18 ;
      RECT 168.38 223.798 168.58 223.918 ;
      RECT 170.54 223.798 170.74 223.918 ;
      RECT 171.98 223.798 172.18 223.918 ;
      RECT 166.94 223.798 167.14 223.918 ;
      RECT 164.06 223.558 164.26 223.678 ;
      RECT 164.78 223.558 164.98 223.678 ;
      RECT 165.5 223.558 165.7 223.678 ;
      RECT 166.22 223.558 166.42 223.678 ;
      RECT 167.66 223.558 167.86 223.678 ;
      RECT 169.46 222.84 169.66 222.96 ;
      RECT 166.58 222.84 166.78 222.96 ;
      RECT 171.26 222.885 171.46 223.005 ;
      RECT 171.26 223.558 171.46 223.678 ;
      RECT 169.82 223.558 170.02 223.678 ;
      RECT 169.1 223.558 169.3 223.678 ;
      RECT 169.46 258.99 169.66 259.11 ;
      RECT 166.58 258.75 166.78 258.87 ;
      RECT 171.98 261.9 172.18 262.02 ;
      RECT 171.26 261.9 171.46 262.02 ;
      RECT 170.54 261.9 170.74 262.02 ;
      RECT 169.82 261.9 170.02 262.02 ;
      RECT 169.1 261.9 169.3 262.02 ;
      RECT 167.66 261.9 167.86 262.02 ;
      RECT 166.94 261.9 167.14 262.02 ;
      RECT 166.22 261.9 166.42 262.02 ;
      RECT 164.78 261.9 164.98 262.02 ;
      RECT 166.58 261.51 166.78 261.63 ;
      RECT 169.46 261.27 169.66 261.39 ;
      RECT 166.58 260.25 166.78 260.37 ;
      RECT 169.46 260.01 169.66 260.13 ;
      RECT 169.82 264.66 170.02 264.78 ;
      RECT 168.38 264.66 168.58 264.78 ;
      RECT 166.94 264.66 167.14 264.78 ;
      RECT 165.5 264.66 165.7 264.78 ;
      RECT 164.78 264.66 164.98 264.78 ;
      RECT 170.54 264.42 170.74 264.54 ;
      RECT 169.1 264.42 169.3 264.54 ;
      RECT 167.66 264.42 167.86 264.54 ;
      RECT 166.22 264.42 166.42 264.54 ;
      RECT 164.06 264.42 164.26 264.54 ;
      RECT 171.98 264.42 172.18 264.54 ;
      RECT 171.26 264.42 171.46 264.54 ;
      RECT 169.46 263.79 169.66 263.91 ;
      RECT 166.58 263.79 166.78 263.91 ;
      RECT 169.46 262.77 169.66 262.89 ;
      RECT 166.58 262.53 166.78 262.65 ;
      RECT 168.38 262.14 168.58 262.26 ;
      RECT 165.5 262.14 165.7 262.26 ;
      RECT 164.06 262.14 164.26 262.26 ;
      RECT 166.22 267.18 166.42 267.3 ;
      RECT 164.06 267.18 164.26 267.3 ;
      RECT 171.98 266.94 172.18 267.06 ;
      RECT 171.26 266.94 171.46 267.06 ;
      RECT 170.54 266.94 170.74 267.06 ;
      RECT 169.82 266.94 170.02 267.06 ;
      RECT 169.1 266.94 169.3 267.06 ;
      RECT 168.38 266.94 168.58 267.06 ;
      RECT 167.66 266.94 167.86 267.06 ;
      RECT 166.94 266.94 167.14 267.06 ;
      RECT 165.5 266.94 165.7 267.06 ;
      RECT 164.78 266.94 164.98 267.06 ;
      RECT 169.46 266.2885 169.66 266.4085 ;
      RECT 166.58 266.2885 166.78 266.4085 ;
      RECT 169.46 270.09 169.66 270.21 ;
      RECT 166.58 270.09 166.78 270.21 ;
      RECT 170.54 269.7 170.74 269.82 ;
      RECT 167.66 269.7 167.86 269.82 ;
      RECT 166.22 269.7 166.42 269.82 ;
      RECT 164.06 269.7 164.26 269.82 ;
      RECT 171.98 269.46 172.18 269.58 ;
      RECT 171.26 269.46 171.46 269.58 ;
      RECT 169.82 269.46 170.02 269.58 ;
      RECT 169.1 269.46 169.3 269.58 ;
      RECT 168.38 269.46 168.58 269.58 ;
      RECT 166.94 269.46 167.14 269.58 ;
      RECT 165.5 269.46 165.7 269.58 ;
      RECT 164.78 269.46 164.98 269.58 ;
      RECT 169.46 268.83 169.66 268.95 ;
      RECT 166.58 268.83 166.78 268.95 ;
      RECT 169.46 267.81 169.66 267.93 ;
      RECT 166.58 267.81 166.78 267.93 ;
      RECT 169.46 271.35 169.66 271.47 ;
      RECT 166.58 271.35 166.78 271.47 ;
      RECT 164.06 272.22 164.26 272.34 ;
      RECT 165.5 272.22 165.7 272.34 ;
      RECT 171.98 271.98 172.18 272.1 ;
      RECT 171.26 271.98 171.46 272.1 ;
      RECT 170.54 271.98 170.74 272.1 ;
      RECT 169.82 271.98 170.02 272.1 ;
      RECT 169.1 271.98 169.3 272.1 ;
      RECT 168.38 271.98 168.58 272.1 ;
      RECT 167.66 271.98 167.86 272.1 ;
      RECT 166.94 271.98 167.14 272.1 ;
      RECT 166.22 271.98 166.42 272.1 ;
      RECT 164.78 271.98 164.98 272.1 ;
      RECT 167.3 275.3695 167.5 275.4895 ;
      RECT 165.86 275.3695 166.06 275.4895 ;
      RECT 165.14 275.3695 165.34 275.4895 ;
      RECT 164.42 275.3695 164.62 275.4895 ;
      RECT 171.62 275.1295 171.82 275.2495 ;
      RECT 165.5 196.38 165.7 196.5 ;
      RECT 164.78 196.38 164.98 196.5 ;
      RECT 164.06 196.38 164.26 196.5 ;
      RECT 166.58 195.12 166.78 195.24 ;
      RECT 169.46 195.12 169.66 195.24 ;
      RECT 168.38 199.14 168.58 199.26 ;
      RECT 166.94 199.14 167.14 199.26 ;
      RECT 165.5 199.14 165.7 199.26 ;
      RECT 164.06 199.14 164.26 199.26 ;
      RECT 164.78 198.9 164.98 199.02 ;
      RECT 166.22 198.9 166.42 199.02 ;
      RECT 167.66 198.9 167.86 199.02 ;
      RECT 169.1 198.9 169.3 199.02 ;
      RECT 169.82 198.9 170.02 199.02 ;
      RECT 169.46 197.64 169.66 197.76 ;
      RECT 166.58 197.64 166.78 197.76 ;
      RECT 168.38 196.62 168.58 196.74 ;
      RECT 166.22 196.62 166.42 196.74 ;
      RECT 164.06 201.66 164.26 201.78 ;
      RECT 165.5 201.66 165.7 201.78 ;
      RECT 168.38 201.66 168.58 201.78 ;
      RECT 164.78 201.42 164.98 201.54 ;
      RECT 166.22 201.42 166.42 201.54 ;
      RECT 166.94 201.42 167.14 201.54 ;
      RECT 169.82 201.42 170.02 201.54 ;
      RECT 169.1 201.42 169.3 201.54 ;
      RECT 167.66 201.42 167.86 201.54 ;
      RECT 169.46 200.16 169.66 200.28 ;
      RECT 166.58 200.16 166.78 200.28 ;
      RECT 168.38 204.18 168.58 204.3 ;
      RECT 166.94 204.18 167.14 204.3 ;
      RECT 164.06 204.18 164.26 204.3 ;
      RECT 164.78 203.94 164.98 204.06 ;
      RECT 165.5 203.94 165.7 204.06 ;
      RECT 166.22 203.94 166.42 204.06 ;
      RECT 167.66 203.94 167.86 204.06 ;
      RECT 169.1 203.94 169.3 204.06 ;
      RECT 169.82 203.94 170.02 204.06 ;
      RECT 166.58 202.68 166.78 202.8 ;
      RECT 169.46 202.68 169.66 202.8 ;
      RECT 164.06 206.7 164.26 206.82 ;
      RECT 166.94 206.7 167.14 206.82 ;
      RECT 168.38 206.7 168.58 206.82 ;
      RECT 169.82 206.46 170.02 206.58 ;
      RECT 169.1 206.46 169.3 206.58 ;
      RECT 167.66 206.46 167.86 206.58 ;
      RECT 166.22 206.46 166.42 206.58 ;
      RECT 165.5 206.46 165.7 206.58 ;
      RECT 164.78 206.46 164.98 206.58 ;
      RECT 166.58 205.2 166.78 205.32 ;
      RECT 169.46 205.2 169.66 205.32 ;
      RECT 166.58 210.24 166.78 210.36 ;
      RECT 169.46 210.24 169.66 210.36 ;
      RECT 167.66 209.22 167.86 209.34 ;
      RECT 166.22 209.22 166.42 209.34 ;
      RECT 164.78 209.22 164.98 209.34 ;
      RECT 169.82 208.98 170.02 209.1 ;
      RECT 169.1 208.98 169.3 209.1 ;
      RECT 168.38 208.98 168.58 209.1 ;
      RECT 166.94 208.98 167.14 209.1 ;
      RECT 165.5 208.98 165.7 209.1 ;
      RECT 164.06 208.98 164.26 209.1 ;
      RECT 166.58 207.72 166.78 207.84 ;
      RECT 169.46 207.72 169.66 207.84 ;
      RECT 166.58 212.76 166.78 212.88 ;
      RECT 169.46 212.76 169.66 212.88 ;
      RECT 169.1 211.74 169.3 211.86 ;
      RECT 166.94 211.74 167.14 211.86 ;
      RECT 164.78 211.74 164.98 211.86 ;
      RECT 169.82 211.5 170.02 211.62 ;
      RECT 168.38 211.5 168.58 211.62 ;
      RECT 167.66 211.5 167.86 211.62 ;
      RECT 166.22 211.5 166.42 211.62 ;
      RECT 165.5 211.5 165.7 211.62 ;
      RECT 164.06 211.5 164.26 211.62 ;
      RECT 166.58 215.28 166.78 215.4 ;
      RECT 169.46 215.28 169.66 215.4 ;
      RECT 168.38 214.26 168.58 214.38 ;
      RECT 166.94 214.26 167.14 214.38 ;
      RECT 165.5 214.26 165.7 214.38 ;
      RECT 164.06 214.26 164.26 214.38 ;
      RECT 169.82 214.02 170.02 214.14 ;
      RECT 169.1 214.02 169.3 214.14 ;
      RECT 167.66 214.02 167.86 214.14 ;
      RECT 166.22 214.02 166.42 214.14 ;
      RECT 164.78 214.02 164.98 214.14 ;
      RECT 168.38 216.78 168.58 216.9 ;
      RECT 166.94 216.78 167.14 216.9 ;
      RECT 165.5 216.78 165.7 216.9 ;
      RECT 164.78 216.78 164.98 216.9 ;
      RECT 164.06 216.54 164.26 216.66 ;
      RECT 169.82 216.54 170.02 216.66 ;
      RECT 169.1 216.54 169.3 216.66 ;
      RECT 167.66 216.54 167.86 216.66 ;
      RECT 166.22 216.54 166.42 216.66 ;
      RECT 164.78 219.3 164.98 219.42 ;
      RECT 168.38 219.3 168.58 219.42 ;
      RECT 169.82 219.06 170.02 219.18 ;
      RECT 169.1 219.06 169.3 219.18 ;
      RECT 167.66 219.06 167.86 219.18 ;
      RECT 166.94 219.06 167.14 219.18 ;
      RECT 166.22 219.06 166.42 219.18 ;
      RECT 171.26 118.324 171.46 118.444 ;
      RECT 170.54 118.324 170.74 118.444 ;
      RECT 169.82 118.324 170.02 118.444 ;
      RECT 166.94 118.324 167.14 118.444 ;
      RECT 165.5 118.324 165.7 118.444 ;
      RECT 164.78 118.324 164.98 118.444 ;
      RECT 171.98 118.084 172.18 118.204 ;
      RECT 164.06 118.084 164.26 118.204 ;
      RECT 166.22 118.084 166.42 118.204 ;
      RECT 167.66 118.084 167.86 118.204 ;
      RECT 168.38 118.084 168.58 118.204 ;
      RECT 169.1 118.084 169.3 118.204 ;
      RECT 166.58 155.04 166.78 155.16 ;
      RECT 169.46 154.8 169.66 154.92 ;
      RECT 168.38 156.3 168.58 156.42 ;
      RECT 166.94 156.3 167.14 156.42 ;
      RECT 164.78 156.3 164.98 156.42 ;
      RECT 169.82 156.06 170.02 156.18 ;
      RECT 164.06 156.06 164.26 156.18 ;
      RECT 165.5 156.06 165.7 156.18 ;
      RECT 166.22 156.06 166.42 156.18 ;
      RECT 167.66 156.06 167.86 156.18 ;
      RECT 169.1 156.06 169.3 156.18 ;
      RECT 164.78 166.38 164.98 166.5 ;
      RECT 166.94 166.38 167.14 166.5 ;
      RECT 168.38 166.38 168.58 166.5 ;
      RECT 169.1 166.14 169.3 166.26 ;
      RECT 167.66 166.14 167.86 166.26 ;
      RECT 166.22 166.14 166.42 166.26 ;
      RECT 165.5 166.14 165.7 166.26 ;
      RECT 164.06 166.14 164.26 166.26 ;
      RECT 168.38 168.9 168.58 169.02 ;
      RECT 166.94 168.9 167.14 169.02 ;
      RECT 169.1 168.66 169.3 168.78 ;
      RECT 167.66 168.66 167.86 168.78 ;
      RECT 166.22 168.66 166.42 168.78 ;
      RECT 165.5 168.66 165.7 168.78 ;
      RECT 164.78 168.66 164.98 168.78 ;
      RECT 164.06 168.66 164.26 168.78 ;
      RECT 166.58 167.4 166.78 167.52 ;
      RECT 164.78 171.42 164.98 171.54 ;
      RECT 166.94 171.42 167.14 171.54 ;
      RECT 168.38 171.42 168.58 171.54 ;
      RECT 169.1 171.18 169.3 171.3 ;
      RECT 167.66 171.18 167.86 171.3 ;
      RECT 166.22 171.18 166.42 171.3 ;
      RECT 165.5 171.18 165.7 171.3 ;
      RECT 164.06 171.18 164.26 171.3 ;
      RECT 169.46 170.505 169.66 170.625 ;
      RECT 166.58 170.505 166.78 170.625 ;
      RECT 166.58 169.92 166.78 170.04 ;
      RECT 164.78 173.94 164.98 174.06 ;
      RECT 166.94 173.94 167.14 174.06 ;
      RECT 168.38 173.94 168.58 174.06 ;
      RECT 169.1 173.7 169.3 173.82 ;
      RECT 167.66 173.7 167.86 173.82 ;
      RECT 166.22 173.7 166.42 173.82 ;
      RECT 165.5 173.7 165.7 173.82 ;
      RECT 164.06 173.7 164.26 173.82 ;
      RECT 166.58 172.44 166.78 172.56 ;
      RECT 166.58 177.48 166.78 177.6 ;
      RECT 164.06 176.46 164.26 176.58 ;
      RECT 166.94 176.46 167.14 176.58 ;
      RECT 168.38 176.46 168.58 176.58 ;
      RECT 169.1 176.22 169.3 176.34 ;
      RECT 167.66 176.22 167.86 176.34 ;
      RECT 166.22 176.22 166.42 176.34 ;
      RECT 165.5 176.22 165.7 176.34 ;
      RECT 164.78 176.22 164.98 176.34 ;
      RECT 166.58 174.96 166.78 175.08 ;
      RECT 168.38 178.98 168.58 179.1 ;
      RECT 166.94 178.98 167.14 179.1 ;
      RECT 165.5 178.98 165.7 179.1 ;
      RECT 164.06 178.98 164.26 179.1 ;
      RECT 164.78 178.74 164.98 178.86 ;
      RECT 166.22 178.74 166.42 178.86 ;
      RECT 167.66 178.74 167.86 178.86 ;
      RECT 169.1 178.74 169.3 178.86 ;
      RECT 169.82 193.86 170.02 193.98 ;
      RECT 169.1 193.86 169.3 193.98 ;
      RECT 167.66 193.86 167.86 193.98 ;
      RECT 166.22 193.86 166.42 193.98 ;
      RECT 165.5 193.86 165.7 193.98 ;
      RECT 164.78 193.86 164.98 193.98 ;
      RECT 166.58 192.6 166.78 192.72 ;
      RECT 169.46 192.6 169.66 192.72 ;
      RECT 168.38 191.58 168.58 191.7 ;
      RECT 169.82 191.34 170.02 191.46 ;
      RECT 169.1 191.34 169.3 191.46 ;
      RECT 167.66 191.34 167.86 191.46 ;
      RECT 166.94 191.34 167.14 191.46 ;
      RECT 166.22 191.34 166.42 191.46 ;
      RECT 165.5 191.34 165.7 191.46 ;
      RECT 164.78 191.34 164.98 191.46 ;
      RECT 164.06 191.34 164.26 191.46 ;
      RECT 168.38 194.1 168.58 194.22 ;
      RECT 166.94 194.1 167.14 194.22 ;
      RECT 164.06 194.1 164.26 194.22 ;
      RECT 169.82 196.38 170.02 196.5 ;
      RECT 169.1 196.38 169.3 196.5 ;
      RECT 167.66 196.38 167.86 196.5 ;
      RECT 166.94 196.38 167.14 196.5 ;
      RECT 157.94 261.27 158.14 261.39 ;
      RECT 157.94 260.01 158.14 260.13 ;
      RECT 160.46 264.66 160.66 264.78 ;
      RECT 159.74 264.66 159.94 264.78 ;
      RECT 158.3 264.66 158.5 264.78 ;
      RECT 156.86 264.66 157.06 264.78 ;
      RECT 157.58 264.42 157.78 264.54 ;
      RECT 159.02 264.42 159.22 264.54 ;
      RECT 157.94 264.03 158.14 264.15 ;
      RECT 157.94 262.77 158.14 262.89 ;
      RECT 159.74 262.14 159.94 262.26 ;
      RECT 156.86 262.14 157.06 262.26 ;
      RECT 156.14 264.42 156.34 264.54 ;
      RECT 156.14 262.14 156.34 262.26 ;
      RECT 159.74 267.18 159.94 267.3 ;
      RECT 159.02 267.18 159.22 267.3 ;
      RECT 158.3 267.18 158.5 267.3 ;
      RECT 160.46 266.94 160.66 267.06 ;
      RECT 157.58 266.94 157.78 267.06 ;
      RECT 156.86 266.94 157.06 267.06 ;
      RECT 157.94 266.2885 158.14 266.4085 ;
      RECT 156.14 267.18 156.34 267.3 ;
      RECT 159.74 269.7 159.94 269.82 ;
      RECT 159.02 269.7 159.22 269.82 ;
      RECT 156.86 269.7 157.06 269.82 ;
      RECT 160.46 269.46 160.66 269.58 ;
      RECT 158.3 269.46 158.5 269.58 ;
      RECT 157.58 269.46 157.78 269.58 ;
      RECT 157.94 269.07 158.14 269.19 ;
      RECT 157.94 267.81 158.14 267.93 ;
      RECT 156.14 269.46 156.34 269.58 ;
      RECT 157.94 271.59 158.14 271.71 ;
      RECT 157.94 270.33 158.14 270.45 ;
      RECT 159.74 272.22 159.94 272.34 ;
      RECT 158.3 272.22 158.5 272.34 ;
      RECT 157.58 272.22 157.78 272.34 ;
      RECT 160.46 271.98 160.66 272.1 ;
      RECT 159.02 271.98 159.22 272.1 ;
      RECT 156.86 271.98 157.06 272.1 ;
      RECT 156.14 272.22 156.34 272.34 ;
      RECT 160.1 275.3695 160.3 275.4895 ;
      RECT 159.38 275.1295 159.58 275.2495 ;
      RECT 158.66 275.1295 158.86 275.2495 ;
      RECT 157.22 275.1295 157.42 275.2495 ;
      RECT 160.46 274.74 160.66 274.86 ;
      RECT 158.3 274.74 158.5 274.86 ;
      RECT 157.58 274.74 157.78 274.86 ;
      RECT 159.74 274.5 159.94 274.62 ;
      RECT 159.02 274.5 159.22 274.62 ;
      RECT 156.86 274.5 157.06 274.62 ;
      RECT 155.78 275.1295 155.98 275.2495 ;
      RECT 156.14 274.74 156.34 274.86 ;
      RECT 156.5 275.1295 156.7 275.2495 ;
      RECT 160.1 277.858 160.3 277.978 ;
      RECT 159.38 277.618 159.58 277.738 ;
      RECT 158.66 277.618 158.86 277.738 ;
      RECT 157.22 277.618 157.42 277.738 ;
      RECT 159.74 277.26 159.94 277.38 ;
      RECT 158.3 277.26 158.5 277.38 ;
      RECT 157.58 277.26 157.78 277.38 ;
      RECT 160.46 277.02 160.66 277.14 ;
      RECT 159.02 277.02 159.22 277.14 ;
      RECT 156.86 277.02 157.06 277.14 ;
      RECT 156.14 277.26 156.34 277.38 ;
      RECT 155.78 277.618 155.98 277.738 ;
      RECT 156.5 277.618 156.7 277.738 ;
      RECT 160.1 279.78 160.3 279.9 ;
      RECT 159.38 279.54 159.58 279.66 ;
      RECT 158.66 279.54 158.86 279.66 ;
      RECT 157.22 279.54 157.42 279.66 ;
      RECT 155.78 279.54 155.98 279.66 ;
      RECT 156.5 279.54 156.7 279.66 ;
      RECT 160.1 282.3 160.3 282.42 ;
      RECT 159.38 282.06 159.58 282.18 ;
      RECT 158.66 282.06 158.86 282.18 ;
      RECT 157.22 282.06 157.42 282.18 ;
      RECT 155.78 282.06 155.98 282.18 ;
      RECT 156.5 282.06 156.7 282.18 ;
      RECT 160.46 285.8245 160.66 285.9445 ;
      RECT 159.74 285.8245 159.94 285.9445 ;
      RECT 159.02 285.8245 159.22 285.9445 ;
      RECT 158.3 285.8245 158.5 285.9445 ;
      RECT 157.58 285.8245 157.78 285.9445 ;
      RECT 156.86 285.8245 157.06 285.9445 ;
      RECT 156.14 285.8245 156.34 285.9445 ;
      RECT 157.94 305.625 158.14 305.745 ;
      RECT 156.14 306.041 156.34 306.161 ;
      RECT 160.46 306.041 160.66 306.161 ;
      RECT 156.86 306.041 157.06 306.161 ;
      RECT 157.58 306.041 157.78 306.161 ;
      RECT 159.02 306.041 159.22 306.161 ;
      RECT 158.3 306.041 158.5 306.161 ;
      RECT 159.74 306.041 159.94 306.161 ;
      RECT 157.94 323.3835 158.14 323.5035 ;
      RECT 156.14 325.9425 156.34 326.0625 ;
      RECT 156.86 325.9425 157.06 326.0625 ;
      RECT 157.58 325.9425 157.78 326.0625 ;
      RECT 158.3 325.9425 158.5 326.0625 ;
      RECT 159.02 325.9425 159.22 326.0625 ;
      RECT 159.74 325.9425 159.94 326.0625 ;
      RECT 160.46 325.9425 160.66 326.0625 ;
      RECT 157.94 348.339 158.14 348.459 ;
      RECT 158.3 191.58 158.5 191.7 ;
      RECT 156.86 191.58 157.06 191.7 ;
      RECT 160.46 191.34 160.66 191.46 ;
      RECT 157.58 191.34 157.78 191.46 ;
      RECT 156.14 191.34 156.34 191.46 ;
      RECT 156.14 193.86 156.34 193.98 ;
      RECT 159.74 194.1 159.94 194.22 ;
      RECT 158.3 194.1 158.5 194.22 ;
      RECT 157.58 194.1 157.78 194.22 ;
      RECT 156.86 194.1 157.06 194.22 ;
      RECT 157.94 195.36 158.14 195.48 ;
      RECT 156.86 196.38 157.06 196.5 ;
      RECT 159.02 196.38 159.22 196.5 ;
      RECT 160.46 196.38 160.66 196.5 ;
      RECT 157.58 196.62 157.78 196.74 ;
      RECT 158.3 196.62 158.5 196.74 ;
      RECT 159.74 196.62 159.94 196.74 ;
      RECT 157.94 197.88 158.14 198 ;
      RECT 160.46 198.9 160.66 199.02 ;
      RECT 159.74 198.9 159.94 199.02 ;
      RECT 158.3 198.9 158.5 199.02 ;
      RECT 156.86 198.9 157.06 199.02 ;
      RECT 157.58 199.14 157.78 199.26 ;
      RECT 159.02 199.14 159.22 199.26 ;
      RECT 156.14 196.62 156.34 196.74 ;
      RECT 156.14 199.14 156.34 199.26 ;
      RECT 157.94 200.4 158.14 200.52 ;
      RECT 160.46 201.42 160.66 201.54 ;
      RECT 159.74 201.42 159.94 201.54 ;
      RECT 158.3 201.42 158.5 201.54 ;
      RECT 159.02 201.66 159.22 201.78 ;
      RECT 157.58 201.66 157.78 201.78 ;
      RECT 156.86 201.66 157.06 201.78 ;
      RECT 156.14 201.42 156.34 201.54 ;
      RECT 156.14 204.18 156.34 204.3 ;
      RECT 157.94 202.92 158.14 203.04 ;
      RECT 160.46 203.94 160.66 204.06 ;
      RECT 159.74 203.94 159.94 204.06 ;
      RECT 156.86 203.94 157.06 204.06 ;
      RECT 157.58 204.18 157.78 204.3 ;
      RECT 158.3 204.18 158.5 204.3 ;
      RECT 159.02 204.18 159.22 204.3 ;
      RECT 156.14 206.7 156.34 206.82 ;
      RECT 157.94 205.44 158.14 205.56 ;
      RECT 156.86 206.46 157.06 206.58 ;
      RECT 158.3 206.46 158.5 206.58 ;
      RECT 159.02 206.46 159.22 206.58 ;
      RECT 160.46 206.7 160.66 206.82 ;
      RECT 159.74 206.7 159.94 206.82 ;
      RECT 157.58 206.7 157.78 206.82 ;
      RECT 156.14 208.98 156.34 209.1 ;
      RECT 157.94 207.96 158.14 208.08 ;
      RECT 157.58 208.98 157.78 209.1 ;
      RECT 159.02 208.98 159.22 209.1 ;
      RECT 156.86 209.22 157.06 209.34 ;
      RECT 158.3 209.22 158.5 209.34 ;
      RECT 159.74 209.22 159.94 209.34 ;
      RECT 160.46 209.22 160.66 209.34 ;
      RECT 157.94 210.24 158.14 210.36 ;
      RECT 156.14 211.5 156.34 211.62 ;
      RECT 157.58 211.5 157.78 211.62 ;
      RECT 159.02 211.5 159.22 211.62 ;
      RECT 156.86 211.74 157.06 211.86 ;
      RECT 158.3 211.74 158.5 211.86 ;
      RECT 159.74 211.74 159.94 211.86 ;
      RECT 160.46 211.74 160.66 211.86 ;
      RECT 157.94 212.76 158.14 212.88 ;
      RECT 156.14 214.26 156.34 214.38 ;
      RECT 156.86 214.02 157.06 214.14 ;
      RECT 159.02 214.02 159.22 214.14 ;
      RECT 159.74 214.02 159.94 214.14 ;
      RECT 160.46 214.02 160.66 214.14 ;
      RECT 157.58 214.26 157.78 214.38 ;
      RECT 158.3 214.26 158.5 214.38 ;
      RECT 157.94 215.28 158.14 215.4 ;
      RECT 156.14 216.78 156.34 216.9 ;
      RECT 157.58 216.54 157.78 216.66 ;
      RECT 158.3 216.54 158.5 216.66 ;
      RECT 159.02 216.54 159.22 216.66 ;
      RECT 160.46 216.54 160.66 216.66 ;
      RECT 156.86 216.78 157.06 216.9 ;
      RECT 159.74 216.78 159.94 216.9 ;
      RECT 156.14 219.06 156.34 219.18 ;
      RECT 157.58 219.06 157.78 219.18 ;
      RECT 159.02 219.06 159.22 219.18 ;
      RECT 160.46 219.06 160.66 219.18 ;
      RECT 156.86 219.3 157.06 219.42 ;
      RECT 158.3 219.3 158.5 219.42 ;
      RECT 159.74 219.3 159.94 219.42 ;
      RECT 156.14 223.558 156.34 223.678 ;
      RECT 156.86 223.798 157.06 223.918 ;
      RECT 157.58 223.798 157.78 223.918 ;
      RECT 158.3 223.798 158.5 223.918 ;
      RECT 159.02 223.798 159.22 223.918 ;
      RECT 160.46 223.798 160.66 223.918 ;
      RECT 159.74 223.558 159.94 223.678 ;
      RECT 157.94 222.84 158.14 222.96 ;
      RECT 157.94 258.99 158.14 259.11 ;
      RECT 160.46 261.9 160.66 262.02 ;
      RECT 159.02 261.9 159.22 262.02 ;
      RECT 158.3 261.9 158.5 262.02 ;
      RECT 157.58 261.9 157.78 262.02 ;
      RECT 153.62 279.78 153.82 279.9 ;
      RECT 154.34 279.78 154.54 279.9 ;
      RECT 147.86 282.3 148.06 282.42 ;
      RECT 148.58 282.3 148.78 282.42 ;
      RECT 152.9 282.3 153.1 282.42 ;
      RECT 153.62 282.3 153.82 282.42 ;
      RECT 154.34 282.3 154.54 282.42 ;
      RECT 147.5 285.8245 147.7 285.9445 ;
      RECT 148.22 285.8245 148.42 285.9445 ;
      RECT 148.94 285.8245 149.14 285.9445 ;
      RECT 152.54 285.8245 152.74 285.9445 ;
      RECT 153.26 285.8245 153.46 285.9445 ;
      RECT 153.98 285.8245 154.18 285.9445 ;
      RECT 154.7 285.8245 154.9 285.9445 ;
      RECT 155.42 285.8245 155.62 285.9445 ;
      RECT 155.06 305.625 155.26 305.745 ;
      RECT 148.94 306.041 149.14 306.161 ;
      RECT 148.22 306.041 148.42 306.161 ;
      RECT 147.5 306.041 147.7 306.161 ;
      RECT 152.54 306.041 152.74 306.161 ;
      RECT 153.26 306.041 153.46 306.161 ;
      RECT 153.98 306.041 154.18 306.161 ;
      RECT 154.7 306.041 154.9 306.161 ;
      RECT 155.42 306.041 155.62 306.161 ;
      RECT 155.06 323.3835 155.26 323.5035 ;
      RECT 153.26 325.9425 153.46 326.0625 ;
      RECT 152.54 325.9425 152.74 326.0625 ;
      RECT 148.94 325.9425 149.14 326.0625 ;
      RECT 148.22 325.9425 148.42 326.0625 ;
      RECT 147.5 325.9425 147.7 326.0625 ;
      RECT 155.42 325.9425 155.62 326.0625 ;
      RECT 154.7 325.9425 154.9 326.0625 ;
      RECT 153.98 325.9425 154.18 326.0625 ;
      RECT 155.06 348.339 155.26 348.459 ;
      RECT 156.14 118.324 156.34 118.444 ;
      RECT 160.46 118.324 160.66 118.444 ;
      RECT 159.02 118.324 159.22 118.444 ;
      RECT 157.58 118.324 157.78 118.444 ;
      RECT 156.86 118.084 157.06 118.204 ;
      RECT 158.3 118.084 158.5 118.204 ;
      RECT 159.74 118.084 159.94 118.204 ;
      RECT 157.94 155.04 158.14 155.16 ;
      RECT 156.14 156.06 156.34 156.18 ;
      RECT 159.74 156.06 159.94 156.18 ;
      RECT 158.3 156.06 158.5 156.18 ;
      RECT 156.86 156.06 157.06 156.18 ;
      RECT 157.58 156.3 157.78 156.42 ;
      RECT 159.02 156.3 159.22 156.42 ;
      RECT 160.46 156.3 160.66 156.42 ;
      RECT 156.14 166.14 156.34 166.26 ;
      RECT 156.86 166.14 157.06 166.26 ;
      RECT 157.58 166.14 157.78 166.26 ;
      RECT 159.02 166.14 159.22 166.26 ;
      RECT 160.46 166.14 160.66 166.26 ;
      RECT 159.74 166.38 159.94 166.5 ;
      RECT 158.3 166.38 158.5 166.5 ;
      RECT 156.14 168.66 156.34 168.78 ;
      RECT 157.94 167.4 158.14 167.52 ;
      RECT 159.02 168.66 159.22 168.78 ;
      RECT 160.46 168.66 160.66 168.78 ;
      RECT 157.58 168.66 157.78 168.78 ;
      RECT 156.86 168.66 157.06 168.78 ;
      RECT 158.3 168.9 158.5 169.02 ;
      RECT 159.74 168.9 159.94 169.02 ;
      RECT 156.86 171.42 157.06 171.54 ;
      RECT 157.58 171.42 157.78 171.54 ;
      RECT 159.74 171.42 159.94 171.54 ;
      RECT 160.46 171.18 160.66 171.3 ;
      RECT 159.02 171.18 159.22 171.3 ;
      RECT 158.3 171.18 158.5 171.3 ;
      RECT 157.94 170.505 158.14 170.625 ;
      RECT 157.94 169.92 158.14 170.04 ;
      RECT 156.14 171.18 156.34 171.3 ;
      RECT 156.86 173.94 157.06 174.06 ;
      RECT 157.58 173.94 157.78 174.06 ;
      RECT 159.02 173.94 159.22 174.06 ;
      RECT 160.46 173.7 160.66 173.82 ;
      RECT 159.74 173.7 159.94 173.82 ;
      RECT 158.3 173.7 158.5 173.82 ;
      RECT 157.94 172.44 158.14 172.56 ;
      RECT 156.14 173.94 156.34 174.06 ;
      RECT 157.94 177.48 158.14 177.6 ;
      RECT 157.58 176.46 157.78 176.58 ;
      RECT 158.3 176.46 158.5 176.58 ;
      RECT 160.46 176.46 160.66 176.58 ;
      RECT 159.74 176.22 159.94 176.34 ;
      RECT 159.02 176.22 159.22 176.34 ;
      RECT 156.86 176.22 157.06 176.34 ;
      RECT 157.94 174.96 158.14 175.08 ;
      RECT 156.14 176.46 156.34 176.58 ;
      RECT 156.86 178.98 157.06 179.1 ;
      RECT 158.3 178.98 158.5 179.1 ;
      RECT 159.74 178.98 159.94 179.1 ;
      RECT 157.58 178.74 157.78 178.86 ;
      RECT 159.02 178.74 159.22 178.86 ;
      RECT 160.46 178.74 160.66 178.86 ;
      RECT 156.14 178.74 156.34 178.86 ;
      RECT 160.46 193.86 160.66 193.98 ;
      RECT 159.02 193.86 159.22 193.98 ;
      RECT 157.94 192.84 158.14 192.96 ;
      RECT 159.74 191.58 159.94 191.7 ;
      RECT 159.02 191.58 159.22 191.7 ;
      RECT 148.22 234.42 148.42 234.54 ;
      RECT 147.5 234.18 147.7 234.3 ;
      RECT 147.5 236.94 147.7 237.06 ;
      RECT 148.94 236.94 149.14 237.06 ;
      RECT 148.22 236.7 148.42 236.82 ;
      RECT 147.5 239.46 147.7 239.58 ;
      RECT 148.94 239.22 149.14 239.34 ;
      RECT 148.22 239.22 148.42 239.34 ;
      RECT 147.5 241.98 147.7 242.1 ;
      RECT 148.22 241.74 148.42 241.86 ;
      RECT 148.94 241.74 149.14 241.86 ;
      RECT 148.94 244.5 149.14 244.62 ;
      RECT 148.22 244.26 148.42 244.38 ;
      RECT 147.5 244.26 147.7 244.38 ;
      RECT 148.22 247.02 148.42 247.14 ;
      RECT 148.94 246.78 149.14 246.9 ;
      RECT 147.5 246.78 147.7 246.9 ;
      RECT 148.22 249.54 148.42 249.66 ;
      RECT 148.94 249.3 149.14 249.42 ;
      RECT 147.5 249.3 147.7 249.42 ;
      RECT 148.22 252.06 148.42 252.18 ;
      RECT 148.94 251.82 149.14 251.94 ;
      RECT 147.5 251.82 147.7 251.94 ;
      RECT 155.06 258.75 155.26 258.87 ;
      RECT 155.42 261.9 155.62 262.02 ;
      RECT 154.7 261.9 154.9 262.02 ;
      RECT 153.26 261.9 153.46 262.02 ;
      RECT 148.22 261.9 148.42 262.02 ;
      RECT 155.06 261.27 155.26 261.39 ;
      RECT 155.06 260.25 155.26 260.37 ;
      RECT 155.42 264.66 155.62 264.78 ;
      RECT 153.98 264.66 154.18 264.78 ;
      RECT 152.54 264.66 152.74 264.78 ;
      RECT 147.5 264.66 147.7 264.78 ;
      RECT 148.94 264.42 149.14 264.54 ;
      RECT 148.22 264.42 148.42 264.54 ;
      RECT 154.7 264.42 154.9 264.54 ;
      RECT 153.26 264.42 153.46 264.54 ;
      RECT 155.06 263.79 155.26 263.91 ;
      RECT 155.06 262.53 155.26 262.65 ;
      RECT 153.98 262.14 154.18 262.26 ;
      RECT 152.54 262.14 152.74 262.26 ;
      RECT 148.94 262.14 149.14 262.26 ;
      RECT 147.5 262.14 147.7 262.26 ;
      RECT 155.42 267.18 155.62 267.3 ;
      RECT 154.7 267.18 154.9 267.3 ;
      RECT 153.98 267.18 154.18 267.3 ;
      RECT 152.54 267.18 152.74 267.3 ;
      RECT 148.94 267.18 149.14 267.3 ;
      RECT 153.26 266.94 153.46 267.06 ;
      RECT 148.22 266.94 148.42 267.06 ;
      RECT 147.5 266.94 147.7 267.06 ;
      RECT 155.06 266.2885 155.26 266.4085 ;
      RECT 155.06 270.09 155.26 270.21 ;
      RECT 154.7 269.7 154.9 269.82 ;
      RECT 153.98 269.7 154.18 269.82 ;
      RECT 153.26 269.7 153.46 269.82 ;
      RECT 152.54 269.7 152.74 269.82 ;
      RECT 148.22 269.7 148.42 269.82 ;
      RECT 147.5 269.7 147.7 269.82 ;
      RECT 155.42 269.46 155.62 269.58 ;
      RECT 148.94 269.46 149.14 269.58 ;
      RECT 155.06 268.83 155.26 268.95 ;
      RECT 155.06 267.81 155.26 267.93 ;
      RECT 155.06 271.35 155.26 271.47 ;
      RECT 155.42 272.22 155.62 272.34 ;
      RECT 153.26 272.22 153.46 272.34 ;
      RECT 148.94 272.22 149.14 272.34 ;
      RECT 147.5 272.22 147.7 272.34 ;
      RECT 154.7 271.98 154.9 272.1 ;
      RECT 153.98 271.98 154.18 272.1 ;
      RECT 152.54 271.98 152.74 272.1 ;
      RECT 148.22 271.98 148.42 272.1 ;
      RECT 153.98 274.74 154.18 274.86 ;
      RECT 148.94 274.74 149.14 274.86 ;
      RECT 152.54 274.74 152.74 274.86 ;
      RECT 153.26 274.5 153.46 274.62 ;
      RECT 148.22 274.5 148.42 274.62 ;
      RECT 147.5 274.5 147.7 274.62 ;
      RECT 155.42 274.5 155.62 274.62 ;
      RECT 154.7 274.5 154.9 274.62 ;
      RECT 147.86 275.3695 148.06 275.4895 ;
      RECT 148.58 275.3695 148.78 275.4895 ;
      RECT 152.9 275.3695 153.1 275.4895 ;
      RECT 153.62 275.3695 153.82 275.4895 ;
      RECT 154.34 275.3695 154.54 275.4895 ;
      RECT 147.5 277.02 147.7 277.14 ;
      RECT 148.94 277.02 149.14 277.14 ;
      RECT 153.26 277.02 153.46 277.14 ;
      RECT 154.7 277.02 154.9 277.14 ;
      RECT 155.42 277.02 155.62 277.14 ;
      RECT 148.22 277.26 148.42 277.38 ;
      RECT 152.54 277.26 152.74 277.38 ;
      RECT 153.98 277.26 154.18 277.38 ;
      RECT 147.86 277.858 148.06 277.978 ;
      RECT 148.58 277.858 148.78 277.978 ;
      RECT 152.9 277.858 153.1 277.978 ;
      RECT 153.62 277.858 153.82 277.978 ;
      RECT 154.34 277.858 154.54 277.978 ;
      RECT 147.86 279.78 148.06 279.9 ;
      RECT 148.58 279.78 148.78 279.9 ;
      RECT 152.9 279.78 153.1 279.9 ;
      RECT 148.94 196.38 149.14 196.5 ;
      RECT 148.22 196.38 148.42 196.5 ;
      RECT 147.5 196.62 147.7 196.74 ;
      RECT 152.54 196.62 152.74 196.74 ;
      RECT 153.98 196.62 154.18 196.74 ;
      RECT 154.7 196.62 154.9 196.74 ;
      RECT 155.06 197.64 155.26 197.76 ;
      RECT 155.42 198.9 155.62 199.02 ;
      RECT 153.26 198.9 153.46 199.02 ;
      RECT 148.94 198.9 149.14 199.02 ;
      RECT 148.22 198.9 148.42 199.02 ;
      RECT 147.5 198.9 147.7 199.02 ;
      RECT 152.54 199.14 152.74 199.26 ;
      RECT 153.98 199.14 154.18 199.26 ;
      RECT 154.7 199.14 154.9 199.26 ;
      RECT 155.06 200.16 155.26 200.28 ;
      RECT 154.7 201.42 154.9 201.54 ;
      RECT 153.26 201.42 153.46 201.54 ;
      RECT 152.54 201.42 152.74 201.54 ;
      RECT 148.94 201.42 149.14 201.54 ;
      RECT 147.5 201.42 147.7 201.54 ;
      RECT 155.42 201.66 155.62 201.78 ;
      RECT 153.98 201.66 154.18 201.78 ;
      RECT 148.22 201.66 148.42 201.78 ;
      RECT 155.42 204.18 155.62 204.3 ;
      RECT 152.54 204.18 152.74 204.3 ;
      RECT 148.22 204.18 148.42 204.3 ;
      RECT 147.5 203.94 147.7 204.06 ;
      RECT 148.94 203.94 149.14 204.06 ;
      RECT 153.26 203.94 153.46 204.06 ;
      RECT 153.98 203.94 154.18 204.06 ;
      RECT 155.06 202.92 155.26 203.04 ;
      RECT 154.7 203.94 154.9 204.06 ;
      RECT 148.22 206.7 148.42 206.82 ;
      RECT 152.54 206.7 152.74 206.82 ;
      RECT 153.98 206.7 154.18 206.82 ;
      RECT 155.42 206.7 155.62 206.82 ;
      RECT 154.7 206.46 154.9 206.58 ;
      RECT 153.26 206.46 153.46 206.58 ;
      RECT 148.94 206.46 149.14 206.58 ;
      RECT 147.5 206.46 147.7 206.58 ;
      RECT 155.06 205.2 155.26 205.32 ;
      RECT 155.42 209.22 155.62 209.34 ;
      RECT 153.26 209.22 153.46 209.34 ;
      RECT 154.7 208.98 154.9 209.1 ;
      RECT 153.98 208.98 154.18 209.1 ;
      RECT 152.54 208.98 152.74 209.1 ;
      RECT 148.94 208.98 149.14 209.1 ;
      RECT 148.22 208.98 148.42 209.1 ;
      RECT 147.5 208.98 147.7 209.1 ;
      RECT 155.06 207.72 155.26 207.84 ;
      RECT 155.42 211.74 155.62 211.86 ;
      RECT 153.26 211.74 153.46 211.86 ;
      RECT 152.54 211.74 152.74 211.86 ;
      RECT 148.94 211.74 149.14 211.86 ;
      RECT 154.7 211.5 154.9 211.62 ;
      RECT 153.98 211.5 154.18 211.62 ;
      RECT 148.22 211.5 148.42 211.62 ;
      RECT 147.5 211.5 147.7 211.62 ;
      RECT 155.06 210.48 155.26 210.6 ;
      RECT 155.06 215.52 155.26 215.64 ;
      RECT 153.98 214.26 154.18 214.38 ;
      RECT 152.54 214.26 152.74 214.38 ;
      RECT 148.94 214.26 149.14 214.38 ;
      RECT 148.22 214.26 148.42 214.38 ;
      RECT 147.5 214.26 147.7 214.38 ;
      RECT 155.42 214.02 155.62 214.14 ;
      RECT 154.7 214.02 154.9 214.14 ;
      RECT 153.26 214.02 153.46 214.14 ;
      RECT 155.06 213 155.26 213.12 ;
      RECT 153.98 216.78 154.18 216.9 ;
      RECT 152.54 216.78 152.74 216.9 ;
      RECT 155.42 216.54 155.62 216.66 ;
      RECT 154.7 216.54 154.9 216.66 ;
      RECT 153.26 216.54 153.46 216.66 ;
      RECT 148.94 216.54 149.14 216.66 ;
      RECT 148.22 216.54 148.42 216.66 ;
      RECT 147.5 216.54 147.7 216.66 ;
      RECT 155.42 219.3 155.62 219.42 ;
      RECT 153.26 219.3 153.46 219.42 ;
      RECT 148.22 219.3 148.42 219.42 ;
      RECT 154.7 219.06 154.9 219.18 ;
      RECT 153.98 219.06 154.18 219.18 ;
      RECT 152.54 219.06 152.74 219.18 ;
      RECT 148.94 219.06 149.14 219.18 ;
      RECT 147.5 219.06 147.7 219.18 ;
      RECT 147.5 223.798 147.7 223.918 ;
      RECT 148.22 223.798 148.42 223.918 ;
      RECT 148.94 223.798 149.14 223.918 ;
      RECT 152.54 223.798 152.74 223.918 ;
      RECT 153.98 223.798 154.18 223.918 ;
      RECT 155.42 223.798 155.62 223.918 ;
      RECT 153.26 223.558 153.46 223.678 ;
      RECT 154.7 223.558 154.9 223.678 ;
      RECT 155.06 223.08 155.26 223.2 ;
      RECT 148.22 229.14 148.42 229.26 ;
      RECT 148.94 229.14 149.14 229.26 ;
      RECT 148.94 231.9 149.14 232.02 ;
      RECT 147.5 231.9 147.7 232.02 ;
      RECT 148.22 231.66 148.42 231.78 ;
      RECT 147.5 229.38 147.7 229.5 ;
      RECT 148.94 234.42 149.14 234.54 ;
      RECT 143.9 325.9425 144.1 326.0625 ;
      RECT 143.18 325.9425 143.38 326.0625 ;
      RECT 142.46 325.9425 142.66 326.0625 ;
      RECT 141.74 325.9425 141.94 326.0625 ;
      RECT 141.02 325.9425 141.22 326.0625 ;
      RECT 146.78 325.9425 146.98 326.0625 ;
      RECT 146.06 325.9425 146.26 326.0625 ;
      RECT 145.34 325.9425 145.54 326.0625 ;
      RECT 144.62 325.9425 144.82 326.0625 ;
      RECT 146.42 348.339 146.62 348.459 ;
      RECT 143.54 348.339 143.74 348.459 ;
      RECT 155.42 118.324 155.62 118.444 ;
      RECT 153.26 118.324 153.46 118.444 ;
      RECT 148.22 118.324 148.42 118.444 ;
      RECT 147.5 118.324 147.7 118.444 ;
      RECT 148.94 118.084 149.14 118.204 ;
      RECT 152.54 118.084 152.74 118.204 ;
      RECT 153.98 118.084 154.18 118.204 ;
      RECT 154.7 118.084 154.9 118.204 ;
      RECT 155.06 154.8 155.26 154.92 ;
      RECT 153.98 156.3 154.18 156.42 ;
      RECT 153.26 156.3 153.46 156.42 ;
      RECT 148.22 156.3 148.42 156.42 ;
      RECT 147.5 156.06 147.7 156.18 ;
      RECT 148.94 156.06 149.14 156.18 ;
      RECT 152.54 156.06 152.74 156.18 ;
      RECT 154.7 156.06 154.9 156.18 ;
      RECT 155.42 156.06 155.62 156.18 ;
      RECT 147.5 166.38 147.7 166.5 ;
      RECT 152.54 166.38 152.74 166.5 ;
      RECT 153.98 166.38 154.18 166.5 ;
      RECT 155.42 166.38 155.62 166.5 ;
      RECT 154.7 166.14 154.9 166.26 ;
      RECT 153.26 166.14 153.46 166.26 ;
      RECT 148.94 166.14 149.14 166.26 ;
      RECT 148.22 166.14 148.42 166.26 ;
      RECT 155.42 168.9 155.62 169.02 ;
      RECT 153.98 168.9 154.18 169.02 ;
      RECT 152.54 168.9 152.74 169.02 ;
      RECT 147.5 168.66 147.7 168.78 ;
      RECT 148.22 168.66 148.42 168.78 ;
      RECT 148.94 168.66 149.14 168.78 ;
      RECT 153.26 168.66 153.46 168.78 ;
      RECT 154.7 168.66 154.9 168.78 ;
      RECT 155.06 167.4 155.26 167.52 ;
      RECT 155.06 169.92 155.26 170.04 ;
      RECT 155.06 170.505 155.26 170.625 ;
      RECT 148.94 171.18 149.14 171.3 ;
      RECT 153.98 171.18 154.18 171.3 ;
      RECT 152.54 171.18 152.74 171.3 ;
      RECT 148.22 171.18 148.42 171.3 ;
      RECT 155.42 171.42 155.62 171.54 ;
      RECT 154.7 171.42 154.9 171.54 ;
      RECT 153.26 171.42 153.46 171.54 ;
      RECT 147.5 171.42 147.7 171.54 ;
      RECT 155.06 172.68 155.26 172.8 ;
      RECT 148.22 173.7 148.42 173.82 ;
      RECT 148.94 173.7 149.14 173.82 ;
      RECT 152.54 173.7 152.74 173.82 ;
      RECT 153.26 173.7 153.46 173.82 ;
      RECT 153.98 173.7 154.18 173.82 ;
      RECT 155.42 173.7 155.62 173.82 ;
      RECT 154.7 173.94 154.9 174.06 ;
      RECT 147.5 173.94 147.7 174.06 ;
      RECT 155.06 175.2 155.26 175.32 ;
      RECT 147.5 176.22 147.7 176.34 ;
      RECT 148.22 176.22 148.42 176.34 ;
      RECT 148.94 176.22 149.14 176.34 ;
      RECT 152.54 176.22 152.74 176.34 ;
      RECT 153.98 176.22 154.18 176.34 ;
      RECT 155.42 176.22 155.62 176.34 ;
      RECT 154.7 176.46 154.9 176.58 ;
      RECT 153.26 176.46 153.46 176.58 ;
      RECT 155.06 177.72 155.26 177.84 ;
      RECT 154.7 178.74 154.9 178.86 ;
      RECT 153.26 178.74 153.46 178.86 ;
      RECT 148.94 178.74 149.14 178.86 ;
      RECT 148.22 178.74 148.42 178.86 ;
      RECT 155.42 178.98 155.62 179.1 ;
      RECT 153.98 178.98 154.18 179.1 ;
      RECT 152.54 178.98 152.74 179.1 ;
      RECT 147.5 178.98 147.7 179.1 ;
      RECT 147.5 191.34 147.7 191.46 ;
      RECT 148.94 191.34 149.14 191.46 ;
      RECT 152.54 191.34 152.74 191.46 ;
      RECT 153.98 191.34 154.18 191.46 ;
      RECT 154.7 191.34 154.9 191.46 ;
      RECT 148.22 191.58 148.42 191.7 ;
      RECT 153.26 191.58 153.46 191.7 ;
      RECT 155.42 191.58 155.62 191.7 ;
      RECT 155.06 192.6 155.26 192.72 ;
      RECT 148.22 193.86 148.42 193.98 ;
      RECT 148.94 193.86 149.14 193.98 ;
      RECT 153.98 193.86 154.18 193.98 ;
      RECT 155.42 193.86 155.62 193.98 ;
      RECT 147.5 194.1 147.7 194.22 ;
      RECT 152.54 194.1 152.74 194.22 ;
      RECT 153.26 194.1 153.46 194.22 ;
      RECT 154.7 194.1 154.9 194.22 ;
      RECT 155.06 195.12 155.26 195.24 ;
      RECT 153.26 196.38 153.46 196.5 ;
      RECT 155.42 196.38 155.62 196.5 ;
      RECT 142.46 267.18 142.66 267.3 ;
      RECT 141.02 267.18 141.22 267.3 ;
      RECT 145.34 266.94 145.54 267.06 ;
      RECT 144.62 266.94 144.82 267.06 ;
      RECT 143.18 266.94 143.38 267.06 ;
      RECT 141.74 266.94 141.94 267.06 ;
      RECT 146.42 266.2885 146.62 266.4085 ;
      RECT 143.54 266.2885 143.74 266.4085 ;
      RECT 143.54 270.09 143.74 270.21 ;
      RECT 145.34 269.7 145.54 269.82 ;
      RECT 143.9 269.7 144.1 269.82 ;
      RECT 143.18 269.7 143.38 269.82 ;
      RECT 141.02 269.7 141.22 269.82 ;
      RECT 146.78 269.46 146.98 269.58 ;
      RECT 146.06 269.46 146.26 269.58 ;
      RECT 144.62 269.46 144.82 269.58 ;
      RECT 142.46 269.46 142.66 269.58 ;
      RECT 141.74 269.46 141.94 269.58 ;
      RECT 146.42 269.07 146.62 269.19 ;
      RECT 143.54 269.07 143.74 269.19 ;
      RECT 146.42 267.81 146.62 267.93 ;
      RECT 143.54 267.81 143.74 267.93 ;
      RECT 146.42 271.35 146.62 271.47 ;
      RECT 143.54 271.35 143.74 271.47 ;
      RECT 146.42 270.33 146.62 270.45 ;
      RECT 143.9 272.22 144.1 272.34 ;
      RECT 142.46 272.22 142.66 272.34 ;
      RECT 141.74 272.22 141.94 272.34 ;
      RECT 141.02 272.22 141.22 272.34 ;
      RECT 146.78 272.22 146.98 272.34 ;
      RECT 145.34 272.22 145.54 272.34 ;
      RECT 146.06 271.98 146.26 272.1 ;
      RECT 144.62 271.98 144.82 272.1 ;
      RECT 143.18 271.98 143.38 272.1 ;
      RECT 142.82 275.1295 143.02 275.2495 ;
      RECT 142.1 275.1295 142.3 275.2495 ;
      RECT 141.38 275.1295 141.58 275.2495 ;
      RECT 144.62 274.74 144.82 274.86 ;
      RECT 146.06 274.74 146.26 274.86 ;
      RECT 146.78 274.74 146.98 274.86 ;
      RECT 143.9 274.74 144.1 274.86 ;
      RECT 143.18 274.74 143.38 274.86 ;
      RECT 141.74 274.74 141.94 274.86 ;
      RECT 145.34 274.5 145.54 274.62 ;
      RECT 142.46 274.5 142.66 274.62 ;
      RECT 141.02 274.5 141.22 274.62 ;
      RECT 144.26 275.3695 144.46 275.4895 ;
      RECT 144.98 275.3695 145.18 275.4895 ;
      RECT 145.7 275.3695 145.9 275.4895 ;
      RECT 147.14 275.3695 147.34 275.4895 ;
      RECT 141.02 277.02 141.22 277.14 ;
      RECT 143.18 277.02 143.38 277.14 ;
      RECT 145.34 277.02 145.54 277.14 ;
      RECT 146.06 277.02 146.26 277.14 ;
      RECT 141.74 277.26 141.94 277.38 ;
      RECT 142.46 277.26 142.66 277.38 ;
      RECT 143.9 277.26 144.1 277.38 ;
      RECT 144.62 277.26 144.82 277.38 ;
      RECT 146.78 277.26 146.98 277.38 ;
      RECT 141.38 277.618 141.58 277.738 ;
      RECT 142.82 277.618 143.02 277.738 ;
      RECT 144.26 277.618 144.46 277.738 ;
      RECT 144.98 277.618 145.18 277.738 ;
      RECT 142.1 277.858 142.3 277.978 ;
      RECT 145.7 277.858 145.9 277.978 ;
      RECT 147.14 277.858 147.34 277.978 ;
      RECT 142.1 279.54 142.3 279.66 ;
      RECT 144.98 279.54 145.18 279.66 ;
      RECT 145.7 279.54 145.9 279.66 ;
      RECT 147.14 279.54 147.34 279.66 ;
      RECT 141.38 279.78 141.58 279.9 ;
      RECT 144.26 279.78 144.46 279.9 ;
      RECT 142.82 279.78 143.02 279.9 ;
      RECT 141.38 282.06 141.58 282.18 ;
      RECT 142.82 282.06 143.02 282.18 ;
      RECT 144.98 282.06 145.18 282.18 ;
      RECT 147.14 282.06 147.34 282.18 ;
      RECT 142.1 282.3 142.3 282.42 ;
      RECT 144.26 282.3 144.46 282.42 ;
      RECT 145.7 282.3 145.9 282.42 ;
      RECT 141.02 285.8245 141.22 285.9445 ;
      RECT 141.74 285.8245 141.94 285.9445 ;
      RECT 142.46 285.8245 142.66 285.9445 ;
      RECT 143.18 285.8245 143.38 285.9445 ;
      RECT 143.9 285.8245 144.1 285.9445 ;
      RECT 144.62 285.8245 144.82 285.9445 ;
      RECT 145.34 285.8245 145.54 285.9445 ;
      RECT 146.06 285.8245 146.26 285.9445 ;
      RECT 146.78 285.8245 146.98 285.9445 ;
      RECT 143.54 305.625 143.74 305.745 ;
      RECT 146.42 305.625 146.62 305.745 ;
      RECT 143.18 306.041 143.38 306.161 ;
      RECT 143.9 306.041 144.1 306.161 ;
      RECT 144.62 306.041 144.82 306.161 ;
      RECT 145.34 306.041 145.54 306.161 ;
      RECT 146.06 306.041 146.26 306.161 ;
      RECT 146.78 306.041 146.98 306.161 ;
      RECT 141.02 306.041 141.22 306.161 ;
      RECT 141.74 306.041 141.94 306.161 ;
      RECT 142.46 306.041 142.66 306.161 ;
      RECT 146.42 323.3835 146.62 323.5035 ;
      RECT 143.54 323.3835 143.74 323.5035 ;
      RECT 143.9 236.7 144.1 236.82 ;
      RECT 143.18 236.7 143.38 236.82 ;
      RECT 141.74 236.7 141.94 236.82 ;
      RECT 143.54 235.68 143.74 235.8 ;
      RECT 146.42 235.44 146.62 235.56 ;
      RECT 146.78 239.46 146.98 239.58 ;
      RECT 144.62 239.46 144.82 239.58 ;
      RECT 142.46 239.46 142.66 239.58 ;
      RECT 141.02 239.46 141.22 239.58 ;
      RECT 146.06 239.22 146.26 239.34 ;
      RECT 145.34 239.22 145.54 239.34 ;
      RECT 143.9 239.22 144.1 239.34 ;
      RECT 143.18 239.22 143.38 239.34 ;
      RECT 141.74 239.22 141.94 239.34 ;
      RECT 143.54 238.2 143.74 238.32 ;
      RECT 146.42 237.96 146.62 238.08 ;
      RECT 143.54 243 143.74 243.12 ;
      RECT 141.02 241.98 141.22 242.1 ;
      RECT 142.46 241.98 142.66 242.1 ;
      RECT 143.9 241.98 144.1 242.1 ;
      RECT 144.62 241.98 144.82 242.1 ;
      RECT 145.34 241.98 145.54 242.1 ;
      RECT 141.74 241.74 141.94 241.86 ;
      RECT 143.18 241.74 143.38 241.86 ;
      RECT 146.06 241.74 146.26 241.86 ;
      RECT 146.78 241.74 146.98 241.86 ;
      RECT 143.54 240.72 143.74 240.84 ;
      RECT 146.42 240.48 146.62 240.6 ;
      RECT 146.42 245.52 146.62 245.64 ;
      RECT 146.78 244.5 146.98 244.62 ;
      RECT 141.02 244.5 141.22 244.62 ;
      RECT 143.18 244.5 143.38 244.62 ;
      RECT 143.9 244.5 144.1 244.62 ;
      RECT 145.34 244.5 145.54 244.62 ;
      RECT 146.06 244.26 146.26 244.38 ;
      RECT 144.62 244.26 144.82 244.38 ;
      RECT 142.46 244.26 142.66 244.38 ;
      RECT 141.74 244.26 141.94 244.38 ;
      RECT 146.42 243.24 146.62 243.36 ;
      RECT 143.54 248.28 143.74 248.4 ;
      RECT 146.42 248.04 146.62 248.16 ;
      RECT 146.78 247.02 146.98 247.14 ;
      RECT 145.34 247.02 145.54 247.14 ;
      RECT 143.9 247.02 144.1 247.14 ;
      RECT 144.62 246.78 144.82 246.9 ;
      RECT 143.18 246.78 143.38 246.9 ;
      RECT 142.46 246.78 142.66 246.9 ;
      RECT 141.74 246.78 141.94 246.9 ;
      RECT 146.06 246.78 146.26 246.9 ;
      RECT 141.02 246.78 141.22 246.9 ;
      RECT 143.54 245.76 143.74 245.88 ;
      RECT 143.54 250.8 143.74 250.92 ;
      RECT 146.42 250.56 146.62 250.68 ;
      RECT 144.62 249.54 144.82 249.66 ;
      RECT 142.46 249.54 142.66 249.66 ;
      RECT 141.74 249.54 141.94 249.66 ;
      RECT 146.78 249.54 146.98 249.66 ;
      RECT 146.06 249.3 146.26 249.42 ;
      RECT 145.34 249.3 145.54 249.42 ;
      RECT 143.9 249.3 144.1 249.42 ;
      RECT 143.18 249.3 143.38 249.42 ;
      RECT 141.02 249.3 141.22 249.42 ;
      RECT 146.78 252.06 146.98 252.18 ;
      RECT 145.34 252.06 145.54 252.18 ;
      RECT 143.9 252.06 144.1 252.18 ;
      RECT 146.06 251.82 146.26 251.94 ;
      RECT 144.62 251.82 144.82 251.94 ;
      RECT 143.18 251.82 143.38 251.94 ;
      RECT 142.46 251.82 142.66 251.94 ;
      RECT 141.74 251.82 141.94 251.94 ;
      RECT 141.02 251.82 141.22 251.94 ;
      RECT 146.42 258.75 146.62 258.87 ;
      RECT 143.54 258.75 143.74 258.87 ;
      RECT 146.78 261.9 146.98 262.02 ;
      RECT 145.34 261.9 145.54 262.02 ;
      RECT 144.62 261.9 144.82 262.02 ;
      RECT 141.74 261.9 141.94 262.02 ;
      RECT 146.42 261.51 146.62 261.63 ;
      RECT 143.54 261.27 143.74 261.39 ;
      RECT 146.42 260.01 146.62 260.13 ;
      RECT 143.54 260.01 143.74 260.13 ;
      RECT 145.34 264.66 145.54 264.78 ;
      RECT 144.62 264.66 144.82 264.78 ;
      RECT 143.18 264.66 143.38 264.78 ;
      RECT 142.46 264.66 142.66 264.78 ;
      RECT 141.02 264.66 141.22 264.78 ;
      RECT 146.78 264.42 146.98 264.54 ;
      RECT 146.06 264.42 146.26 264.54 ;
      RECT 143.9 264.42 144.1 264.54 ;
      RECT 141.74 264.42 141.94 264.54 ;
      RECT 146.42 263.79 146.62 263.91 ;
      RECT 143.54 263.79 143.74 263.91 ;
      RECT 146.42 262.53 146.62 262.65 ;
      RECT 143.54 262.53 143.74 262.65 ;
      RECT 146.06 262.14 146.26 262.26 ;
      RECT 143.9 262.14 144.1 262.26 ;
      RECT 143.18 262.14 143.38 262.26 ;
      RECT 142.46 262.14 142.66 262.26 ;
      RECT 141.02 262.14 141.22 262.26 ;
      RECT 146.78 267.18 146.98 267.3 ;
      RECT 146.06 267.18 146.26 267.3 ;
      RECT 143.9 267.18 144.1 267.3 ;
      RECT 146.78 209.22 146.98 209.34 ;
      RECT 145.34 209.22 145.54 209.34 ;
      RECT 143.9 209.22 144.1 209.34 ;
      RECT 143.18 209.22 143.38 209.34 ;
      RECT 141.74 209.22 141.94 209.34 ;
      RECT 146.06 208.98 146.26 209.1 ;
      RECT 144.62 208.98 144.82 209.1 ;
      RECT 142.46 208.98 142.66 209.1 ;
      RECT 141.02 208.98 141.22 209.1 ;
      RECT 143.54 207.96 143.74 208.08 ;
      RECT 146.42 207.72 146.62 207.84 ;
      RECT 146.42 212.76 146.62 212.88 ;
      RECT 146.78 211.74 146.98 211.86 ;
      RECT 146.06 211.74 146.26 211.86 ;
      RECT 144.62 211.74 144.82 211.86 ;
      RECT 143.18 211.74 143.38 211.86 ;
      RECT 141.74 211.74 141.94 211.86 ;
      RECT 145.34 211.5 145.54 211.62 ;
      RECT 143.9 211.5 144.1 211.62 ;
      RECT 142.46 211.5 142.66 211.62 ;
      RECT 141.02 211.5 141.22 211.62 ;
      RECT 143.54 210.48 143.74 210.6 ;
      RECT 143.54 215.52 143.74 215.64 ;
      RECT 146.42 215.28 146.62 215.4 ;
      RECT 146.06 214.26 146.26 214.38 ;
      RECT 144.62 214.26 144.82 214.38 ;
      RECT 143.18 214.26 143.38 214.38 ;
      RECT 141.74 214.26 141.94 214.38 ;
      RECT 146.78 214.02 146.98 214.14 ;
      RECT 145.34 214.02 145.54 214.14 ;
      RECT 143.9 214.02 144.1 214.14 ;
      RECT 142.46 214.02 142.66 214.14 ;
      RECT 141.02 214.02 141.22 214.14 ;
      RECT 143.54 213 143.74 213.12 ;
      RECT 146.78 216.78 146.98 216.9 ;
      RECT 146.06 216.78 146.26 216.9 ;
      RECT 145.34 216.78 145.54 216.9 ;
      RECT 144.62 216.78 144.82 216.9 ;
      RECT 143.9 216.78 144.1 216.9 ;
      RECT 143.18 216.78 143.38 216.9 ;
      RECT 141.02 216.78 141.22 216.9 ;
      RECT 142.46 216.54 142.66 216.66 ;
      RECT 141.74 216.54 141.94 216.66 ;
      RECT 146.78 219.3 146.98 219.42 ;
      RECT 146.06 219.3 146.26 219.42 ;
      RECT 144.62 219.3 144.82 219.42 ;
      RECT 143.9 219.3 144.1 219.42 ;
      RECT 143.18 219.3 143.38 219.42 ;
      RECT 141.74 219.3 141.94 219.42 ;
      RECT 145.34 219.06 145.54 219.18 ;
      RECT 142.46 219.06 142.66 219.18 ;
      RECT 141.02 219.06 141.22 219.18 ;
      RECT 141.02 223.798 141.22 223.918 ;
      RECT 143.18 223.798 143.38 223.918 ;
      RECT 144.62 223.798 144.82 223.918 ;
      RECT 145.34 223.798 145.54 223.918 ;
      RECT 141.74 223.558 141.94 223.678 ;
      RECT 142.46 223.558 142.66 223.678 ;
      RECT 143.9 223.558 144.1 223.678 ;
      RECT 146.06 223.558 146.26 223.678 ;
      RECT 146.78 223.558 146.98 223.678 ;
      RECT 143.54 223.08 143.74 223.2 ;
      RECT 146.42 222.84 146.62 222.96 ;
      RECT 141.02 229.14 141.22 229.26 ;
      RECT 143.18 229.14 143.38 229.26 ;
      RECT 143.9 229.14 144.1 229.26 ;
      RECT 145.34 229.14 145.54 229.26 ;
      RECT 146.78 229.14 146.98 229.26 ;
      RECT 143.54 228.12 143.74 228.24 ;
      RECT 146.42 227.88 146.62 228 ;
      RECT 146.78 231.9 146.98 232.02 ;
      RECT 145.34 231.9 145.54 232.02 ;
      RECT 143.9 231.9 144.1 232.02 ;
      RECT 141.02 231.9 141.22 232.02 ;
      RECT 146.06 231.66 146.26 231.78 ;
      RECT 144.62 231.66 144.82 231.78 ;
      RECT 143.18 231.66 143.38 231.78 ;
      RECT 142.46 231.66 142.66 231.78 ;
      RECT 141.74 231.66 141.94 231.78 ;
      RECT 143.54 230.64 143.74 230.76 ;
      RECT 146.42 230.4 146.62 230.52 ;
      RECT 141.74 229.38 141.94 229.5 ;
      RECT 142.46 229.38 142.66 229.5 ;
      RECT 144.62 229.38 144.82 229.5 ;
      RECT 146.06 229.38 146.26 229.5 ;
      RECT 146.78 234.42 146.98 234.54 ;
      RECT 145.34 234.42 145.54 234.54 ;
      RECT 143.18 234.42 143.38 234.54 ;
      RECT 142.46 234.42 142.66 234.54 ;
      RECT 141.02 234.42 141.22 234.54 ;
      RECT 141.74 234.18 141.94 234.3 ;
      RECT 143.9 234.18 144.1 234.3 ;
      RECT 144.62 234.18 144.82 234.3 ;
      RECT 146.06 234.18 146.26 234.3 ;
      RECT 143.54 233.16 143.74 233.28 ;
      RECT 146.42 232.92 146.62 233.04 ;
      RECT 141.02 236.94 141.22 237.06 ;
      RECT 142.46 236.94 142.66 237.06 ;
      RECT 146.78 236.7 146.98 236.82 ;
      RECT 146.06 236.7 146.26 236.82 ;
      RECT 145.34 236.7 145.54 236.82 ;
      RECT 144.62 236.7 144.82 236.82 ;
      RECT 142.46 173.7 142.66 173.82 ;
      RECT 141.74 173.7 141.94 173.82 ;
      RECT 146.42 172.44 146.62 172.56 ;
      RECT 143.54 172.68 143.74 172.8 ;
      RECT 146.42 177.48 146.62 177.6 ;
      RECT 141.74 176.46 141.94 176.58 ;
      RECT 142.46 176.46 142.66 176.58 ;
      RECT 143.9 176.46 144.1 176.58 ;
      RECT 145.34 176.46 145.54 176.58 ;
      RECT 146.78 176.46 146.98 176.58 ;
      RECT 146.06 176.22 146.26 176.34 ;
      RECT 144.62 176.22 144.82 176.34 ;
      RECT 143.18 176.22 143.38 176.34 ;
      RECT 141.02 176.22 141.22 176.34 ;
      RECT 143.54 175.2 143.74 175.32 ;
      RECT 146.42 174.96 146.62 175.08 ;
      RECT 141.02 178.98 141.22 179.1 ;
      RECT 142.46 178.98 142.66 179.1 ;
      RECT 143.18 178.98 143.38 179.1 ;
      RECT 143.9 178.98 144.1 179.1 ;
      RECT 146.78 178.98 146.98 179.1 ;
      RECT 141.74 178.74 141.94 178.86 ;
      RECT 144.62 178.74 144.82 178.86 ;
      RECT 145.34 178.74 145.54 178.86 ;
      RECT 146.06 178.74 146.26 178.86 ;
      RECT 143.54 177.72 143.74 177.84 ;
      RECT 146.78 193.86 146.98 193.98 ;
      RECT 145.34 193.86 145.54 193.98 ;
      RECT 143.9 193.86 144.1 193.98 ;
      RECT 143.18 193.86 143.38 193.98 ;
      RECT 141.74 193.86 141.94 193.98 ;
      RECT 143.54 192.6 143.74 192.72 ;
      RECT 146.42 192.6 146.62 192.72 ;
      RECT 144.62 191.58 144.82 191.7 ;
      RECT 142.46 191.58 142.66 191.7 ;
      RECT 141.02 191.58 141.22 191.7 ;
      RECT 146.78 191.34 146.98 191.46 ;
      RECT 146.06 191.34 146.26 191.46 ;
      RECT 145.34 191.34 145.54 191.46 ;
      RECT 143.9 191.34 144.1 191.46 ;
      RECT 143.18 191.34 143.38 191.46 ;
      RECT 141.74 191.34 141.94 191.46 ;
      RECT 141.74 196.38 141.94 196.5 ;
      RECT 143.18 196.38 143.38 196.5 ;
      RECT 143.9 196.38 144.1 196.5 ;
      RECT 145.34 196.38 145.54 196.5 ;
      RECT 146.78 196.38 146.98 196.5 ;
      RECT 146.42 195.36 146.62 195.48 ;
      RECT 143.54 195.36 143.74 195.48 ;
      RECT 146.06 194.1 146.26 194.22 ;
      RECT 144.62 194.1 144.82 194.22 ;
      RECT 142.46 194.1 142.66 194.22 ;
      RECT 141.02 194.1 141.22 194.22 ;
      RECT 146.78 199.14 146.98 199.26 ;
      RECT 145.34 199.14 145.54 199.26 ;
      RECT 143.9 199.14 144.1 199.26 ;
      RECT 143.18 199.14 143.38 199.26 ;
      RECT 141.02 199.14 141.22 199.26 ;
      RECT 141.74 198.9 141.94 199.02 ;
      RECT 142.46 198.9 142.66 199.02 ;
      RECT 144.62 198.9 144.82 199.02 ;
      RECT 146.06 198.9 146.26 199.02 ;
      RECT 143.54 197.88 143.74 198 ;
      RECT 146.42 197.64 146.62 197.76 ;
      RECT 146.06 196.62 146.26 196.74 ;
      RECT 144.62 196.62 144.82 196.74 ;
      RECT 142.46 196.62 142.66 196.74 ;
      RECT 141.02 196.62 141.22 196.74 ;
      RECT 142.46 201.66 142.66 201.78 ;
      RECT 143.9 201.66 144.1 201.78 ;
      RECT 145.34 201.66 145.54 201.78 ;
      RECT 146.78 201.66 146.98 201.78 ;
      RECT 141.02 201.42 141.22 201.54 ;
      RECT 141.74 201.42 141.94 201.54 ;
      RECT 143.18 201.42 143.38 201.54 ;
      RECT 144.62 201.42 144.82 201.54 ;
      RECT 146.06 201.42 146.26 201.54 ;
      RECT 143.54 200.4 143.74 200.52 ;
      RECT 146.42 200.16 146.62 200.28 ;
      RECT 146.78 204.18 146.98 204.3 ;
      RECT 145.34 204.18 145.54 204.3 ;
      RECT 143.9 204.18 144.1 204.3 ;
      RECT 143.18 204.18 143.38 204.3 ;
      RECT 141.74 204.18 141.94 204.3 ;
      RECT 142.46 203.94 142.66 204.06 ;
      RECT 144.62 203.94 144.82 204.06 ;
      RECT 146.06 203.94 146.26 204.06 ;
      RECT 141.02 203.94 141.22 204.06 ;
      RECT 143.54 202.92 143.74 203.04 ;
      RECT 146.42 202.68 146.62 202.8 ;
      RECT 141.74 206.7 141.94 206.82 ;
      RECT 143.18 206.7 143.38 206.82 ;
      RECT 144.62 206.7 144.82 206.82 ;
      RECT 145.34 206.7 145.54 206.82 ;
      RECT 146.78 206.7 146.98 206.82 ;
      RECT 146.06 206.46 146.26 206.58 ;
      RECT 143.9 206.46 144.1 206.58 ;
      RECT 142.46 206.46 142.66 206.58 ;
      RECT 141.02 206.46 141.22 206.58 ;
      RECT 143.54 205.44 143.74 205.56 ;
      RECT 146.42 205.2 146.62 205.32 ;
      RECT 146.42 210.24 146.62 210.36 ;
      RECT 132.02 271.35 132.22 271.47 ;
      RECT 131.66 270.96 131.86 271.08 ;
      RECT 133.82 270.72 134.02 270.84 ;
      RECT 133.1 270.72 133.3 270.84 ;
      RECT 132.38 270.72 132.58 270.84 ;
      RECT 134.18 270.33 134.38 270.45 ;
      RECT 133.46 270.33 133.66 270.45 ;
      RECT 131.3 270.33 131.5 270.45 ;
      RECT 135.26 273.24 135.46 273.36 ;
      RECT 134.54 273.24 134.74 273.36 ;
      RECT 135.26 275.76 135.46 275.88 ;
      RECT 132.38 273.24 132.58 273.36 ;
      RECT 133.1 273.24 133.3 273.36 ;
      RECT 131.66 273.48 131.86 273.6 ;
      RECT 133.82 273.48 134.02 273.6 ;
      RECT 132.38 275.76 132.58 275.88 ;
      RECT 133.82 275.76 134.02 275.88 ;
      RECT 134.54 276 134.74 276.12 ;
      RECT 135.26 278.28 135.46 278.4 ;
      RECT 131.66 276 131.86 276.12 ;
      RECT 133.1 276 133.3 276.12 ;
      RECT 132.38 278.28 132.58 278.4 ;
      RECT 133.82 278.28 134.02 278.4 ;
      RECT 134.54 278.52 134.74 278.64 ;
      RECT 133.1 278.52 133.3 278.64 ;
      RECT 131.66 278.52 131.86 278.64 ;
      RECT 134.18 305.625 134.38 305.745 ;
      RECT 133.46 305.625 133.66 305.745 ;
      RECT 132.74 305.625 132.94 305.745 ;
      RECT 132.02 305.625 132.22 305.745 ;
      RECT 131.3 305.625 131.5 305.745 ;
      RECT 134.9 305.625 135.1 305.745 ;
      RECT 134.18 323.3835 134.38 323.5035 ;
      RECT 133.46 323.3835 133.66 323.5035 ;
      RECT 132.74 323.3835 132.94 323.5035 ;
      RECT 132.02 323.3835 132.22 323.5035 ;
      RECT 131.3 323.3835 131.5 323.5035 ;
      RECT 134.9 323.3835 135.1 323.5035 ;
      RECT 134.18 348.339 134.38 348.459 ;
      RECT 133.46 348.339 133.66 348.459 ;
      RECT 132.74 348.339 132.94 348.459 ;
      RECT 132.02 348.339 132.22 348.459 ;
      RECT 131.3 348.339 131.5 348.459 ;
      RECT 134.9 348.339 135.1 348.459 ;
      RECT 146.78 118.324 146.98 118.444 ;
      RECT 144.62 118.324 144.82 118.444 ;
      RECT 143.9 118.324 144.1 118.444 ;
      RECT 141.74 118.324 141.94 118.444 ;
      RECT 141.02 118.084 141.22 118.204 ;
      RECT 142.46 118.084 142.66 118.204 ;
      RECT 143.18 118.084 143.38 118.204 ;
      RECT 145.34 118.084 145.54 118.204 ;
      RECT 146.06 118.084 146.26 118.204 ;
      RECT 143.54 155.04 143.74 155.16 ;
      RECT 146.42 154.8 146.62 154.92 ;
      RECT 146.78 156.3 146.98 156.42 ;
      RECT 145.34 156.3 145.54 156.42 ;
      RECT 144.62 156.3 144.82 156.42 ;
      RECT 143.18 156.3 143.38 156.42 ;
      RECT 142.46 156.3 142.66 156.42 ;
      RECT 141.02 156.3 141.22 156.42 ;
      RECT 146.06 156.06 146.26 156.18 ;
      RECT 143.9 156.06 144.1 156.18 ;
      RECT 141.74 156.06 141.94 156.18 ;
      RECT 143.9 166.38 144.1 166.5 ;
      RECT 145.34 166.38 145.54 166.5 ;
      RECT 146.78 166.38 146.98 166.5 ;
      RECT 141.02 166.14 141.22 166.26 ;
      RECT 141.74 166.14 141.94 166.26 ;
      RECT 142.46 166.14 142.66 166.26 ;
      RECT 143.18 166.14 143.38 166.26 ;
      RECT 144.62 166.14 144.82 166.26 ;
      RECT 146.06 166.14 146.26 166.26 ;
      RECT 146.78 168.9 146.98 169.02 ;
      RECT 146.06 168.9 146.26 169.02 ;
      RECT 143.9 168.9 144.1 169.02 ;
      RECT 142.46 168.9 142.66 169.02 ;
      RECT 141.02 168.9 141.22 169.02 ;
      RECT 141.74 168.66 141.94 168.78 ;
      RECT 143.18 168.66 143.38 168.78 ;
      RECT 144.62 168.66 144.82 168.78 ;
      RECT 145.34 168.66 145.54 168.78 ;
      RECT 143.54 167.64 143.74 167.76 ;
      RECT 146.42 167.4 146.62 167.52 ;
      RECT 146.42 169.92 146.62 170.04 ;
      RECT 143.54 170.16 143.74 170.28 ;
      RECT 141.74 171.18 141.94 171.3 ;
      RECT 143.18 171.18 143.38 171.3 ;
      RECT 144.62 171.18 144.82 171.3 ;
      RECT 145.34 171.18 145.54 171.3 ;
      RECT 146.78 171.18 146.98 171.3 ;
      RECT 146.06 171.42 146.26 171.54 ;
      RECT 143.9 171.42 144.1 171.54 ;
      RECT 142.46 171.42 142.66 171.54 ;
      RECT 141.02 171.42 141.22 171.54 ;
      RECT 146.78 173.94 146.98 174.06 ;
      RECT 145.34 173.94 145.54 174.06 ;
      RECT 143.9 173.94 144.1 174.06 ;
      RECT 141.02 173.94 141.22 174.06 ;
      RECT 146.06 173.7 146.26 173.82 ;
      RECT 144.62 173.7 144.82 173.82 ;
      RECT 143.18 173.7 143.38 173.82 ;
      RECT 132.02 213 132.22 213.12 ;
      RECT 134.9 215.28 135.1 215.4 ;
      RECT 134.9 222.84 135.1 222.96 ;
      RECT 134.54 222.122 134.74 222.242 ;
      RECT 135.26 222.122 135.46 222.242 ;
      RECT 132.02 223.08 132.22 223.2 ;
      RECT 134.18 223.08 134.38 223.2 ;
      RECT 131.3 222.84 131.5 222.96 ;
      RECT 132.74 222.84 132.94 222.96 ;
      RECT 133.46 222.84 133.66 222.96 ;
      RECT 131.66 222.362 131.86 222.482 ;
      RECT 133.1 222.362 133.3 222.482 ;
      RECT 133.82 222.362 134.02 222.482 ;
      RECT 132.38 222.122 132.58 222.242 ;
      RECT 134.18 243 134.38 243.12 ;
      RECT 133.46 243 133.66 243.12 ;
      RECT 132.02 243 132.22 243.12 ;
      RECT 134.9 245.52 135.1 245.64 ;
      RECT 134.9 243.24 135.1 243.36 ;
      RECT 132.02 245.52 132.22 245.64 ;
      RECT 133.46 245.52 133.66 245.64 ;
      RECT 132.74 243.24 132.94 243.36 ;
      RECT 131.3 243.24 131.5 243.36 ;
      RECT 134.9 248.04 135.1 248.16 ;
      RECT 134.18 248.28 134.38 248.4 ;
      RECT 132.74 248.28 132.94 248.4 ;
      RECT 131.3 248.28 131.5 248.4 ;
      RECT 133.46 248.04 133.66 248.16 ;
      RECT 132.02 248.04 132.22 248.16 ;
      RECT 131.3 245.76 131.5 245.88 ;
      RECT 132.74 245.76 132.94 245.88 ;
      RECT 134.18 245.76 134.38 245.88 ;
      RECT 134.9 258.75 135.1 258.87 ;
      RECT 132.74 258.99 132.94 259.11 ;
      RECT 134.18 258.75 134.38 258.87 ;
      RECT 133.46 258.75 133.66 258.87 ;
      RECT 132.02 258.75 132.22 258.87 ;
      RECT 131.3 258.75 131.5 258.87 ;
      RECT 134.9 261.27 135.1 261.39 ;
      RECT 134.9 260.25 135.1 260.37 ;
      RECT 134.18 261.51 134.38 261.63 ;
      RECT 132.74 261.51 132.94 261.63 ;
      RECT 133.46 261.27 133.66 261.39 ;
      RECT 132.02 261.27 132.22 261.39 ;
      RECT 131.3 261.27 131.5 261.39 ;
      RECT 134.18 260.25 134.38 260.37 ;
      RECT 131.3 260.25 131.5 260.37 ;
      RECT 133.46 260.01 133.66 260.13 ;
      RECT 132.74 260.01 132.94 260.13 ;
      RECT 132.02 260.01 132.22 260.13 ;
      RECT 134.9 264.03 135.1 264.15 ;
      RECT 135.26 263.4 135.46 263.52 ;
      RECT 134.54 263.16 134.74 263.28 ;
      RECT 134.9 262.53 135.1 262.65 ;
      RECT 132.74 264.03 132.94 264.15 ;
      RECT 131.3 264.03 131.5 264.15 ;
      RECT 134.18 263.79 134.38 263.91 ;
      RECT 133.46 263.79 133.66 263.91 ;
      RECT 132.02 263.79 132.22 263.91 ;
      RECT 133.82 263.4 134.02 263.52 ;
      RECT 133.1 263.4 133.3 263.52 ;
      RECT 131.66 263.4 131.86 263.52 ;
      RECT 132.38 263.16 132.58 263.28 ;
      RECT 131.3 262.77 131.5 262.89 ;
      RECT 132.74 262.77 132.94 262.89 ;
      RECT 134.18 262.53 134.38 262.65 ;
      RECT 133.46 262.53 133.66 262.65 ;
      RECT 132.02 262.53 132.22 262.65 ;
      RECT 134.9 266.2885 135.1 266.4085 ;
      RECT 135.26 265.92 135.46 266.04 ;
      RECT 134.54 265.68 134.74 265.8 ;
      RECT 134.18 266.2885 134.38 266.4085 ;
      RECT 133.46 266.2885 133.66 266.4085 ;
      RECT 132.74 266.2885 132.94 266.4085 ;
      RECT 132.02 266.2885 132.22 266.4085 ;
      RECT 131.3 266.2885 131.5 266.4085 ;
      RECT 133.82 265.92 134.02 266.04 ;
      RECT 133.1 265.92 133.3 266.04 ;
      RECT 132.38 265.68 132.58 265.8 ;
      RECT 131.66 265.68 131.86 265.8 ;
      RECT 134.9 270.09 135.1 270.21 ;
      RECT 135.26 268.44 135.46 268.56 ;
      RECT 134.54 268.2 134.74 268.32 ;
      RECT 134.9 267.81 135.1 267.93 ;
      RECT 132.74 270.09 132.94 270.21 ;
      RECT 132.02 270.09 132.22 270.21 ;
      RECT 133.82 268.44 134.02 268.56 ;
      RECT 132.38 268.44 132.58 268.56 ;
      RECT 133.1 268.2 133.3 268.32 ;
      RECT 131.66 268.2 131.86 268.32 ;
      RECT 134.18 267.81 134.38 267.93 ;
      RECT 133.46 267.81 133.66 267.93 ;
      RECT 132.74 267.81 132.94 267.93 ;
      RECT 132.02 267.81 132.22 267.93 ;
      RECT 131.3 267.81 131.5 267.93 ;
      RECT 134.9 271.35 135.1 271.47 ;
      RECT 134.54 270.96 134.74 271.08 ;
      RECT 135.26 270.72 135.46 270.84 ;
      RECT 131.3 271.59 131.5 271.71 ;
      RECT 134.18 271.59 134.38 271.71 ;
      RECT 132.74 271.59 132.94 271.71 ;
      RECT 133.46 271.35 133.66 271.47 ;
      RECT 131.3 169.92 131.5 170.04 ;
      RECT 134.9 169.92 135.1 170.04 ;
      RECT 134.54 171.18 134.74 171.3 ;
      RECT 135.26 171.42 135.46 171.54 ;
      RECT 133.1 173.94 133.3 174.06 ;
      RECT 131.66 173.94 131.86 174.06 ;
      RECT 133.82 173.7 134.02 173.82 ;
      RECT 132.38 173.7 132.58 173.82 ;
      RECT 134.18 172.68 134.38 172.8 ;
      RECT 132.02 172.68 132.22 172.8 ;
      RECT 131.3 172.68 131.5 172.8 ;
      RECT 132.74 172.44 132.94 172.56 ;
      RECT 133.46 172.44 133.66 172.56 ;
      RECT 135.26 173.94 135.46 174.06 ;
      RECT 134.54 173.94 134.74 174.06 ;
      RECT 134.9 172.44 135.1 172.56 ;
      RECT 133.46 177.48 133.66 177.6 ;
      RECT 132.74 177.48 132.94 177.6 ;
      RECT 131.3 177.48 131.5 177.6 ;
      RECT 133.1 176.46 133.3 176.58 ;
      RECT 131.66 176.46 131.86 176.58 ;
      RECT 133.82 176.22 134.02 176.34 ;
      RECT 132.38 176.22 132.58 176.34 ;
      RECT 134.18 175.2 134.38 175.32 ;
      RECT 132.74 175.2 132.94 175.32 ;
      RECT 132.02 175.2 132.22 175.32 ;
      RECT 131.3 174.96 131.5 175.08 ;
      RECT 133.46 174.96 133.66 175.08 ;
      RECT 134.9 177.48 135.1 177.6 ;
      RECT 135.26 176.46 135.46 176.58 ;
      RECT 134.54 176.22 134.74 176.34 ;
      RECT 134.9 174.96 135.1 175.08 ;
      RECT 133.46 180 133.66 180.12 ;
      RECT 132.02 180 132.22 180.12 ;
      RECT 131.66 178.98 131.86 179.1 ;
      RECT 133.1 178.98 133.3 179.1 ;
      RECT 132.38 178.74 132.58 178.86 ;
      RECT 133.82 178.74 134.02 178.86 ;
      RECT 134.18 177.72 134.38 177.84 ;
      RECT 132.02 177.72 132.22 177.84 ;
      RECT 134.54 178.98 134.74 179.1 ;
      RECT 135.26 178.74 135.46 178.86 ;
      RECT 132.74 180.24 132.94 180.36 ;
      RECT 131.3 180.24 131.5 180.36 ;
      RECT 131.3 192.84 131.5 192.96 ;
      RECT 132.02 192.84 132.22 192.96 ;
      RECT 132.74 192.84 132.94 192.96 ;
      RECT 133.46 192.6 133.66 192.72 ;
      RECT 134.18 192.6 134.38 192.72 ;
      RECT 134.9 192.6 135.1 192.72 ;
      RECT 132.74 195.36 132.94 195.48 ;
      RECT 131.3 195.12 131.5 195.24 ;
      RECT 132.02 195.12 132.22 195.24 ;
      RECT 133.46 195.12 133.66 195.24 ;
      RECT 134.18 195.12 134.38 195.24 ;
      RECT 134.9 195.12 135.1 195.24 ;
      RECT 131.3 197.88 131.5 198 ;
      RECT 134.18 197.88 134.38 198 ;
      RECT 133.46 197.64 133.66 197.76 ;
      RECT 132.74 197.64 132.94 197.76 ;
      RECT 132.02 197.64 132.22 197.76 ;
      RECT 134.9 197.64 135.1 197.76 ;
      RECT 134.18 200.4 134.38 200.52 ;
      RECT 133.46 200.16 133.66 200.28 ;
      RECT 132.74 200.16 132.94 200.28 ;
      RECT 132.02 200.16 132.22 200.28 ;
      RECT 131.3 200.16 131.5 200.28 ;
      RECT 134.9 200.16 135.1 200.28 ;
      RECT 134.18 202.92 134.38 203.04 ;
      RECT 131.3 202.92 131.5 203.04 ;
      RECT 132.02 202.68 132.22 202.8 ;
      RECT 132.74 202.68 132.94 202.8 ;
      RECT 133.46 202.68 133.66 202.8 ;
      RECT 134.9 202.68 135.1 202.8 ;
      RECT 132.74 205.44 132.94 205.56 ;
      RECT 134.18 205.44 134.38 205.56 ;
      RECT 131.3 205.2 131.5 205.32 ;
      RECT 132.02 205.2 132.22 205.32 ;
      RECT 133.46 205.2 133.66 205.32 ;
      RECT 134.9 205.2 135.1 205.32 ;
      RECT 132.02 210.24 132.22 210.36 ;
      RECT 133.46 210.24 133.66 210.36 ;
      RECT 131.3 207.96 131.5 208.08 ;
      RECT 134.18 207.96 134.38 208.08 ;
      RECT 132.02 207.72 132.22 207.84 ;
      RECT 132.74 207.72 132.94 207.84 ;
      RECT 133.46 207.72 133.66 207.84 ;
      RECT 134.9 210.24 135.1 210.36 ;
      RECT 134.9 207.72 135.1 207.84 ;
      RECT 131.3 212.76 131.5 212.88 ;
      RECT 132.74 212.76 132.94 212.88 ;
      RECT 133.46 212.76 133.66 212.88 ;
      RECT 131.3 210.48 131.5 210.6 ;
      RECT 132.74 210.48 132.94 210.6 ;
      RECT 134.18 210.48 134.38 210.6 ;
      RECT 134.9 212.76 135.1 212.88 ;
      RECT 132.74 215.52 132.94 215.64 ;
      RECT 134.18 215.52 134.38 215.64 ;
      RECT 131.3 215.28 131.5 215.4 ;
      RECT 132.02 215.28 132.22 215.4 ;
      RECT 133.46 215.28 133.66 215.4 ;
      RECT 134.18 213 134.38 213.12 ;
      RECT 133.46 139.92 133.66 140.04 ;
      RECT 132.02 139.92 132.22 140.04 ;
      RECT 132.74 139.68 132.94 139.8 ;
      RECT 131.3 139.68 131.5 139.8 ;
      RECT 134.54 143.7 134.74 143.82 ;
      RECT 135.26 143.7 135.46 143.82 ;
      RECT 134.9 142.2 135.1 142.32 ;
      RECT 133.82 143.46 134.02 143.58 ;
      RECT 132.38 143.46 132.58 143.58 ;
      RECT 131.66 143.46 131.86 143.58 ;
      RECT 134.18 142.44 134.38 142.56 ;
      RECT 132.02 142.44 132.22 142.56 ;
      RECT 133.46 142.2 133.66 142.32 ;
      RECT 132.74 142.2 132.94 142.32 ;
      RECT 131.3 142.2 131.5 142.32 ;
      RECT 133.1 143.7 133.3 143.82 ;
      RECT 134.9 147.24 135.1 147.36 ;
      RECT 134.54 146.22 134.74 146.34 ;
      RECT 135.26 145.98 135.46 146.1 ;
      RECT 134.9 144.72 135.1 144.84 ;
      RECT 132.74 147.24 132.94 147.36 ;
      RECT 131.3 147.24 131.5 147.36 ;
      RECT 132.38 146.22 132.58 146.34 ;
      RECT 133.82 145.98 134.02 146.1 ;
      RECT 133.1 145.98 133.3 146.1 ;
      RECT 131.66 145.98 131.86 146.1 ;
      RECT 134.18 144.96 134.38 145.08 ;
      RECT 132.02 144.96 132.22 145.08 ;
      RECT 131.3 144.96 131.5 145.08 ;
      RECT 132.74 144.72 132.94 144.84 ;
      RECT 133.46 144.72 133.66 144.84 ;
      RECT 134.9 149.76 135.1 149.88 ;
      RECT 134.54 148.74 134.74 148.86 ;
      RECT 135.26 148.5 135.46 148.62 ;
      RECT 134.18 150 134.38 150.12 ;
      RECT 132.74 150 132.94 150.12 ;
      RECT 131.3 150 131.5 150.12 ;
      RECT 133.46 149.76 133.66 149.88 ;
      RECT 132.02 149.76 132.22 149.88 ;
      RECT 133.1 148.74 133.3 148.86 ;
      RECT 131.66 148.74 131.86 148.86 ;
      RECT 132.38 148.5 132.58 148.62 ;
      RECT 133.82 148.5 134.02 148.62 ;
      RECT 133.46 147.48 133.66 147.6 ;
      RECT 132.02 147.48 132.22 147.6 ;
      RECT 134.18 147.48 134.38 147.6 ;
      RECT 134.9 152.28 135.1 152.4 ;
      RECT 134.54 151.26 134.74 151.38 ;
      RECT 135.26 151.02 135.46 151.14 ;
      RECT 134.18 152.52 134.38 152.64 ;
      RECT 132.74 152.52 132.94 152.64 ;
      RECT 131.3 152.52 131.5 152.64 ;
      RECT 133.46 152.28 133.66 152.4 ;
      RECT 132.02 152.28 132.22 152.4 ;
      RECT 133.1 151.26 133.3 151.38 ;
      RECT 131.66 151.26 131.86 151.38 ;
      RECT 133.82 151.02 134.02 151.14 ;
      RECT 132.38 151.02 132.58 151.14 ;
      RECT 134.9 154.8 135.1 154.92 ;
      RECT 134.54 153.78 134.74 153.9 ;
      RECT 135.26 153.54 135.46 153.66 ;
      RECT 132.74 155.04 132.94 155.16 ;
      RECT 134.18 154.8 134.38 154.92 ;
      RECT 133.46 154.8 133.66 154.92 ;
      RECT 132.02 154.8 132.22 154.92 ;
      RECT 131.3 154.8 131.5 154.92 ;
      RECT 133.1 153.78 133.3 153.9 ;
      RECT 131.66 153.78 131.86 153.9 ;
      RECT 132.38 153.54 132.58 153.66 ;
      RECT 133.82 153.54 134.02 153.66 ;
      RECT 134.54 156.3 134.74 156.42 ;
      RECT 135.26 156.06 135.46 156.18 ;
      RECT 133.1 156.3 133.3 156.42 ;
      RECT 131.66 156.3 131.86 156.42 ;
      RECT 133.82 156.06 134.02 156.18 ;
      RECT 132.38 156.06 132.58 156.18 ;
      RECT 134.54 166.14 134.74 166.26 ;
      RECT 135.26 166.14 135.46 166.26 ;
      RECT 133.82 166.38 134.02 166.5 ;
      RECT 131.66 166.14 131.86 166.26 ;
      RECT 132.38 166.14 132.58 166.26 ;
      RECT 133.1 166.14 133.3 166.26 ;
      RECT 134.54 168.66 134.74 168.78 ;
      RECT 135.26 168.66 135.46 168.78 ;
      RECT 134.9 167.4 135.1 167.52 ;
      RECT 133.82 168.9 134.02 169.02 ;
      RECT 133.1 168.9 133.3 169.02 ;
      RECT 131.66 168.66 131.86 168.78 ;
      RECT 132.38 168.66 132.58 168.78 ;
      RECT 134.18 167.64 134.38 167.76 ;
      RECT 133.46 167.64 133.66 167.76 ;
      RECT 132.74 167.4 132.94 167.52 ;
      RECT 132.02 167.4 132.22 167.52 ;
      RECT 131.3 167.4 131.5 167.52 ;
      RECT 133.1 171.42 133.3 171.54 ;
      RECT 133.82 171.18 134.02 171.3 ;
      RECT 132.38 171.18 132.58 171.3 ;
      RECT 131.66 171.18 131.86 171.3 ;
      RECT 134.18 170.16 134.38 170.28 ;
      RECT 132.74 170.16 132.94 170.28 ;
      RECT 133.46 169.92 133.66 170.04 ;
      RECT 132.02 169.92 132.22 170.04 ;
      RECT 134.18 119.52 134.38 119.64 ;
      RECT 132.74 119.52 132.94 119.64 ;
      RECT 133.82 118.324 134.02 118.444 ;
      RECT 133.1 118.324 133.3 118.444 ;
      RECT 134.9 122.28 135.1 122.4 ;
      RECT 134.54 121.02 134.74 121.14 ;
      RECT 135.26 120.78 135.46 120.9 ;
      RECT 131.3 122.28 131.5 122.4 ;
      RECT 132.74 122.28 132.94 122.4 ;
      RECT 133.46 122.28 133.66 122.4 ;
      RECT 132.02 122.04 132.22 122.16 ;
      RECT 134.18 122.04 134.38 122.16 ;
      RECT 133.82 121.02 134.02 121.14 ;
      RECT 131.66 120.78 131.86 120.9 ;
      RECT 132.38 120.78 132.58 120.9 ;
      RECT 133.1 120.78 133.3 120.9 ;
      RECT 134.9 124.56 135.1 124.68 ;
      RECT 135.26 123.54 135.46 123.66 ;
      RECT 134.54 123.3 134.74 123.42 ;
      RECT 132.02 124.8 132.22 124.92 ;
      RECT 132.74 124.8 132.94 124.92 ;
      RECT 131.3 124.56 131.5 124.68 ;
      RECT 133.46 124.56 133.66 124.68 ;
      RECT 134.18 124.56 134.38 124.68 ;
      RECT 133.1 123.54 133.3 123.66 ;
      RECT 131.66 123.3 131.86 123.42 ;
      RECT 132.38 123.3 132.58 123.42 ;
      RECT 133.82 123.3 134.02 123.42 ;
      RECT 134.9 127.08 135.1 127.2 ;
      RECT 134.54 125.82 134.74 125.94 ;
      RECT 135.26 125.82 135.46 125.94 ;
      RECT 133.46 127.32 133.66 127.44 ;
      RECT 132.02 127.32 132.22 127.44 ;
      RECT 131.3 127.32 131.5 127.44 ;
      RECT 134.18 127.08 134.38 127.2 ;
      RECT 132.74 127.08 132.94 127.2 ;
      RECT 133.82 126.06 134.02 126.18 ;
      RECT 131.66 125.82 131.86 125.94 ;
      RECT 132.38 125.82 132.58 125.94 ;
      RECT 133.1 125.82 133.3 125.94 ;
      RECT 135.26 130.86 135.46 130.98 ;
      RECT 134.9 129.6 135.1 129.72 ;
      RECT 134.54 128.58 134.74 128.7 ;
      RECT 135.26 128.34 135.46 128.46 ;
      RECT 133.82 130.86 134.02 130.98 ;
      RECT 132.38 130.86 132.58 130.98 ;
      RECT 132.02 129.84 132.22 129.96 ;
      RECT 133.46 129.84 133.66 129.96 ;
      RECT 134.18 129.6 134.38 129.72 ;
      RECT 132.74 129.6 132.94 129.72 ;
      RECT 131.3 129.6 131.5 129.72 ;
      RECT 133.1 128.58 133.3 128.7 ;
      RECT 131.66 128.58 131.86 128.7 ;
      RECT 133.82 128.34 134.02 128.46 ;
      RECT 132.38 128.34 132.58 128.46 ;
      RECT 134.54 133.62 134.74 133.74 ;
      RECT 135.26 133.38 135.46 133.5 ;
      RECT 134.9 132.12 135.1 132.24 ;
      RECT 134.54 131.1 134.74 131.22 ;
      RECT 133.1 133.62 133.3 133.74 ;
      RECT 131.66 133.38 131.86 133.5 ;
      RECT 132.38 133.38 132.58 133.5 ;
      RECT 133.82 133.38 134.02 133.5 ;
      RECT 134.18 132.36 134.38 132.48 ;
      RECT 132.74 132.36 132.94 132.48 ;
      RECT 131.3 132.36 131.5 132.48 ;
      RECT 133.46 132.12 133.66 132.24 ;
      RECT 132.02 132.12 132.22 132.24 ;
      RECT 131.66 131.1 131.86 131.22 ;
      RECT 133.1 131.1 133.3 131.22 ;
      RECT 134.54 136.14 134.74 136.26 ;
      RECT 135.26 135.9 135.46 136.02 ;
      RECT 134.9 134.64 135.1 134.76 ;
      RECT 133.82 136.14 134.02 136.26 ;
      RECT 133.1 135.9 133.3 136.02 ;
      RECT 131.66 135.9 131.86 136.02 ;
      RECT 132.38 135.9 132.58 136.02 ;
      RECT 134.18 134.88 134.38 135 ;
      RECT 132.74 134.88 132.94 135 ;
      RECT 131.3 134.88 131.5 135 ;
      RECT 133.46 134.64 133.66 134.76 ;
      RECT 132.02 134.64 132.22 134.76 ;
      RECT 135.26 138.66 135.46 138.78 ;
      RECT 134.54 138.66 134.74 138.78 ;
      RECT 134.9 137.4 135.1 137.52 ;
      RECT 131.66 138.66 131.86 138.78 ;
      RECT 132.38 138.42 132.58 138.54 ;
      RECT 133.1 138.42 133.3 138.54 ;
      RECT 133.82 138.42 134.02 138.54 ;
      RECT 132.02 137.4 132.22 137.52 ;
      RECT 131.3 137.4 131.5 137.52 ;
      RECT 132.74 137.16 132.94 137.28 ;
      RECT 133.46 137.16 133.66 137.28 ;
      RECT 134.18 137.16 134.38 137.28 ;
      RECT 135.26 140.94 135.46 141.06 ;
      RECT 134.54 140.94 134.74 141.06 ;
      RECT 134.9 139.68 135.1 139.8 ;
      RECT 133.1 141.18 133.3 141.3 ;
      RECT 132.38 141.18 132.58 141.3 ;
      RECT 131.66 140.94 131.86 141.06 ;
      RECT 133.82 140.94 134.02 141.06 ;
      RECT 134.18 139.92 134.38 140.04 ;
      RECT 129.14 261.27 129.34 261.39 ;
      RECT 130.58 261.27 130.78 261.39 ;
      RECT 126.98 261.51 127.18 261.63 ;
      RECT 129.86 261.51 130.06 261.63 ;
      RECT 126.98 262.53 127.18 262.65 ;
      RECT 127.7 262.53 127.9 262.65 ;
      RECT 129.14 262.53 129.34 262.65 ;
      RECT 129.86 262.53 130.06 262.65 ;
      RECT 128.42 262.77 128.62 262.89 ;
      RECT 130.58 262.77 130.78 262.89 ;
      RECT 127.34 263.16 127.54 263.28 ;
      RECT 128.78 263.16 128.98 263.28 ;
      RECT 129.5 263.16 129.7 263.28 ;
      RECT 130.94 263.16 131.14 263.28 ;
      RECT 130.22 263.4 130.42 263.52 ;
      RECT 128.06 263.4 128.26 263.52 ;
      RECT 129.14 263.79 129.34 263.91 ;
      RECT 130.58 263.79 130.78 263.91 ;
      RECT 126.98 263.79 127.18 263.91 ;
      RECT 128.42 264.03 128.62 264.15 ;
      RECT 129.86 264.03 130.06 264.15 ;
      RECT 127.7 264.03 127.9 264.15 ;
      RECT 128.06 265.68 128.26 265.8 ;
      RECT 129.5 265.68 129.7 265.8 ;
      RECT 130.22 265.68 130.42 265.8 ;
      RECT 127.34 265.92 127.54 266.04 ;
      RECT 128.78 265.92 128.98 266.04 ;
      RECT 130.94 265.92 131.14 266.04 ;
      RECT 126.98 266.2885 127.18 266.4085 ;
      RECT 127.7 266.2885 127.9 266.4085 ;
      RECT 128.42 266.2885 128.62 266.4085 ;
      RECT 129.14 266.2885 129.34 266.4085 ;
      RECT 129.86 266.2885 130.06 266.4085 ;
      RECT 130.58 266.2885 130.78 266.4085 ;
      RECT 126.98 267.81 127.18 267.93 ;
      RECT 127.7 267.81 127.9 267.93 ;
      RECT 128.42 267.81 128.62 267.93 ;
      RECT 129.14 267.81 129.34 267.93 ;
      RECT 129.86 267.81 130.06 267.93 ;
      RECT 130.58 267.81 130.78 267.93 ;
      RECT 128.06 268.2 128.26 268.32 ;
      RECT 129.5 268.2 129.7 268.32 ;
      RECT 130.94 268.2 131.14 268.32 ;
      RECT 127.34 268.44 127.54 268.56 ;
      RECT 128.78 268.44 128.98 268.56 ;
      RECT 130.22 268.44 130.42 268.56 ;
      RECT 127.7 270.09 127.9 270.21 ;
      RECT 129.14 270.09 129.34 270.21 ;
      RECT 130.58 270.09 130.78 270.21 ;
      RECT 126.98 270.33 127.18 270.45 ;
      RECT 128.42 270.33 128.62 270.45 ;
      RECT 129.86 270.33 130.06 270.45 ;
      RECT 127.34 270.72 127.54 270.84 ;
      RECT 128.78 270.72 128.98 270.84 ;
      RECT 130.94 270.72 131.14 270.84 ;
      RECT 129.5 270.96 129.7 271.08 ;
      RECT 128.06 270.96 128.26 271.08 ;
      RECT 130.22 270.96 130.42 271.08 ;
      RECT 126.98 271.35 127.18 271.47 ;
      RECT 128.42 271.35 128.62 271.47 ;
      RECT 130.58 271.35 130.78 271.47 ;
      RECT 127.7 271.59 127.9 271.71 ;
      RECT 129.14 271.59 129.34 271.71 ;
      RECT 129.86 271.59 130.06 271.71 ;
      RECT 130.22 273.48 130.42 273.6 ;
      RECT 129.5 273.48 129.7 273.6 ;
      RECT 128.78 273.48 128.98 273.6 ;
      RECT 127.34 273.48 127.54 273.6 ;
      RECT 130.94 273.24 131.14 273.36 ;
      RECT 128.06 273.24 128.26 273.36 ;
      RECT 130.22 276 130.42 276.12 ;
      RECT 128.78 276 128.98 276.12 ;
      RECT 127.34 276 127.54 276.12 ;
      RECT 130.94 275.76 131.14 275.88 ;
      RECT 129.5 275.76 129.7 275.88 ;
      RECT 128.06 275.76 128.26 275.88 ;
      RECT 130.94 278.28 131.14 278.4 ;
      RECT 129.5 278.28 129.7 278.4 ;
      RECT 128.06 278.28 128.26 278.4 ;
      RECT 130.22 278.52 130.42 278.64 ;
      RECT 128.78 278.52 128.98 278.64 ;
      RECT 127.34 278.52 127.54 278.64 ;
      RECT 129.86 305.625 130.06 305.745 ;
      RECT 130.58 305.625 130.78 305.745 ;
      RECT 130.58 323.3835 130.78 323.5035 ;
      RECT 129.86 323.3835 130.06 323.5035 ;
      RECT 129.14 323.3835 129.34 323.5035 ;
      RECT 128.42 323.3835 128.62 323.5035 ;
      RECT 127.7 323.3835 127.9 323.5035 ;
      RECT 126.98 323.3835 127.18 323.5035 ;
      RECT 128.42 348.339 128.62 348.459 ;
      RECT 127.7 348.339 127.9 348.459 ;
      RECT 126.98 348.339 127.18 348.459 ;
      RECT 129.14 348.339 129.34 348.459 ;
      RECT 129.86 348.339 130.06 348.459 ;
      RECT 130.58 348.339 130.78 348.459 ;
      RECT 134.9 119.52 135.1 119.64 ;
      RECT 134.54 118.324 134.74 118.444 ;
      RECT 135.26 118.084 135.46 118.204 ;
      RECT 132.02 119.76 132.22 119.88 ;
      RECT 133.46 119.76 133.66 119.88 ;
      RECT 131.3 119.76 131.5 119.88 ;
      RECT 127.7 192.6 127.9 192.72 ;
      RECT 129.14 192.6 129.34 192.72 ;
      RECT 129.86 192.6 130.06 192.72 ;
      RECT 130.58 192.6 130.78 192.72 ;
      RECT 127.7 195.12 127.9 195.24 ;
      RECT 129.14 195.12 129.34 195.24 ;
      RECT 130.58 195.36 130.78 195.48 ;
      RECT 129.86 195.36 130.06 195.48 ;
      RECT 128.42 195.36 128.62 195.48 ;
      RECT 126.98 195.36 127.18 195.48 ;
      RECT 127.7 197.88 127.9 198 ;
      RECT 128.42 197.88 128.62 198 ;
      RECT 129.86 197.88 130.06 198 ;
      RECT 130.58 197.64 130.78 197.76 ;
      RECT 129.14 197.64 129.34 197.76 ;
      RECT 126.98 197.64 127.18 197.76 ;
      RECT 129.86 200.4 130.06 200.52 ;
      RECT 129.14 200.4 129.34 200.52 ;
      RECT 130.58 200.16 130.78 200.28 ;
      RECT 128.42 200.16 128.62 200.28 ;
      RECT 127.7 200.16 127.9 200.28 ;
      RECT 126.98 200.16 127.18 200.28 ;
      RECT 129.86 202.92 130.06 203.04 ;
      RECT 128.42 202.92 128.62 203.04 ;
      RECT 126.98 202.68 127.18 202.8 ;
      RECT 127.7 202.68 127.9 202.8 ;
      RECT 129.14 202.68 129.34 202.8 ;
      RECT 130.58 202.68 130.78 202.8 ;
      RECT 126.98 205.44 127.18 205.56 ;
      RECT 129.14 205.44 129.34 205.56 ;
      RECT 129.86 205.44 130.06 205.56 ;
      RECT 127.7 205.2 127.9 205.32 ;
      RECT 128.42 205.2 128.62 205.32 ;
      RECT 130.58 205.2 130.78 205.32 ;
      RECT 127.7 207.96 127.9 208.08 ;
      RECT 128.42 207.96 128.62 208.08 ;
      RECT 129.86 207.96 130.06 208.08 ;
      RECT 126.98 207.72 127.18 207.84 ;
      RECT 129.14 207.72 129.34 207.84 ;
      RECT 130.58 207.72 130.78 207.84 ;
      RECT 126.98 210.48 127.18 210.6 ;
      RECT 128.42 210.48 128.62 210.6 ;
      RECT 129.86 210.48 130.06 210.6 ;
      RECT 127.7 210.24 127.9 210.36 ;
      RECT 129.14 210.24 129.34 210.36 ;
      RECT 130.58 210.24 130.78 210.36 ;
      RECT 126.98 212.76 127.18 212.88 ;
      RECT 127.7 212.76 127.9 212.88 ;
      RECT 128.42 212.76 128.62 212.88 ;
      RECT 130.58 213 130.78 213.12 ;
      RECT 129.86 213 130.06 213.12 ;
      RECT 129.14 213 129.34 213.12 ;
      RECT 129.14 215.52 129.34 215.64 ;
      RECT 130.58 215.52 130.78 215.64 ;
      RECT 126.98 215.28 127.18 215.4 ;
      RECT 127.7 215.28 127.9 215.4 ;
      RECT 128.42 215.28 128.62 215.4 ;
      RECT 129.86 215.28 130.06 215.4 ;
      RECT 128.06 222.362 128.26 222.482 ;
      RECT 128.78 222.362 128.98 222.482 ;
      RECT 130.22 222.362 130.42 222.482 ;
      RECT 130.94 222.362 131.14 222.482 ;
      RECT 127.34 222.122 127.54 222.242 ;
      RECT 129.5 222.122 129.7 222.242 ;
      RECT 126.98 223.08 127.18 223.2 ;
      RECT 128.42 223.08 128.62 223.2 ;
      RECT 129.86 223.08 130.06 223.2 ;
      RECT 130.58 223.08 130.78 223.2 ;
      RECT 127.7 222.84 127.9 222.96 ;
      RECT 129.14 222.84 129.34 222.96 ;
      RECT 129.86 243.24 130.06 243.36 ;
      RECT 128.42 243.24 128.62 243.36 ;
      RECT 126.98 243.24 127.18 243.36 ;
      RECT 130.58 243 130.78 243.12 ;
      RECT 129.14 243 129.34 243.12 ;
      RECT 127.7 243 127.9 243.12 ;
      RECT 127.7 245.52 127.9 245.64 ;
      RECT 129.86 245.52 130.06 245.64 ;
      RECT 130.58 245.52 130.78 245.64 ;
      RECT 126.98 245.76 127.18 245.88 ;
      RECT 128.42 245.76 128.62 245.88 ;
      RECT 129.14 245.76 129.34 245.88 ;
      RECT 126.98 248.04 127.18 248.16 ;
      RECT 128.42 248.04 128.62 248.16 ;
      RECT 129.86 248.04 130.06 248.16 ;
      RECT 127.7 248.28 127.9 248.4 ;
      RECT 129.14 248.28 129.34 248.4 ;
      RECT 130.58 248.28 130.78 248.4 ;
      RECT 127.7 258.75 127.9 258.87 ;
      RECT 129.14 258.75 129.34 258.87 ;
      RECT 129.86 258.75 130.06 258.87 ;
      RECT 126.98 258.99 127.18 259.11 ;
      RECT 128.42 258.99 128.62 259.11 ;
      RECT 130.58 258.99 130.78 259.11 ;
      RECT 126.98 260.01 127.18 260.13 ;
      RECT 127.7 260.01 127.9 260.13 ;
      RECT 129.14 260.01 129.34 260.13 ;
      RECT 130.58 260.01 130.78 260.13 ;
      RECT 128.42 260.25 128.62 260.37 ;
      RECT 129.86 260.25 130.06 260.37 ;
      RECT 127.7 261.27 127.9 261.39 ;
      RECT 128.42 261.27 128.62 261.39 ;
      RECT 128.42 152.28 128.62 152.4 ;
      RECT 129.86 152.28 130.06 152.4 ;
      RECT 130.58 152.28 130.78 152.4 ;
      RECT 127.7 152.52 127.9 152.64 ;
      RECT 129.14 152.52 129.34 152.64 ;
      RECT 130.94 153.54 131.14 153.66 ;
      RECT 129.5 153.54 129.7 153.66 ;
      RECT 128.06 153.54 128.26 153.66 ;
      RECT 127.34 153.78 127.54 153.9 ;
      RECT 128.78 153.78 128.98 153.9 ;
      RECT 130.22 153.78 130.42 153.9 ;
      RECT 128.42 154.8 128.62 154.92 ;
      RECT 130.58 154.8 130.78 154.92 ;
      RECT 126.98 155.04 127.18 155.16 ;
      RECT 127.7 155.04 127.9 155.16 ;
      RECT 129.86 155.04 130.06 155.16 ;
      RECT 129.14 155.04 129.34 155.16 ;
      RECT 128.06 156.06 128.26 156.18 ;
      RECT 129.5 156.06 129.7 156.18 ;
      RECT 130.94 156.06 131.14 156.18 ;
      RECT 127.34 156.3 127.54 156.42 ;
      RECT 128.78 156.3 128.98 156.42 ;
      RECT 130.22 156.3 130.42 156.42 ;
      RECT 126.98 164.88 127.18 165 ;
      RECT 130.94 166.14 131.14 166.26 ;
      RECT 130.22 166.14 130.42 166.26 ;
      RECT 129.5 166.14 129.7 166.26 ;
      RECT 128.06 166.14 128.26 166.26 ;
      RECT 128.78 166.38 128.98 166.5 ;
      RECT 127.34 166.38 127.54 166.5 ;
      RECT 126.98 167.4 127.18 167.52 ;
      RECT 127.7 167.4 127.9 167.52 ;
      RECT 129.14 167.4 129.34 167.52 ;
      RECT 129.86 167.4 130.06 167.52 ;
      RECT 130.58 167.4 130.78 167.52 ;
      RECT 128.42 167.64 128.62 167.76 ;
      RECT 130.22 168.66 130.42 168.78 ;
      RECT 129.5 168.66 129.7 168.78 ;
      RECT 127.34 168.9 127.54 169.02 ;
      RECT 128.06 168.9 128.26 169.02 ;
      RECT 128.78 168.9 128.98 169.02 ;
      RECT 130.94 168.9 131.14 169.02 ;
      RECT 127.7 169.92 127.9 170.04 ;
      RECT 129.14 169.92 129.34 170.04 ;
      RECT 130.58 169.92 130.78 170.04 ;
      RECT 126.98 170.16 127.18 170.28 ;
      RECT 128.42 170.16 128.62 170.28 ;
      RECT 129.86 170.16 130.06 170.28 ;
      RECT 128.06 171.18 128.26 171.3 ;
      RECT 128.78 171.18 128.98 171.3 ;
      RECT 130.94 171.18 131.14 171.3 ;
      RECT 130.22 171.42 130.42 171.54 ;
      RECT 129.5 171.42 129.7 171.54 ;
      RECT 127.34 171.42 127.54 171.54 ;
      RECT 130.58 172.44 130.78 172.56 ;
      RECT 129.86 172.44 130.06 172.56 ;
      RECT 129.14 172.44 129.34 172.56 ;
      RECT 127.7 172.44 127.9 172.56 ;
      RECT 126.98 172.44 127.18 172.56 ;
      RECT 128.42 172.68 128.62 172.8 ;
      RECT 129.5 173.7 129.7 173.82 ;
      RECT 130.22 173.7 130.42 173.82 ;
      RECT 130.94 173.7 131.14 173.82 ;
      RECT 127.34 173.94 127.54 174.06 ;
      RECT 128.06 173.94 128.26 174.06 ;
      RECT 128.78 173.94 128.98 174.06 ;
      RECT 130.58 174.96 130.78 175.08 ;
      RECT 129.14 174.96 129.34 175.08 ;
      RECT 127.7 174.96 127.9 175.08 ;
      RECT 126.98 174.96 127.18 175.08 ;
      RECT 128.42 175.2 128.62 175.32 ;
      RECT 129.86 175.2 130.06 175.32 ;
      RECT 129.5 176.22 129.7 176.34 ;
      RECT 130.94 176.22 131.14 176.34 ;
      RECT 128.06 176.22 128.26 176.34 ;
      RECT 128.78 176.22 128.98 176.34 ;
      RECT 127.34 176.46 127.54 176.58 ;
      RECT 130.22 176.46 130.42 176.58 ;
      RECT 127.7 177.72 127.9 177.84 ;
      RECT 128.42 177.72 128.62 177.84 ;
      RECT 129.86 177.72 130.06 177.84 ;
      RECT 130.94 178.74 131.14 178.86 ;
      RECT 129.5 178.74 129.7 178.86 ;
      RECT 128.06 178.74 128.26 178.86 ;
      RECT 126.98 177.48 127.18 177.6 ;
      RECT 129.14 177.48 129.34 177.6 ;
      RECT 130.58 177.48 130.78 177.6 ;
      RECT 130.22 178.98 130.42 179.1 ;
      RECT 128.78 178.98 128.98 179.1 ;
      RECT 127.34 178.98 127.54 179.1 ;
      RECT 126.98 180 127.18 180.12 ;
      RECT 127.7 180 127.9 180.12 ;
      RECT 129.14 180 129.34 180.12 ;
      RECT 130.58 180 130.78 180.12 ;
      RECT 129.86 180.24 130.06 180.36 ;
      RECT 128.42 180.24 128.62 180.36 ;
      RECT 126.98 182.52 127.18 182.64 ;
      RECT 126.98 185.04 127.18 185.16 ;
      RECT 126.98 187.56 127.18 187.68 ;
      RECT 126.98 190.08 127.18 190.2 ;
      RECT 128.42 192.84 128.62 192.96 ;
      RECT 126.98 192.84 127.18 192.96 ;
      RECT 129.5 130.86 129.7 130.98 ;
      RECT 130.94 131.1 131.14 131.22 ;
      RECT 130.22 131.1 130.42 131.22 ;
      RECT 128.06 131.1 128.26 131.22 ;
      RECT 127.34 131.1 127.54 131.22 ;
      RECT 127.7 132.12 127.9 132.24 ;
      RECT 129.14 132.12 129.34 132.24 ;
      RECT 130.58 132.12 130.78 132.24 ;
      RECT 126.98 132.36 127.18 132.48 ;
      RECT 128.42 132.36 128.62 132.48 ;
      RECT 129.86 132.36 130.06 132.48 ;
      RECT 130.94 133.38 131.14 133.5 ;
      RECT 130.22 133.38 130.42 133.5 ;
      RECT 127.34 133.62 127.54 133.74 ;
      RECT 128.06 133.62 128.26 133.74 ;
      RECT 128.78 133.62 128.98 133.74 ;
      RECT 129.5 133.62 129.7 133.74 ;
      RECT 126.98 134.64 127.18 134.76 ;
      RECT 128.42 134.64 128.62 134.76 ;
      RECT 129.14 134.64 129.34 134.76 ;
      RECT 130.58 134.64 130.78 134.76 ;
      RECT 127.7 134.88 127.9 135 ;
      RECT 129.86 134.88 130.06 135 ;
      RECT 127.34 135.9 127.54 136.02 ;
      RECT 128.78 135.9 128.98 136.02 ;
      RECT 130.94 135.9 131.14 136.02 ;
      RECT 130.22 136.14 130.42 136.26 ;
      RECT 129.5 136.14 129.7 136.26 ;
      RECT 128.06 136.14 128.26 136.26 ;
      RECT 130.58 137.16 130.78 137.28 ;
      RECT 128.42 137.16 128.62 137.28 ;
      RECT 127.7 137.16 127.9 137.28 ;
      RECT 126.98 137.4 127.18 137.52 ;
      RECT 129.14 137.4 129.34 137.52 ;
      RECT 129.86 137.4 130.06 137.52 ;
      RECT 128.06 138.42 128.26 138.54 ;
      RECT 130.94 138.42 131.14 138.54 ;
      RECT 129.5 138.42 129.7 138.54 ;
      RECT 127.34 138.66 127.54 138.78 ;
      RECT 128.78 138.66 128.98 138.78 ;
      RECT 130.22 138.66 130.42 138.78 ;
      RECT 126.98 139.68 127.18 139.8 ;
      RECT 127.7 139.68 127.9 139.8 ;
      RECT 129.86 139.68 130.06 139.8 ;
      RECT 128.42 139.92 128.62 140.04 ;
      RECT 129.14 139.92 129.34 140.04 ;
      RECT 130.58 139.92 130.78 140.04 ;
      RECT 130.94 140.94 131.14 141.06 ;
      RECT 129.5 140.94 129.7 141.06 ;
      RECT 128.06 140.94 128.26 141.06 ;
      RECT 127.34 141.18 127.54 141.3 ;
      RECT 128.78 141.18 128.98 141.3 ;
      RECT 130.22 141.18 130.42 141.3 ;
      RECT 127.7 142.2 127.9 142.32 ;
      RECT 129.86 142.2 130.06 142.32 ;
      RECT 126.98 142.44 127.18 142.56 ;
      RECT 128.42 142.44 128.62 142.56 ;
      RECT 129.14 142.44 129.34 142.56 ;
      RECT 130.58 142.44 130.78 142.56 ;
      RECT 128.78 143.7 128.98 143.82 ;
      RECT 130.22 143.7 130.42 143.82 ;
      RECT 130.94 143.7 131.14 143.82 ;
      RECT 127.34 143.46 127.54 143.58 ;
      RECT 128.06 143.46 128.26 143.58 ;
      RECT 129.5 143.46 129.7 143.58 ;
      RECT 129.5 145.98 129.7 146.1 ;
      RECT 128.78 145.98 128.98 146.1 ;
      RECT 128.06 145.98 128.26 146.1 ;
      RECT 127.7 144.96 127.9 145.08 ;
      RECT 129.86 144.96 130.06 145.08 ;
      RECT 129.14 144.96 129.34 145.08 ;
      RECT 126.98 144.72 127.18 144.84 ;
      RECT 128.42 144.72 128.62 144.84 ;
      RECT 130.58 144.72 130.78 144.84 ;
      RECT 129.86 147.24 130.06 147.36 ;
      RECT 128.42 147.24 128.62 147.36 ;
      RECT 126.98 147.24 127.18 147.36 ;
      RECT 130.94 146.22 131.14 146.34 ;
      RECT 130.22 146.22 130.42 146.34 ;
      RECT 127.34 146.22 127.54 146.34 ;
      RECT 130.22 148.74 130.42 148.86 ;
      RECT 128.78 148.74 128.98 148.86 ;
      RECT 127.34 148.74 127.54 148.86 ;
      RECT 128.06 148.5 128.26 148.62 ;
      RECT 129.5 148.5 129.7 148.62 ;
      RECT 130.94 148.5 131.14 148.62 ;
      RECT 130.58 147.48 130.78 147.6 ;
      RECT 129.14 147.48 129.34 147.6 ;
      RECT 127.7 147.48 127.9 147.6 ;
      RECT 129.86 150 130.06 150.12 ;
      RECT 126.98 150 127.18 150.12 ;
      RECT 130.58 149.76 130.78 149.88 ;
      RECT 129.14 149.76 129.34 149.88 ;
      RECT 128.42 149.76 128.62 149.88 ;
      RECT 127.7 149.76 127.9 149.88 ;
      RECT 128.78 151.26 128.98 151.38 ;
      RECT 128.06 151.26 128.26 151.38 ;
      RECT 127.34 151.26 127.54 151.38 ;
      RECT 130.94 151.02 131.14 151.14 ;
      RECT 130.22 151.02 130.42 151.14 ;
      RECT 129.5 151.02 129.7 151.14 ;
      RECT 126.98 152.28 127.18 152.4 ;
      RECT 125.54 266.2885 125.74 266.4085 ;
      RECT 126.26 266.2885 126.46 266.4085 ;
      RECT 124.1 267.81 124.3 267.93 ;
      RECT 124.82 267.81 125.02 267.93 ;
      RECT 125.54 267.81 125.74 267.93 ;
      RECT 126.26 267.81 126.46 267.93 ;
      RECT 125.18 268.2 125.38 268.32 ;
      RECT 125.9 268.2 126.1 268.32 ;
      RECT 123.74 268.44 123.94 268.56 ;
      RECT 124.46 268.44 124.66 268.56 ;
      RECT 126.62 268.44 126.82 268.56 ;
      RECT 124.1 270.09 124.3 270.21 ;
      RECT 125.54 270.09 125.74 270.21 ;
      RECT 124.82 270.33 125.02 270.45 ;
      RECT 126.26 270.33 126.46 270.45 ;
      RECT 123.74 270.72 123.94 270.84 ;
      RECT 125.18 270.72 125.38 270.84 ;
      RECT 126.62 270.72 126.82 270.84 ;
      RECT 125.9 270.96 126.1 271.08 ;
      RECT 124.46 270.96 124.66 271.08 ;
      RECT 125.54 271.35 125.74 271.47 ;
      RECT 126.26 271.35 126.46 271.47 ;
      RECT 124.1 271.59 124.3 271.71 ;
      RECT 124.82 271.59 125.02 271.71 ;
      RECT 125.9 273.48 126.1 273.6 ;
      RECT 124.46 273.48 124.66 273.6 ;
      RECT 126.62 273.24 126.82 273.36 ;
      RECT 125.18 273.24 125.38 273.36 ;
      RECT 123.74 273.24 123.94 273.36 ;
      RECT 125.9 276 126.1 276.12 ;
      RECT 124.46 276 124.66 276.12 ;
      RECT 126.62 275.76 126.82 275.88 ;
      RECT 125.18 275.76 125.38 275.88 ;
      RECT 123.74 275.76 123.94 275.88 ;
      RECT 126.62 278.28 126.82 278.4 ;
      RECT 125.18 278.28 125.38 278.4 ;
      RECT 123.74 278.28 123.94 278.4 ;
      RECT 125.9 278.52 126.1 278.64 ;
      RECT 124.46 278.52 124.66 278.64 ;
      RECT 126.26 323.3835 126.46 323.5035 ;
      RECT 125.54 323.3835 125.74 323.5035 ;
      RECT 124.82 323.3835 125.02 323.5035 ;
      RECT 124.1 323.3835 124.3 323.5035 ;
      RECT 126.26 348.339 126.46 348.459 ;
      RECT 125.54 348.339 125.74 348.459 ;
      RECT 124.82 348.339 125.02 348.459 ;
      RECT 124.1 348.339 124.3 348.459 ;
      RECT 129.86 119.52 130.06 119.64 ;
      RECT 127.7 119.52 127.9 119.64 ;
      RECT 130.58 119.76 130.78 119.88 ;
      RECT 129.14 119.76 129.34 119.88 ;
      RECT 128.42 119.76 128.62 119.88 ;
      RECT 126.98 119.76 127.18 119.88 ;
      RECT 130.22 120.78 130.42 120.9 ;
      RECT 129.5 120.78 129.7 120.9 ;
      RECT 127.34 120.78 127.54 120.9 ;
      RECT 130.94 121.02 131.14 121.14 ;
      RECT 128.78 121.02 128.98 121.14 ;
      RECT 128.06 121.02 128.26 121.14 ;
      RECT 129.86 122.04 130.06 122.16 ;
      RECT 129.14 122.04 129.34 122.16 ;
      RECT 128.42 122.04 128.62 122.16 ;
      RECT 127.7 122.04 127.9 122.16 ;
      RECT 126.98 122.28 127.18 122.4 ;
      RECT 130.58 122.28 130.78 122.4 ;
      RECT 130.22 123.3 130.42 123.42 ;
      RECT 128.78 123.3 128.98 123.42 ;
      RECT 128.06 123.3 128.26 123.42 ;
      RECT 130.94 123.54 131.14 123.66 ;
      RECT 129.5 123.54 129.7 123.66 ;
      RECT 127.34 123.54 127.54 123.66 ;
      RECT 129.14 124.56 129.34 124.68 ;
      RECT 127.7 124.56 127.9 124.68 ;
      RECT 130.58 124.8 130.78 124.92 ;
      RECT 129.86 124.8 130.06 124.92 ;
      RECT 128.42 124.8 128.62 124.92 ;
      RECT 126.98 124.8 127.18 124.92 ;
      RECT 129.5 125.82 129.7 125.94 ;
      RECT 128.06 125.82 128.26 125.94 ;
      RECT 127.34 125.82 127.54 125.94 ;
      RECT 130.94 126.06 131.14 126.18 ;
      RECT 130.22 126.06 130.42 126.18 ;
      RECT 128.78 126.06 128.98 126.18 ;
      RECT 127.7 127.08 127.9 127.2 ;
      RECT 129.86 127.08 130.06 127.2 ;
      RECT 130.58 127.08 130.78 127.2 ;
      RECT 126.98 127.32 127.18 127.44 ;
      RECT 128.42 127.32 128.62 127.44 ;
      RECT 129.14 127.32 129.34 127.44 ;
      RECT 127.34 128.34 127.54 128.46 ;
      RECT 128.78 128.34 128.98 128.46 ;
      RECT 129.5 128.34 129.7 128.46 ;
      RECT 130.22 128.34 130.42 128.46 ;
      RECT 128.06 128.58 128.26 128.7 ;
      RECT 130.94 128.58 131.14 128.7 ;
      RECT 126.98 129.6 127.18 129.72 ;
      RECT 127.7 129.6 127.9 129.72 ;
      RECT 129.14 129.6 129.34 129.72 ;
      RECT 130.58 129.84 130.78 129.96 ;
      RECT 129.86 129.84 130.06 129.96 ;
      RECT 128.42 129.84 128.62 129.96 ;
      RECT 128.78 130.86 128.98 130.98 ;
      RECT 124.82 195.12 125.02 195.24 ;
      RECT 126.26 195.12 126.46 195.24 ;
      RECT 125.54 195.36 125.74 195.48 ;
      RECT 124.1 195.36 124.3 195.48 ;
      RECT 124.82 197.88 125.02 198 ;
      RECT 126.26 197.88 126.46 198 ;
      RECT 125.54 197.64 125.74 197.76 ;
      RECT 124.1 197.64 124.3 197.76 ;
      RECT 124.82 200.4 125.02 200.52 ;
      RECT 126.26 200.16 126.46 200.28 ;
      RECT 125.54 200.16 125.74 200.28 ;
      RECT 124.1 200.16 124.3 200.28 ;
      RECT 124.82 202.92 125.02 203.04 ;
      RECT 124.1 202.92 124.3 203.04 ;
      RECT 125.54 202.68 125.74 202.8 ;
      RECT 126.26 202.68 126.46 202.8 ;
      RECT 124.82 205.44 125.02 205.56 ;
      RECT 124.1 205.2 124.3 205.32 ;
      RECT 125.54 205.2 125.74 205.32 ;
      RECT 126.26 205.2 126.46 205.32 ;
      RECT 124.82 207.96 125.02 208.08 ;
      RECT 124.1 207.72 124.3 207.84 ;
      RECT 125.54 207.72 125.74 207.84 ;
      RECT 126.26 207.72 126.46 207.84 ;
      RECT 125.54 210.48 125.74 210.6 ;
      RECT 124.1 210.24 124.3 210.36 ;
      RECT 124.82 210.24 125.02 210.36 ;
      RECT 126.26 210.24 126.46 210.36 ;
      RECT 124.1 212.76 124.3 212.88 ;
      RECT 124.82 212.76 125.02 212.88 ;
      RECT 126.26 212.76 126.46 212.88 ;
      RECT 125.54 213 125.74 213.12 ;
      RECT 124.82 215.52 125.02 215.64 ;
      RECT 126.26 215.52 126.46 215.64 ;
      RECT 124.1 215.28 124.3 215.4 ;
      RECT 125.54 215.28 125.74 215.4 ;
      RECT 123.74 222.362 123.94 222.482 ;
      RECT 124.46 222.362 124.66 222.482 ;
      RECT 125.18 222.122 125.38 222.242 ;
      RECT 125.9 222.122 126.1 222.242 ;
      RECT 126.62 222.122 126.82 222.242 ;
      RECT 124.1 223.08 124.3 223.2 ;
      RECT 124.82 223.08 125.02 223.2 ;
      RECT 125.54 222.84 125.74 222.96 ;
      RECT 126.26 222.84 126.46 222.96 ;
      RECT 123.74 250.56 123.94 250.68 ;
      RECT 124.46 250.56 124.66 250.68 ;
      RECT 125.18 250.56 125.38 250.68 ;
      RECT 125.9 250.8 126.1 250.92 ;
      RECT 126.62 250.8 126.82 250.92 ;
      RECT 123.74 253.08 123.94 253.2 ;
      RECT 125.18 253.08 125.38 253.2 ;
      RECT 125.9 253.08 126.1 253.2 ;
      RECT 126.62 253.08 126.82 253.2 ;
      RECT 124.46 253.32 124.66 253.44 ;
      RECT 123.74 255.6 123.94 255.72 ;
      RECT 124.46 255.6 124.66 255.72 ;
      RECT 125.18 255.6 125.38 255.72 ;
      RECT 126.62 255.6 126.82 255.72 ;
      RECT 125.9 255.84 126.1 255.96 ;
      RECT 123.74 258.12 123.94 258.24 ;
      RECT 125.18 258.12 125.38 258.24 ;
      RECT 126.62 258.12 126.82 258.24 ;
      RECT 124.46 258.36 124.66 258.48 ;
      RECT 125.9 258.36 126.1 258.48 ;
      RECT 124.1 258.75 124.3 258.87 ;
      RECT 124.82 258.99 125.02 259.11 ;
      RECT 125.54 258.99 125.74 259.11 ;
      RECT 126.26 258.99 126.46 259.11 ;
      RECT 124.1 260.01 124.3 260.13 ;
      RECT 124.82 260.01 125.02 260.13 ;
      RECT 125.54 260.01 125.74 260.13 ;
      RECT 126.26 260.25 126.46 260.37 ;
      RECT 123.74 260.64 123.94 260.76 ;
      RECT 125.18 260.64 125.38 260.76 ;
      RECT 126.62 260.64 126.82 260.76 ;
      RECT 124.46 260.88 124.66 261 ;
      RECT 125.9 260.88 126.1 261 ;
      RECT 125.54 261.27 125.74 261.39 ;
      RECT 124.1 261.51 124.3 261.63 ;
      RECT 124.82 261.51 125.02 261.63 ;
      RECT 126.26 261.51 126.46 261.63 ;
      RECT 124.1 262.53 124.3 262.65 ;
      RECT 125.54 262.53 125.74 262.65 ;
      RECT 124.82 262.77 125.02 262.89 ;
      RECT 126.26 262.77 126.46 262.89 ;
      RECT 123.74 263.16 123.94 263.28 ;
      RECT 124.46 263.16 124.66 263.28 ;
      RECT 126.62 263.16 126.82 263.28 ;
      RECT 125.18 263.4 125.38 263.52 ;
      RECT 125.9 263.4 126.1 263.52 ;
      RECT 124.1 263.79 124.3 263.91 ;
      RECT 125.54 263.79 125.74 263.91 ;
      RECT 126.26 263.79 126.46 263.91 ;
      RECT 124.82 264.03 125.02 264.15 ;
      RECT 123.74 265.68 123.94 265.8 ;
      RECT 125.18 265.68 125.38 265.8 ;
      RECT 126.62 265.68 126.82 265.8 ;
      RECT 124.46 265.92 124.66 266.04 ;
      RECT 125.9 265.92 126.1 266.04 ;
      RECT 124.1 266.2885 124.3 266.4085 ;
      RECT 124.82 266.2885 125.02 266.4085 ;
      RECT 123.74 163.62 123.94 163.74 ;
      RECT 124.46 163.62 124.66 163.74 ;
      RECT 125.9 163.62 126.1 163.74 ;
      RECT 125.18 163.86 125.38 163.98 ;
      RECT 124.1 164.88 124.3 165 ;
      RECT 125.54 164.88 125.74 165 ;
      RECT 126.26 164.88 126.46 165 ;
      RECT 124.82 165.12 125.02 165.24 ;
      RECT 125.9 166.14 126.1 166.26 ;
      RECT 125.18 166.14 125.38 166.26 ;
      RECT 124.46 166.14 124.66 166.26 ;
      RECT 123.74 166.14 123.94 166.26 ;
      RECT 126.62 166.38 126.82 166.5 ;
      RECT 125.54 167.4 125.74 167.52 ;
      RECT 124.1 167.64 124.3 167.76 ;
      RECT 124.82 167.64 125.02 167.76 ;
      RECT 126.26 167.64 126.46 167.76 ;
      RECT 126.62 168.66 126.82 168.78 ;
      RECT 125.18 168.66 125.38 168.78 ;
      RECT 123.74 168.66 123.94 168.78 ;
      RECT 124.46 168.9 124.66 169.02 ;
      RECT 125.9 168.9 126.1 169.02 ;
      RECT 124.1 169.92 124.3 170.04 ;
      RECT 124.82 169.92 125.02 170.04 ;
      RECT 125.54 169.92 125.74 170.04 ;
      RECT 126.26 169.92 126.46 170.04 ;
      RECT 124.46 171.18 124.66 171.3 ;
      RECT 125.18 171.18 125.38 171.3 ;
      RECT 125.9 171.18 126.1 171.3 ;
      RECT 126.62 171.18 126.82 171.3 ;
      RECT 123.74 171.42 123.94 171.54 ;
      RECT 125.54 172.44 125.74 172.56 ;
      RECT 124.1 172.44 124.3 172.56 ;
      RECT 124.82 172.68 125.02 172.8 ;
      RECT 126.26 172.68 126.46 172.8 ;
      RECT 124.46 173.7 124.66 173.82 ;
      RECT 125.9 173.7 126.1 173.82 ;
      RECT 126.62 173.7 126.82 173.82 ;
      RECT 123.74 173.94 123.94 174.06 ;
      RECT 125.18 173.94 125.38 174.06 ;
      RECT 126.26 174.96 126.46 175.08 ;
      RECT 125.54 174.96 125.74 175.08 ;
      RECT 124.1 174.96 124.3 175.08 ;
      RECT 124.82 175.2 125.02 175.32 ;
      RECT 123.74 176.22 123.94 176.34 ;
      RECT 124.46 176.22 124.66 176.34 ;
      RECT 125.18 176.22 125.38 176.34 ;
      RECT 125.9 176.22 126.1 176.34 ;
      RECT 126.62 176.22 126.82 176.34 ;
      RECT 124.82 177.72 125.02 177.84 ;
      RECT 126.62 178.74 126.82 178.86 ;
      RECT 125.9 178.74 126.1 178.86 ;
      RECT 125.18 178.74 125.38 178.86 ;
      RECT 124.46 178.74 124.66 178.86 ;
      RECT 123.74 178.74 123.94 178.86 ;
      RECT 124.1 177.48 124.3 177.6 ;
      RECT 125.54 177.48 125.74 177.6 ;
      RECT 126.26 177.48 126.46 177.6 ;
      RECT 125.54 180 125.74 180.12 ;
      RECT 126.26 180 126.46 180.12 ;
      RECT 123.74 181.26 123.94 181.38 ;
      RECT 124.46 181.26 124.66 181.38 ;
      RECT 125.18 181.26 125.38 181.38 ;
      RECT 125.9 181.26 126.1 181.38 ;
      RECT 126.62 181.26 126.82 181.38 ;
      RECT 124.82 180.24 125.02 180.36 ;
      RECT 124.1 180.24 124.3 180.36 ;
      RECT 124.82 182.76 125.02 182.88 ;
      RECT 126.26 182.52 126.46 182.64 ;
      RECT 125.54 182.52 125.74 182.64 ;
      RECT 124.1 182.52 124.3 182.64 ;
      RECT 123.74 184.02 123.94 184.14 ;
      RECT 126.62 183.78 126.82 183.9 ;
      RECT 125.9 183.78 126.1 183.9 ;
      RECT 125.18 183.78 125.38 183.9 ;
      RECT 124.46 183.78 124.66 183.9 ;
      RECT 124.82 185.28 125.02 185.4 ;
      RECT 126.26 185.04 126.46 185.16 ;
      RECT 125.54 185.04 125.74 185.16 ;
      RECT 124.1 185.04 124.3 185.16 ;
      RECT 123.74 186.3 123.94 186.42 ;
      RECT 126.62 186.3 126.82 186.42 ;
      RECT 125.9 186.3 126.1 186.42 ;
      RECT 125.18 186.3 125.38 186.42 ;
      RECT 124.46 186.3 124.66 186.42 ;
      RECT 124.82 187.8 125.02 187.92 ;
      RECT 126.26 187.56 126.46 187.68 ;
      RECT 125.54 187.56 125.74 187.68 ;
      RECT 124.1 187.56 124.3 187.68 ;
      RECT 124.46 189.06 124.66 189.18 ;
      RECT 125.18 189.06 125.38 189.18 ;
      RECT 126.62 188.82 126.82 188.94 ;
      RECT 125.9 188.82 126.1 188.94 ;
      RECT 123.74 188.82 123.94 188.94 ;
      RECT 124.82 190.32 125.02 190.44 ;
      RECT 126.26 190.08 126.46 190.2 ;
      RECT 125.54 190.08 125.74 190.2 ;
      RECT 124.1 190.08 124.3 190.2 ;
      RECT 125.54 192.84 125.74 192.96 ;
      RECT 124.1 192.84 124.3 192.96 ;
      RECT 124.82 192.6 125.02 192.72 ;
      RECT 126.26 192.6 126.46 192.72 ;
      RECT 123.74 131.1 123.94 131.22 ;
      RECT 124.82 132.12 125.02 132.24 ;
      RECT 125.54 132.12 125.74 132.24 ;
      RECT 126.26 132.12 126.46 132.24 ;
      RECT 124.1 132.36 124.3 132.48 ;
      RECT 125.9 133.38 126.1 133.5 ;
      RECT 124.46 133.38 124.66 133.5 ;
      RECT 123.74 133.62 123.94 133.74 ;
      RECT 125.18 133.62 125.38 133.74 ;
      RECT 126.62 133.62 126.82 133.74 ;
      RECT 124.1 134.64 124.3 134.76 ;
      RECT 124.82 134.64 125.02 134.76 ;
      RECT 126.26 134.64 126.46 134.76 ;
      RECT 125.54 134.88 125.74 135 ;
      RECT 123.74 135.9 123.94 136.02 ;
      RECT 125.18 135.9 125.38 136.02 ;
      RECT 126.62 135.9 126.82 136.02 ;
      RECT 125.9 136.14 126.1 136.26 ;
      RECT 124.46 136.14 124.66 136.26 ;
      RECT 125.54 137.16 125.74 137.28 ;
      RECT 124.82 137.16 125.02 137.28 ;
      RECT 126.26 137.4 126.46 137.52 ;
      RECT 124.1 137.4 124.3 137.52 ;
      RECT 123.74 138.42 123.94 138.54 ;
      RECT 125.18 138.42 125.38 138.54 ;
      RECT 126.62 138.42 126.82 138.54 ;
      RECT 124.46 138.66 124.66 138.78 ;
      RECT 125.9 138.66 126.1 138.78 ;
      RECT 124.82 139.68 125.02 139.8 ;
      RECT 126.26 139.68 126.46 139.8 ;
      RECT 124.1 139.92 124.3 140.04 ;
      RECT 125.54 139.92 125.74 140.04 ;
      RECT 125.9 140.94 126.1 141.06 ;
      RECT 125.18 140.94 125.38 141.06 ;
      RECT 124.46 140.94 124.66 141.06 ;
      RECT 123.74 140.94 123.94 141.06 ;
      RECT 126.62 141.18 126.82 141.3 ;
      RECT 124.1 142.2 124.3 142.32 ;
      RECT 124.82 142.2 125.02 142.32 ;
      RECT 125.54 142.2 125.74 142.32 ;
      RECT 125.9 143.46 126.1 143.58 ;
      RECT 125.18 143.46 125.38 143.58 ;
      RECT 124.46 143.46 124.66 143.58 ;
      RECT 123.74 143.46 123.94 143.58 ;
      RECT 126.62 143.46 126.82 143.58 ;
      RECT 123.74 145.98 123.94 146.1 ;
      RECT 124.46 145.98 124.66 146.1 ;
      RECT 125.18 145.98 125.38 146.1 ;
      RECT 125.9 145.98 126.1 146.1 ;
      RECT 124.82 144.96 125.02 145.08 ;
      RECT 124.1 144.72 124.3 144.84 ;
      RECT 125.54 144.72 125.74 144.84 ;
      RECT 126.62 146.22 126.82 146.34 ;
      RECT 125.9 148.74 126.1 148.86 ;
      RECT 124.46 148.74 124.66 148.86 ;
      RECT 123.74 148.5 123.94 148.62 ;
      RECT 125.18 148.5 125.38 148.62 ;
      RECT 126.62 148.5 126.82 148.62 ;
      RECT 124.1 150 124.3 150.12 ;
      RECT 126.26 149.76 126.46 149.88 ;
      RECT 125.54 149.76 125.74 149.88 ;
      RECT 124.82 149.76 125.02 149.88 ;
      RECT 125.18 151.26 125.38 151.38 ;
      RECT 126.62 151.02 126.82 151.14 ;
      RECT 125.9 151.02 126.1 151.14 ;
      RECT 124.46 151.02 124.66 151.14 ;
      RECT 123.74 151.02 123.94 151.14 ;
      RECT 125.54 152.28 125.74 152.4 ;
      RECT 126.26 152.28 126.46 152.4 ;
      RECT 124.1 152.28 124.3 152.4 ;
      RECT 124.82 152.52 125.02 152.64 ;
      RECT 126.62 153.54 126.82 153.66 ;
      RECT 125.18 153.54 125.38 153.66 ;
      RECT 123.74 153.54 123.94 153.66 ;
      RECT 124.46 153.78 124.66 153.9 ;
      RECT 125.9 153.78 126.1 153.9 ;
      RECT 124.82 154.8 125.02 154.92 ;
      RECT 124.1 155.04 124.3 155.16 ;
      RECT 125.54 155.04 125.74 155.16 ;
      RECT 126.26 155.04 126.46 155.16 ;
      RECT 125.9 156.06 126.1 156.18 ;
      RECT 124.46 156.06 124.66 156.18 ;
      RECT 126.62 156.06 126.82 156.18 ;
      RECT 123.74 156.3 123.94 156.42 ;
      RECT 125.18 156.3 125.38 156.42 ;
      RECT 124.1 157.32 124.3 157.44 ;
      RECT 124.82 157.32 125.02 157.44 ;
      RECT 125.54 157.32 125.74 157.44 ;
      RECT 126.26 157.32 126.46 157.44 ;
      RECT 125.9 158.58 126.1 158.7 ;
      RECT 124.46 158.58 124.66 158.7 ;
      RECT 123.74 158.82 123.94 158.94 ;
      RECT 125.18 158.82 125.38 158.94 ;
      RECT 124.1 159.84 124.3 159.96 ;
      RECT 125.54 159.84 125.74 159.96 ;
      RECT 126.26 159.84 126.46 159.96 ;
      RECT 124.82 160.08 125.02 160.2 ;
      RECT 126.62 161.1 126.82 161.22 ;
      RECT 125.9 161.1 126.1 161.22 ;
      RECT 125.18 161.1 125.38 161.22 ;
      RECT 124.46 161.1 124.66 161.22 ;
      RECT 123.74 161.1 123.94 161.22 ;
      RECT 113.3 267.81 113.5 267.93 ;
      RECT 112.58 267.81 112.78 267.93 ;
      RECT 111.14 270.09 111.34 270.21 ;
      RECT 110.78 269.7 110.98 269.82 ;
      RECT 111.5 269.46 111.7 269.58 ;
      RECT 114.02 270.09 114.22 270.21 ;
      RECT 112.58 270.09 112.78 270.21 ;
      RECT 114.38 269.7 114.58 269.82 ;
      RECT 112.94 269.7 113.14 269.82 ;
      RECT 113.66 269.46 113.86 269.58 ;
      RECT 112.22 269.46 112.42 269.58 ;
      RECT 111.86 271.35 112.06 271.47 ;
      RECT 111.14 271.35 111.34 271.47 ;
      RECT 111.86 270.33 112.06 270.45 ;
      RECT 114.02 271.59 114.22 271.71 ;
      RECT 112.58 271.59 112.78 271.71 ;
      RECT 113.3 271.35 113.5 271.47 ;
      RECT 113.3 270.33 113.5 270.45 ;
      RECT 111.5 272.22 111.7 272.34 ;
      RECT 110.78 271.98 110.98 272.1 ;
      RECT 112.94 271.98 113.14 272.1 ;
      RECT 112.22 272.22 112.42 272.34 ;
      RECT 113.66 272.22 113.86 272.34 ;
      RECT 114.38 272.22 114.58 272.34 ;
      RECT 110.78 274.74 110.98 274.86 ;
      RECT 111.5 274.5 111.7 274.62 ;
      RECT 112.22 274.5 112.42 274.62 ;
      RECT 114.38 274.5 114.58 274.62 ;
      RECT 112.94 274.74 113.14 274.86 ;
      RECT 113.66 274.74 113.86 274.86 ;
      RECT 110.78 277.02 110.98 277.14 ;
      RECT 112.94 277.02 113.14 277.14 ;
      RECT 114.38 277.02 114.58 277.14 ;
      RECT 111.5 277.26 111.7 277.38 ;
      RECT 112.22 277.26 112.42 277.38 ;
      RECT 113.66 277.26 113.86 277.38 ;
      RECT 112.22 308.496 112.42 308.616 ;
      RECT 112.94 308.496 113.14 308.616 ;
      RECT 113.66 308.496 113.86 308.616 ;
      RECT 114.38 308.496 114.58 308.616 ;
      RECT 110.78 308.496 110.98 308.616 ;
      RECT 111.5 308.496 111.7 308.616 ;
      RECT 114.02 323.3835 114.22 323.5035 ;
      RECT 113.3 323.3835 113.5 323.5035 ;
      RECT 112.58 323.3835 112.78 323.5035 ;
      RECT 111.14 323.3835 111.34 323.5035 ;
      RECT 111.86 323.3835 112.06 323.5035 ;
      RECT 114.38 325.9425 114.58 326.0625 ;
      RECT 113.66 325.9425 113.86 326.0625 ;
      RECT 112.94 325.9425 113.14 326.0625 ;
      RECT 112.22 325.9425 112.42 326.0625 ;
      RECT 110.78 325.9425 110.98 326.0625 ;
      RECT 111.5 325.9425 111.7 326.0625 ;
      RECT 114.02 348.339 114.22 348.459 ;
      RECT 113.3 348.339 113.5 348.459 ;
      RECT 112.58 348.339 112.78 348.459 ;
      RECT 111.14 348.339 111.34 348.459 ;
      RECT 111.86 348.339 112.06 348.459 ;
      RECT 126.26 119.52 126.46 119.64 ;
      RECT 125.54 119.52 125.74 119.64 ;
      RECT 124.82 119.52 125.02 119.64 ;
      RECT 124.1 119.76 124.3 119.88 ;
      RECT 126.62 120.78 126.82 120.9 ;
      RECT 125.18 120.78 125.38 120.9 ;
      RECT 125.9 121.02 126.1 121.14 ;
      RECT 124.46 121.02 124.66 121.14 ;
      RECT 123.74 121.02 123.94 121.14 ;
      RECT 126.26 122.04 126.46 122.16 ;
      RECT 125.54 122.04 125.74 122.16 ;
      RECT 124.82 122.04 125.02 122.16 ;
      RECT 124.1 122.28 124.3 122.4 ;
      RECT 125.9 123.3 126.1 123.42 ;
      RECT 123.74 123.3 123.94 123.42 ;
      RECT 126.62 123.54 126.82 123.66 ;
      RECT 125.18 123.54 125.38 123.66 ;
      RECT 124.46 123.54 124.66 123.66 ;
      RECT 126.26 124.56 126.46 124.68 ;
      RECT 125.54 124.56 125.74 124.68 ;
      RECT 124.82 124.56 125.02 124.68 ;
      RECT 124.1 124.8 124.3 124.92 ;
      RECT 125.9 125.82 126.1 125.94 ;
      RECT 124.46 125.82 124.66 125.94 ;
      RECT 126.62 126.06 126.82 126.18 ;
      RECT 125.18 126.06 125.38 126.18 ;
      RECT 123.74 126.06 123.94 126.18 ;
      RECT 124.82 127.08 125.02 127.2 ;
      RECT 125.54 127.08 125.74 127.2 ;
      RECT 126.26 127.08 126.46 127.2 ;
      RECT 124.1 127.32 124.3 127.44 ;
      RECT 124.46 128.34 124.66 128.46 ;
      RECT 125.18 128.34 125.38 128.46 ;
      RECT 125.9 128.34 126.1 128.46 ;
      RECT 123.74 128.58 123.94 128.7 ;
      RECT 126.62 128.58 126.82 128.7 ;
      RECT 124.1 129.6 124.3 129.72 ;
      RECT 126.26 129.6 126.46 129.72 ;
      RECT 125.54 129.84 125.74 129.96 ;
      RECT 124.82 129.84 125.02 129.96 ;
      RECT 125.9 130.86 126.1 130.98 ;
      RECT 126.62 130.86 126.82 130.98 ;
      RECT 125.18 131.1 125.38 131.22 ;
      RECT 124.46 131.1 124.66 131.22 ;
      RECT 112.22 239.46 112.42 239.58 ;
      RECT 114.38 239.22 114.58 239.34 ;
      RECT 112.94 239.22 113.14 239.34 ;
      RECT 110.78 241.98 110.98 242.1 ;
      RECT 111.5 241.74 111.7 241.86 ;
      RECT 112.22 241.98 112.42 242.1 ;
      RECT 114.38 241.98 114.58 242.1 ;
      RECT 112.94 241.74 113.14 241.86 ;
      RECT 113.66 241.74 113.86 241.86 ;
      RECT 111.5 244.26 111.7 244.38 ;
      RECT 114.38 244.26 114.58 244.38 ;
      RECT 112.94 244.26 113.14 244.38 ;
      RECT 110.78 244.5 110.98 244.62 ;
      RECT 112.22 244.5 112.42 244.62 ;
      RECT 113.66 244.5 113.86 244.62 ;
      RECT 110.78 247.02 110.98 247.14 ;
      RECT 111.5 246.78 111.7 246.9 ;
      RECT 113.66 247.02 113.86 247.14 ;
      RECT 112.22 247.02 112.42 247.14 ;
      RECT 114.38 246.78 114.58 246.9 ;
      RECT 112.94 246.78 113.14 246.9 ;
      RECT 110.78 249.54 110.98 249.66 ;
      RECT 111.5 249.3 111.7 249.42 ;
      RECT 113.66 249.54 113.86 249.66 ;
      RECT 112.22 249.54 112.42 249.66 ;
      RECT 114.38 249.3 114.58 249.42 ;
      RECT 112.94 249.3 113.14 249.42 ;
      RECT 110.78 252.06 110.98 252.18 ;
      RECT 111.5 251.82 111.7 251.94 ;
      RECT 113.66 252.06 113.86 252.18 ;
      RECT 112.22 252.06 112.42 252.18 ;
      RECT 114.38 251.82 114.58 251.94 ;
      RECT 112.94 251.82 113.14 251.94 ;
      RECT 111.5 254.58 111.7 254.7 ;
      RECT 110.78 254.34 110.98 254.46 ;
      RECT 113.66 254.58 113.86 254.7 ;
      RECT 112.22 254.58 112.42 254.7 ;
      RECT 114.38 254.34 114.58 254.46 ;
      RECT 112.94 254.34 113.14 254.46 ;
      RECT 111.5 256.86 111.7 256.98 ;
      RECT 110.78 256.86 110.98 256.98 ;
      RECT 113.66 257.1 113.86 257.22 ;
      RECT 112.22 257.1 112.42 257.22 ;
      RECT 114.38 256.86 114.58 256.98 ;
      RECT 112.94 256.86 113.14 256.98 ;
      RECT 111.86 258.99 112.06 259.11 ;
      RECT 111.14 258.99 111.34 259.11 ;
      RECT 113.3 258.99 113.5 259.11 ;
      RECT 114.02 258.75 114.22 258.87 ;
      RECT 112.58 258.75 112.78 258.87 ;
      RECT 111.86 260.25 112.06 260.37 ;
      RECT 111.14 260.25 111.34 260.37 ;
      RECT 111.5 259.38 111.7 259.5 ;
      RECT 110.78 259.38 110.98 259.5 ;
      RECT 114.02 260.25 114.22 260.37 ;
      RECT 113.3 260.25 113.5 260.37 ;
      RECT 112.58 260.01 112.78 260.13 ;
      RECT 113.66 259.62 113.86 259.74 ;
      RECT 112.22 259.62 112.42 259.74 ;
      RECT 114.38 259.38 114.58 259.5 ;
      RECT 112.94 259.38 113.14 259.5 ;
      RECT 111.5 261.9 111.7 262.02 ;
      RECT 111.86 261.51 112.06 261.63 ;
      RECT 111.14 261.27 111.34 261.39 ;
      RECT 114.38 261.9 114.58 262.02 ;
      RECT 112.94 261.9 113.14 262.02 ;
      RECT 113.3 261.51 113.5 261.63 ;
      RECT 114.02 261.27 114.22 261.39 ;
      RECT 112.58 261.27 112.78 261.39 ;
      RECT 111.86 262.77 112.06 262.89 ;
      RECT 111.14 262.53 111.34 262.65 ;
      RECT 110.78 262.14 110.98 262.26 ;
      RECT 114.02 262.77 114.22 262.89 ;
      RECT 113.3 262.53 113.5 262.65 ;
      RECT 112.58 262.53 112.78 262.65 ;
      RECT 113.66 262.14 113.86 262.26 ;
      RECT 112.22 262.14 112.42 262.26 ;
      RECT 110.78 264.66 110.98 264.78 ;
      RECT 111.5 264.42 111.7 264.54 ;
      RECT 111.86 264.03 112.06 264.15 ;
      RECT 111.14 263.79 111.34 263.91 ;
      RECT 113.66 264.66 113.86 264.78 ;
      RECT 112.94 264.66 113.14 264.78 ;
      RECT 114.38 264.42 114.58 264.54 ;
      RECT 112.22 264.42 112.42 264.54 ;
      RECT 113.3 264.03 113.5 264.15 ;
      RECT 114.02 263.79 114.22 263.91 ;
      RECT 112.58 263.79 112.78 263.91 ;
      RECT 111.5 267.18 111.7 267.3 ;
      RECT 110.78 267.18 110.98 267.3 ;
      RECT 111.86 266.2885 112.06 266.4085 ;
      RECT 111.14 266.2885 111.34 266.4085 ;
      RECT 112.94 267.18 113.14 267.3 ;
      RECT 112.22 267.18 112.42 267.3 ;
      RECT 114.38 266.94 114.58 267.06 ;
      RECT 113.66 266.94 113.86 267.06 ;
      RECT 114.02 266.2885 114.22 266.4085 ;
      RECT 113.3 266.2885 113.5 266.4085 ;
      RECT 112.58 266.2885 112.78 266.4085 ;
      RECT 111.86 267.81 112.06 267.93 ;
      RECT 111.14 267.81 111.34 267.93 ;
      RECT 114.02 267.81 114.22 267.93 ;
      RECT 112.22 204.18 112.42 204.3 ;
      RECT 110.78 203.94 110.98 204.06 ;
      RECT 111.5 203.94 111.7 204.06 ;
      RECT 112.58 205.2 112.78 205.32 ;
      RECT 114.02 205.2 114.22 205.32 ;
      RECT 113.3 205.44 113.5 205.56 ;
      RECT 111.86 205.2 112.06 205.32 ;
      RECT 111.14 205.44 111.34 205.56 ;
      RECT 112.94 206.46 113.14 206.58 ;
      RECT 114.38 206.46 114.58 206.58 ;
      RECT 113.66 206.7 113.86 206.82 ;
      RECT 112.22 206.7 112.42 206.82 ;
      RECT 110.78 206.46 110.98 206.58 ;
      RECT 111.5 206.46 111.7 206.58 ;
      RECT 113.3 207.72 113.5 207.84 ;
      RECT 114.02 207.96 114.22 208.08 ;
      RECT 112.58 207.96 112.78 208.08 ;
      RECT 111.14 207.72 111.34 207.84 ;
      RECT 111.86 207.96 112.06 208.08 ;
      RECT 113.66 208.98 113.86 209.1 ;
      RECT 114.38 208.98 114.58 209.1 ;
      RECT 112.22 209.22 112.42 209.34 ;
      RECT 112.94 209.22 113.14 209.34 ;
      RECT 110.78 209.22 110.98 209.34 ;
      RECT 111.5 209.22 111.7 209.34 ;
      RECT 113.3 210.48 113.5 210.6 ;
      RECT 112.94 211.5 113.14 211.62 ;
      RECT 111.86 210.48 112.06 210.6 ;
      RECT 111.5 211.5 111.7 211.62 ;
      RECT 114.02 210.24 114.22 210.36 ;
      RECT 112.58 210.24 112.78 210.36 ;
      RECT 111.14 210.24 111.34 210.36 ;
      RECT 112.22 211.74 112.42 211.86 ;
      RECT 113.66 211.74 113.86 211.86 ;
      RECT 114.38 211.74 114.58 211.86 ;
      RECT 113.3 212.76 113.5 212.88 ;
      RECT 112.58 212.76 112.78 212.88 ;
      RECT 110.78 211.74 110.98 211.86 ;
      RECT 114.02 213 114.22 213.12 ;
      RECT 112.94 214.02 113.14 214.14 ;
      RECT 114.38 214.02 114.58 214.14 ;
      RECT 112.22 214.26 112.42 214.38 ;
      RECT 113.66 214.26 113.86 214.38 ;
      RECT 111.14 213 111.34 213.12 ;
      RECT 111.86 213 112.06 213.12 ;
      RECT 111.5 214.02 111.7 214.14 ;
      RECT 110.78 214.26 110.98 214.38 ;
      RECT 114.02 215.28 114.22 215.4 ;
      RECT 113.3 215.52 113.5 215.64 ;
      RECT 112.58 215.52 112.78 215.64 ;
      RECT 111.86 215.28 112.06 215.4 ;
      RECT 111.14 215.52 111.34 215.64 ;
      RECT 112.94 216.54 113.14 216.66 ;
      RECT 114.38 216.54 114.58 216.66 ;
      RECT 112.22 216.78 112.42 216.9 ;
      RECT 113.66 216.78 113.86 216.9 ;
      RECT 110.78 216.54 110.98 216.66 ;
      RECT 111.5 216.78 111.7 216.9 ;
      RECT 110.78 219.3 110.98 219.42 ;
      RECT 112.94 219.06 113.14 219.18 ;
      RECT 114.38 219.06 114.58 219.18 ;
      RECT 112.22 219.3 112.42 219.42 ;
      RECT 113.66 219.3 113.86 219.42 ;
      RECT 111.5 219.06 111.7 219.18 ;
      RECT 110.78 223.798 110.98 223.918 ;
      RECT 111.5 223.558 111.7 223.678 ;
      RECT 111.86 223.08 112.06 223.2 ;
      RECT 111.14 222.84 111.34 222.96 ;
      RECT 112.22 223.798 112.42 223.918 ;
      RECT 112.94 223.798 113.14 223.918 ;
      RECT 113.66 223.558 113.86 223.678 ;
      RECT 114.38 223.558 114.58 223.678 ;
      RECT 113.3 223.08 113.5 223.2 ;
      RECT 112.58 222.84 112.78 222.96 ;
      RECT 114.02 222.84 114.22 222.96 ;
      RECT 112.94 229.14 113.14 229.26 ;
      RECT 114.38 229.14 114.58 229.26 ;
      RECT 110.78 229.38 110.98 229.5 ;
      RECT 111.5 229.38 111.7 229.5 ;
      RECT 112.22 229.38 112.42 229.5 ;
      RECT 113.66 229.38 113.86 229.5 ;
      RECT 110.78 231.9 110.98 232.02 ;
      RECT 111.5 231.66 111.7 231.78 ;
      RECT 113.66 231.9 113.86 232.02 ;
      RECT 112.94 231.9 113.14 232.02 ;
      RECT 112.22 231.66 112.42 231.78 ;
      RECT 114.38 231.66 114.58 231.78 ;
      RECT 111.5 234.42 111.7 234.54 ;
      RECT 110.78 234.18 110.98 234.3 ;
      RECT 114.38 234.42 114.58 234.54 ;
      RECT 112.22 234.42 112.42 234.54 ;
      RECT 112.94 234.18 113.14 234.3 ;
      RECT 113.66 234.18 113.86 234.3 ;
      RECT 110.78 236.94 110.98 237.06 ;
      RECT 111.5 236.94 111.7 237.06 ;
      RECT 112.22 236.94 112.42 237.06 ;
      RECT 112.94 236.94 113.14 237.06 ;
      RECT 113.66 236.7 113.86 236.82 ;
      RECT 114.38 236.7 114.58 236.82 ;
      RECT 110.78 239.46 110.98 239.58 ;
      RECT 111.5 239.22 111.7 239.34 ;
      RECT 113.66 239.46 113.86 239.58 ;
      RECT 112.22 181.26 112.42 181.38 ;
      RECT 113.66 181.26 113.86 181.38 ;
      RECT 114.38 181.26 114.58 181.38 ;
      RECT 110.78 181.5 110.98 181.62 ;
      RECT 111.5 181.26 111.7 181.38 ;
      RECT 111.86 180.24 112.06 180.36 ;
      RECT 113.3 182.76 113.5 182.88 ;
      RECT 114.02 182.52 114.22 182.64 ;
      RECT 112.58 182.52 112.78 182.64 ;
      RECT 111.14 182.76 111.34 182.88 ;
      RECT 111.86 182.52 112.06 182.64 ;
      RECT 114.38 184.02 114.58 184.14 ;
      RECT 113.66 184.02 113.86 184.14 ;
      RECT 112.22 184.02 112.42 184.14 ;
      RECT 112.94 183.78 113.14 183.9 ;
      RECT 111.5 183.78 111.7 183.9 ;
      RECT 110.78 183.78 110.98 183.9 ;
      RECT 112.58 185.28 112.78 185.4 ;
      RECT 113.3 185.28 113.5 185.4 ;
      RECT 114.02 185.04 114.22 185.16 ;
      RECT 111.86 185.04 112.06 185.16 ;
      RECT 111.14 185.04 111.34 185.16 ;
      RECT 113.66 186.54 113.86 186.66 ;
      RECT 114.38 186.3 114.58 186.42 ;
      RECT 112.94 186.3 113.14 186.42 ;
      RECT 112.22 186.3 112.42 186.42 ;
      RECT 110.78 186.54 110.98 186.66 ;
      RECT 111.5 186.3 111.7 186.42 ;
      RECT 112.58 187.8 112.78 187.92 ;
      RECT 114.02 187.56 114.22 187.68 ;
      RECT 113.3 187.56 113.5 187.68 ;
      RECT 111.86 187.8 112.06 187.92 ;
      RECT 111.14 187.8 111.34 187.92 ;
      RECT 112.94 189.06 113.14 189.18 ;
      RECT 114.38 188.82 114.58 188.94 ;
      RECT 113.66 188.82 113.86 188.94 ;
      RECT 112.22 188.82 112.42 188.94 ;
      RECT 111.5 189.06 111.7 189.18 ;
      RECT 110.78 188.82 110.98 188.94 ;
      RECT 114.02 190.32 114.22 190.44 ;
      RECT 113.3 190.08 113.5 190.2 ;
      RECT 112.58 190.08 112.78 190.2 ;
      RECT 111.14 190.32 111.34 190.44 ;
      RECT 111.86 190.32 112.06 190.44 ;
      RECT 114.38 191.58 114.58 191.7 ;
      RECT 113.66 191.58 113.86 191.7 ;
      RECT 112.22 191.58 112.42 191.7 ;
      RECT 112.94 191.34 113.14 191.46 ;
      RECT 111.5 191.58 111.7 191.7 ;
      RECT 110.78 191.34 110.98 191.46 ;
      RECT 114.02 192.84 114.22 192.96 ;
      RECT 113.3 192.84 113.5 192.96 ;
      RECT 112.58 192.6 112.78 192.72 ;
      RECT 111.14 192.84 111.34 192.96 ;
      RECT 111.86 192.6 112.06 192.72 ;
      RECT 113.66 194.1 113.86 194.22 ;
      RECT 112.22 194.1 112.42 194.22 ;
      RECT 114.38 193.86 114.58 193.98 ;
      RECT 112.94 193.86 113.14 193.98 ;
      RECT 111.5 194.1 111.7 194.22 ;
      RECT 110.78 193.86 110.98 193.98 ;
      RECT 114.02 195.12 114.22 195.24 ;
      RECT 111.86 195.12 112.06 195.24 ;
      RECT 111.14 195.12 111.34 195.24 ;
      RECT 112.58 195.36 112.78 195.48 ;
      RECT 113.3 195.36 113.5 195.48 ;
      RECT 114.38 196.38 114.58 196.5 ;
      RECT 112.94 196.38 113.14 196.5 ;
      RECT 112.22 196.38 112.42 196.5 ;
      RECT 110.78 196.38 110.98 196.5 ;
      RECT 113.66 196.62 113.86 196.74 ;
      RECT 112.58 197.64 112.78 197.76 ;
      RECT 114.02 197.88 114.22 198 ;
      RECT 113.3 197.88 113.5 198 ;
      RECT 111.5 196.62 111.7 196.74 ;
      RECT 111.86 197.64 112.06 197.76 ;
      RECT 111.14 197.88 111.34 198 ;
      RECT 114.38 198.9 114.58 199.02 ;
      RECT 113.66 198.9 113.86 199.02 ;
      RECT 112.94 198.9 113.14 199.02 ;
      RECT 112.22 198.9 112.42 199.02 ;
      RECT 111.5 198.9 111.7 199.02 ;
      RECT 110.78 198.9 110.98 199.02 ;
      RECT 113.3 200.16 113.5 200.28 ;
      RECT 112.58 200.4 112.78 200.52 ;
      RECT 114.02 200.4 114.22 200.52 ;
      RECT 111.86 200.16 112.06 200.28 ;
      RECT 111.14 200.4 111.34 200.52 ;
      RECT 114.38 201.42 114.58 201.54 ;
      RECT 112.22 201.42 112.42 201.54 ;
      RECT 113.66 201.66 113.86 201.78 ;
      RECT 112.94 201.66 113.14 201.78 ;
      RECT 111.5 201.42 111.7 201.54 ;
      RECT 110.78 201.66 110.98 201.78 ;
      RECT 114.02 202.68 114.22 202.8 ;
      RECT 113.3 202.68 113.5 202.8 ;
      RECT 112.58 202.68 112.78 202.8 ;
      RECT 111.14 202.92 111.34 203.04 ;
      RECT 111.86 202.92 112.06 203.04 ;
      RECT 112.94 203.94 113.14 204.06 ;
      RECT 114.38 203.94 114.58 204.06 ;
      RECT 113.66 204.18 113.86 204.3 ;
      RECT 113.3 157.56 113.5 157.68 ;
      RECT 112.58 157.56 112.78 157.68 ;
      RECT 114.02 157.32 114.22 157.44 ;
      RECT 110.78 158.82 110.98 158.94 ;
      RECT 111.5 158.58 111.7 158.7 ;
      RECT 113.66 158.82 113.86 158.94 ;
      RECT 112.22 158.82 112.42 158.94 ;
      RECT 112.94 158.58 113.14 158.7 ;
      RECT 114.38 158.58 114.58 158.7 ;
      RECT 111.86 160.08 112.06 160.2 ;
      RECT 111.14 159.84 111.34 159.96 ;
      RECT 114.02 159.84 114.22 159.96 ;
      RECT 113.3 159.84 113.5 159.96 ;
      RECT 112.58 159.84 112.78 159.96 ;
      RECT 111.86 162.34 112.06 162.46 ;
      RECT 111.14 162.34 111.34 162.46 ;
      RECT 110.78 161.1 110.98 161.22 ;
      RECT 111.5 161.1 111.7 161.22 ;
      RECT 114.02 162.34 114.22 162.46 ;
      RECT 112.58 162.34 112.78 162.46 ;
      RECT 112.22 161.1 112.42 161.22 ;
      RECT 112.94 161.1 113.14 161.22 ;
      RECT 113.66 161.1 113.86 161.22 ;
      RECT 114.38 161.1 114.58 161.22 ;
      RECT 111.5 163.62 111.7 163.74 ;
      RECT 114.38 163.62 114.58 163.74 ;
      RECT 112.94 163.62 113.14 163.74 ;
      RECT 112.22 163.62 112.42 163.74 ;
      RECT 113.3 162.6 113.5 162.72 ;
      RECT 111.86 165.12 112.06 165.24 ;
      RECT 111.14 164.88 111.34 165 ;
      RECT 110.78 163.86 110.98 163.98 ;
      RECT 114.02 164.88 114.22 165 ;
      RECT 113.3 164.88 113.5 165 ;
      RECT 112.58 164.88 112.78 165 ;
      RECT 113.66 163.86 113.86 163.98 ;
      RECT 110.78 166.38 110.98 166.5 ;
      RECT 111.5 166.14 111.7 166.26 ;
      RECT 112.22 166.38 112.42 166.5 ;
      RECT 112.94 166.14 113.14 166.26 ;
      RECT 113.66 166.14 113.86 166.26 ;
      RECT 114.38 166.14 114.58 166.26 ;
      RECT 111.86 167.64 112.06 167.76 ;
      RECT 111.14 167.4 111.34 167.52 ;
      RECT 113.3 167.64 113.5 167.76 ;
      RECT 114.02 167.4 114.22 167.52 ;
      RECT 112.58 167.4 112.78 167.52 ;
      RECT 110.78 168.9 110.98 169.02 ;
      RECT 111.5 168.66 111.7 168.78 ;
      RECT 113.66 168.9 113.86 169.02 ;
      RECT 112.94 168.9 113.14 169.02 ;
      RECT 112.22 168.66 112.42 168.78 ;
      RECT 114.38 168.66 114.58 168.78 ;
      RECT 114.02 169.92 114.22 170.04 ;
      RECT 113.3 169.92 113.5 170.04 ;
      RECT 112.58 169.92 112.78 170.04 ;
      RECT 111.86 170.16 112.06 170.28 ;
      RECT 111.14 170.16 111.34 170.28 ;
      RECT 112.94 171.42 113.14 171.54 ;
      RECT 114.38 171.18 114.58 171.3 ;
      RECT 113.66 171.18 113.86 171.3 ;
      RECT 112.22 171.18 112.42 171.3 ;
      RECT 110.78 171.42 110.98 171.54 ;
      RECT 111.5 171.18 111.7 171.3 ;
      RECT 113.3 172.68 113.5 172.8 ;
      RECT 112.58 172.44 112.78 172.56 ;
      RECT 114.02 172.44 114.22 172.56 ;
      RECT 111.86 172.68 112.06 172.8 ;
      RECT 111.14 172.44 111.34 172.56 ;
      RECT 112.94 173.94 113.14 174.06 ;
      RECT 112.22 173.94 112.42 174.06 ;
      RECT 114.38 173.7 114.58 173.82 ;
      RECT 113.66 173.7 113.86 173.82 ;
      RECT 110.78 173.94 110.98 174.06 ;
      RECT 111.5 173.7 111.7 173.82 ;
      RECT 113.3 175.2 113.5 175.32 ;
      RECT 112.58 174.96 112.78 175.08 ;
      RECT 114.02 174.96 114.22 175.08 ;
      RECT 111.86 175.2 112.06 175.32 ;
      RECT 111.14 175.2 111.34 175.32 ;
      RECT 113.66 176.46 113.86 176.58 ;
      RECT 112.22 176.46 112.42 176.58 ;
      RECT 114.38 176.22 114.58 176.34 ;
      RECT 112.94 176.22 113.14 176.34 ;
      RECT 111.5 176.22 111.7 176.34 ;
      RECT 110.78 176.22 110.98 176.34 ;
      RECT 112.94 178.74 113.14 178.86 ;
      RECT 114.38 178.74 114.58 178.86 ;
      RECT 113.3 177.72 113.5 177.84 ;
      RECT 114.02 177.48 114.22 177.6 ;
      RECT 112.58 177.48 112.78 177.6 ;
      RECT 110.78 178.74 110.98 178.86 ;
      RECT 111.5 178.74 111.7 178.86 ;
      RECT 111.86 177.72 112.06 177.84 ;
      RECT 111.14 177.48 111.34 177.6 ;
      RECT 114.02 180 114.22 180.12 ;
      RECT 113.3 180 113.5 180.12 ;
      RECT 112.58 180 112.78 180.12 ;
      RECT 112.22 178.98 112.42 179.1 ;
      RECT 113.66 178.98 113.86 179.1 ;
      RECT 111.14 180 111.34 180.12 ;
      RECT 112.94 181.5 113.14 181.62 ;
      RECT 113.3 135.598 113.5 135.718 ;
      RECT 114.02 135.358 114.22 135.478 ;
      RECT 112.58 135.358 112.78 135.478 ;
      RECT 111.86 135.598 112.06 135.718 ;
      RECT 111.14 135.358 111.34 135.478 ;
      RECT 113.3 137.4 113.5 137.52 ;
      RECT 112.58 137.16 112.78 137.28 ;
      RECT 114.02 137.16 114.22 137.28 ;
      RECT 112.22 136.858 112.42 136.978 ;
      RECT 112.94 136.858 113.14 136.978 ;
      RECT 113.66 136.618 113.86 136.738 ;
      RECT 114.38 136.618 114.58 136.738 ;
      RECT 111.86 137.4 112.06 137.52 ;
      RECT 113.66 139.138 113.86 139.258 ;
      RECT 112.22 139.138 112.42 139.258 ;
      RECT 113.66 138.66 113.86 138.78 ;
      RECT 112.22 138.66 112.42 138.78 ;
      RECT 114.38 138.42 114.58 138.54 ;
      RECT 112.94 138.42 113.14 138.54 ;
      RECT 114.02 138.118 114.22 138.238 ;
      RECT 113.3 137.878 113.5 137.998 ;
      RECT 112.58 137.878 112.78 137.998 ;
      RECT 111.86 138.118 112.06 138.238 ;
      RECT 114.02 140.398 114.22 140.518 ;
      RECT 112.58 140.398 112.78 140.518 ;
      RECT 113.3 139.92 113.5 140.04 ;
      RECT 114.02 139.68 114.22 139.8 ;
      RECT 112.58 139.68 112.78 139.8 ;
      RECT 114.38 139.378 114.58 139.498 ;
      RECT 112.94 139.378 113.14 139.498 ;
      RECT 111.86 139.92 112.06 140.04 ;
      RECT 113.66 141.18 113.86 141.3 ;
      RECT 112.22 141.18 112.42 141.3 ;
      RECT 112.94 140.94 113.14 141.06 ;
      RECT 114.38 140.94 114.58 141.06 ;
      RECT 113.3 140.638 113.5 140.758 ;
      RECT 110.78 141.18 110.98 141.3 ;
      RECT 111.5 140.94 111.7 141.06 ;
      RECT 111.86 140.638 112.06 140.758 ;
      RECT 113.3 142.44 113.5 142.56 ;
      RECT 114.02 142.2 114.22 142.32 ;
      RECT 112.58 142.2 112.78 142.32 ;
      RECT 111.86 142.44 112.06 142.56 ;
      RECT 111.14 142.44 111.34 142.56 ;
      RECT 112.22 143.46 112.42 143.58 ;
      RECT 112.94 143.46 113.14 143.58 ;
      RECT 113.66 143.46 113.86 143.58 ;
      RECT 114.38 143.46 114.58 143.58 ;
      RECT 110.78 143.46 110.98 143.58 ;
      RECT 111.5 143.46 111.7 143.58 ;
      RECT 110.78 145.98 110.98 146.1 ;
      RECT 111.5 145.98 111.7 146.1 ;
      RECT 111.86 144.96 112.06 145.08 ;
      RECT 111.14 144.72 111.34 144.84 ;
      RECT 112.22 145.98 112.42 146.1 ;
      RECT 112.94 145.98 113.14 146.1 ;
      RECT 113.66 145.98 113.86 146.1 ;
      RECT 114.38 145.98 114.58 146.1 ;
      RECT 113.3 144.96 113.5 145.08 ;
      RECT 112.58 144.72 112.78 144.84 ;
      RECT 114.02 144.72 114.22 144.84 ;
      RECT 110.78 148.5 110.98 148.62 ;
      RECT 111.5 148.5 111.7 148.62 ;
      RECT 112.94 148.74 113.14 148.86 ;
      RECT 112.22 148.5 112.42 148.62 ;
      RECT 113.66 148.5 113.86 148.62 ;
      RECT 114.38 148.5 114.58 148.62 ;
      RECT 111.86 150 112.06 150.12 ;
      RECT 111.14 150 111.34 150.12 ;
      RECT 114.02 150 114.22 150.12 ;
      RECT 113.3 149.76 113.5 149.88 ;
      RECT 112.58 149.76 112.78 149.88 ;
      RECT 110.78 151.26 110.98 151.38 ;
      RECT 111.5 151.02 111.7 151.14 ;
      RECT 112.22 151.26 112.42 151.38 ;
      RECT 114.38 151.02 114.58 151.14 ;
      RECT 113.66 151.02 113.86 151.14 ;
      RECT 112.94 151.02 113.14 151.14 ;
      RECT 111.86 152.52 112.06 152.64 ;
      RECT 111.14 152.28 111.34 152.4 ;
      RECT 114.02 152.52 114.22 152.64 ;
      RECT 113.3 152.52 113.5 152.64 ;
      RECT 112.58 152.28 112.78 152.4 ;
      RECT 110.78 153.78 110.98 153.9 ;
      RECT 111.5 153.54 111.7 153.66 ;
      RECT 113.66 153.78 113.86 153.9 ;
      RECT 112.22 153.78 112.42 153.9 ;
      RECT 112.94 153.54 113.14 153.66 ;
      RECT 114.38 153.54 114.58 153.66 ;
      RECT 111.14 154.8 111.34 154.92 ;
      RECT 111.86 154.8 112.06 154.92 ;
      RECT 114.02 155.04 114.22 155.16 ;
      RECT 113.3 154.8 113.5 154.92 ;
      RECT 112.58 154.8 112.78 154.92 ;
      RECT 111.5 156.3 111.7 156.42 ;
      RECT 110.78 156.3 110.98 156.42 ;
      RECT 113.66 156.3 113.86 156.42 ;
      RECT 112.22 156.3 112.42 156.42 ;
      RECT 112.94 156.06 113.14 156.18 ;
      RECT 114.38 156.06 114.58 156.18 ;
      RECT 111.86 157.32 112.06 157.44 ;
      RECT 111.14 157.32 111.34 157.44 ;
      RECT 106.82 348.339 107.02 348.459 ;
      RECT 107.54 348.339 107.74 348.459 ;
      RECT 108.26 348.339 108.46 348.459 ;
      RECT 108.98 348.339 109.18 348.459 ;
      RECT 109.7 348.339 109.9 348.459 ;
      RECT 110.42 348.339 110.62 348.459 ;
      RECT 113.3 119.76 113.5 119.88 ;
      RECT 114.02 119.76 114.22 119.88 ;
      RECT 112.58 119.52 112.78 119.64 ;
      RECT 113.66 119.218 113.86 119.338 ;
      RECT 112.22 119.218 112.42 119.338 ;
      RECT 114.38 118.978 114.58 119.098 ;
      RECT 112.94 118.978 113.14 119.098 ;
      RECT 111.86 119.52 112.06 119.64 ;
      RECT 112.22 121.02 112.42 121.14 ;
      RECT 113.66 121.02 113.86 121.14 ;
      RECT 112.94 120.78 113.14 120.9 ;
      RECT 114.38 120.78 114.58 120.9 ;
      RECT 113.3 120.478 113.5 120.598 ;
      RECT 112.58 120.238 112.78 120.358 ;
      RECT 114.02 120.238 114.22 120.358 ;
      RECT 111.86 120.478 112.06 120.598 ;
      RECT 112.58 122.758 112.78 122.878 ;
      RECT 114.02 122.758 114.22 122.878 ;
      RECT 112.58 122.28 112.78 122.4 ;
      RECT 114.02 122.28 114.22 122.4 ;
      RECT 113.3 122.04 113.5 122.16 ;
      RECT 112.22 121.738 112.42 121.858 ;
      RECT 113.66 121.738 113.86 121.858 ;
      RECT 112.94 121.498 113.14 121.618 ;
      RECT 114.38 121.498 114.58 121.618 ;
      RECT 111.86 122.28 112.06 122.4 ;
      RECT 112.94 124.018 113.14 124.138 ;
      RECT 114.38 124.018 114.58 124.138 ;
      RECT 112.22 123.54 112.42 123.66 ;
      RECT 113.66 123.54 113.86 123.66 ;
      RECT 112.94 123.3 113.14 123.42 ;
      RECT 114.38 123.3 114.58 123.42 ;
      RECT 113.3 122.998 113.5 123.118 ;
      RECT 111.86 122.998 112.06 123.118 ;
      RECT 113.3 125.518 113.5 125.638 ;
      RECT 112.58 125.278 112.78 125.398 ;
      RECT 114.02 125.278 114.22 125.398 ;
      RECT 112.58 124.8 112.78 124.92 ;
      RECT 114.02 124.8 114.22 124.92 ;
      RECT 113.3 124.56 113.5 124.68 ;
      RECT 112.22 124.258 112.42 124.378 ;
      RECT 113.66 124.258 113.86 124.378 ;
      RECT 111.86 125.518 112.06 125.638 ;
      RECT 111.86 124.8 112.06 124.92 ;
      RECT 112.22 126.06 112.42 126.18 ;
      RECT 113.66 126.06 113.86 126.18 ;
      RECT 114.38 126.06 114.58 126.18 ;
      RECT 112.94 125.82 113.14 125.94 ;
      RECT 114.02 127.32 114.22 127.44 ;
      RECT 113.3 127.32 113.5 127.44 ;
      RECT 112.58 127.08 112.78 127.2 ;
      RECT 111.86 127.32 112.06 127.44 ;
      RECT 111.14 127.08 111.34 127.2 ;
      RECT 114.02 129.6 114.22 129.72 ;
      RECT 112.58 129.6 112.78 129.72 ;
      RECT 113.66 128.58 113.86 128.7 ;
      RECT 112.22 128.58 112.42 128.7 ;
      RECT 114.38 128.34 114.58 128.46 ;
      RECT 112.94 128.34 113.14 128.46 ;
      RECT 111.5 128.58 111.7 128.7 ;
      RECT 110.78 128.58 110.98 128.7 ;
      RECT 114.38 130.86 114.58 130.98 ;
      RECT 112.94 130.86 113.14 130.98 ;
      RECT 112.22 130.86 112.42 130.98 ;
      RECT 113.3 129.84 113.5 129.96 ;
      RECT 111.5 130.86 111.7 130.98 ;
      RECT 111.14 129.84 111.34 129.96 ;
      RECT 111.86 129.84 112.06 129.96 ;
      RECT 113.3 132.36 113.5 132.48 ;
      RECT 114.02 132.12 114.22 132.24 ;
      RECT 112.58 132.12 112.78 132.24 ;
      RECT 113.66 131.1 113.86 131.22 ;
      RECT 111.86 132.36 112.06 132.48 ;
      RECT 111.14 132.36 111.34 132.48 ;
      RECT 110.78 131.1 110.98 131.22 ;
      RECT 113.66 133.62 113.86 133.74 ;
      RECT 112.94 133.62 113.14 133.74 ;
      RECT 112.22 133.38 112.42 133.5 ;
      RECT 114.38 133.38 114.58 133.5 ;
      RECT 110.78 133.38 110.98 133.5 ;
      RECT 111.5 133.38 111.7 133.5 ;
      RECT 113.3 134.88 113.5 135 ;
      RECT 114.02 134.64 114.22 134.76 ;
      RECT 112.58 134.64 112.78 134.76 ;
      RECT 113.66 134.338 113.86 134.458 ;
      RECT 112.22 134.338 112.42 134.458 ;
      RECT 114.38 134.098 114.58 134.218 ;
      RECT 112.94 134.098 113.14 134.218 ;
      RECT 111.86 134.88 112.06 135 ;
      RECT 111.14 134.64 111.34 134.76 ;
      RECT 110.78 134.338 110.98 134.458 ;
      RECT 111.5 134.098 111.7 134.218 ;
      RECT 112.22 136.14 112.42 136.26 ;
      RECT 113.66 136.14 113.86 136.26 ;
      RECT 114.38 136.14 114.58 136.26 ;
      RECT 112.94 135.9 113.14 136.02 ;
      RECT 109.7 260.25 109.9 260.37 ;
      RECT 108.98 260.25 109.18 260.37 ;
      RECT 110.42 260.01 110.62 260.13 ;
      RECT 107.54 260.01 107.74 260.13 ;
      RECT 110.06 259.62 110.26 259.74 ;
      RECT 108.62 259.62 108.82 259.74 ;
      RECT 107.18 259.62 107.38 259.74 ;
      RECT 109.34 259.38 109.54 259.5 ;
      RECT 107.9 259.38 108.1 259.5 ;
      RECT 110.06 261.9 110.26 262.02 ;
      RECT 108.62 261.9 108.82 262.02 ;
      RECT 107.18 261.9 107.38 262.02 ;
      RECT 109.7 261.51 109.9 261.63 ;
      RECT 107.54 261.51 107.74 261.63 ;
      RECT 106.82 261.51 107.02 261.63 ;
      RECT 110.42 261.27 110.62 261.39 ;
      RECT 108.98 261.27 109.18 261.39 ;
      RECT 108.26 261.27 108.46 261.39 ;
      RECT 109.7 262.77 109.9 262.89 ;
      RECT 108.26 262.77 108.46 262.89 ;
      RECT 107.54 262.77 107.74 262.89 ;
      RECT 106.82 262.77 107.02 262.89 ;
      RECT 110.42 262.53 110.62 262.65 ;
      RECT 108.98 262.53 109.18 262.65 ;
      RECT 109.34 262.14 109.54 262.26 ;
      RECT 107.9 262.14 108.1 262.26 ;
      RECT 110.06 264.66 110.26 264.78 ;
      RECT 107.9 264.66 108.1 264.78 ;
      RECT 107.18 264.66 107.38 264.78 ;
      RECT 109.34 264.42 109.54 264.54 ;
      RECT 108.62 264.42 108.82 264.54 ;
      RECT 110.42 264.03 110.62 264.15 ;
      RECT 109.7 264.03 109.9 264.15 ;
      RECT 108.98 264.03 109.18 264.15 ;
      RECT 107.54 264.03 107.74 264.15 ;
      RECT 108.26 263.79 108.46 263.91 ;
      RECT 106.82 263.79 107.02 263.91 ;
      RECT 109.34 267.18 109.54 267.3 ;
      RECT 110.06 266.94 110.26 267.06 ;
      RECT 108.62 266.94 108.82 267.06 ;
      RECT 107.9 266.94 108.1 267.06 ;
      RECT 107.18 266.94 107.38 267.06 ;
      RECT 110.42 266.2885 110.62 266.4085 ;
      RECT 109.7 266.2885 109.9 266.4085 ;
      RECT 108.98 266.2885 109.18 266.4085 ;
      RECT 108.26 266.2885 108.46 266.4085 ;
      RECT 107.54 266.2885 107.74 266.4085 ;
      RECT 106.82 266.2885 107.02 266.4085 ;
      RECT 110.42 267.81 110.62 267.93 ;
      RECT 109.7 267.81 109.9 267.93 ;
      RECT 108.98 267.81 109.18 267.93 ;
      RECT 108.26 267.81 108.46 267.93 ;
      RECT 107.54 267.81 107.74 267.93 ;
      RECT 106.82 267.81 107.02 267.93 ;
      RECT 108.98 270.09 109.18 270.21 ;
      RECT 108.26 270.09 108.46 270.21 ;
      RECT 106.82 270.09 107.02 270.21 ;
      RECT 109.34 269.7 109.54 269.82 ;
      RECT 107.18 269.7 107.38 269.82 ;
      RECT 110.06 269.46 110.26 269.58 ;
      RECT 108.62 269.46 108.82 269.58 ;
      RECT 107.9 269.46 108.1 269.58 ;
      RECT 110.42 271.59 110.62 271.71 ;
      RECT 108.98 271.59 109.18 271.71 ;
      RECT 109.7 271.35 109.9 271.47 ;
      RECT 108.26 271.35 108.46 271.47 ;
      RECT 107.54 271.35 107.74 271.47 ;
      RECT 106.82 271.35 107.02 271.47 ;
      RECT 110.42 270.33 110.62 270.45 ;
      RECT 109.7 270.33 109.9 270.45 ;
      RECT 107.54 270.33 107.74 270.45 ;
      RECT 107.18 272.22 107.38 272.34 ;
      RECT 108.62 272.22 108.82 272.34 ;
      RECT 110.06 271.98 110.26 272.1 ;
      RECT 109.34 271.98 109.54 272.1 ;
      RECT 107.9 271.98 108.1 272.1 ;
      RECT 109.34 274.74 109.54 274.86 ;
      RECT 108.62 274.74 108.82 274.86 ;
      RECT 107.9 274.74 108.1 274.86 ;
      RECT 110.06 274.5 110.26 274.62 ;
      RECT 107.18 274.5 107.38 274.62 ;
      RECT 109.34 277.02 109.54 277.14 ;
      RECT 108.62 277.02 108.82 277.14 ;
      RECT 110.06 277.26 110.26 277.38 ;
      RECT 107.9 277.26 108.1 277.38 ;
      RECT 107.18 277.26 107.38 277.38 ;
      RECT 107.18 308.496 107.38 308.616 ;
      RECT 107.9 308.496 108.1 308.616 ;
      RECT 108.62 308.496 108.82 308.616 ;
      RECT 109.34 308.496 109.54 308.616 ;
      RECT 110.06 308.496 110.26 308.616 ;
      RECT 108.26 323.3835 108.46 323.5035 ;
      RECT 107.54 323.3835 107.74 323.5035 ;
      RECT 106.82 323.3835 107.02 323.5035 ;
      RECT 108.98 323.3835 109.18 323.5035 ;
      RECT 109.7 323.3835 109.9 323.5035 ;
      RECT 110.42 323.3835 110.62 323.5035 ;
      RECT 107.18 325.9425 107.38 326.0625 ;
      RECT 107.9 325.9425 108.1 326.0625 ;
      RECT 109.34 325.9425 109.54 326.0625 ;
      RECT 110.06 325.9425 110.26 326.0625 ;
      RECT 108.62 325.9425 108.82 326.0625 ;
      RECT 108.26 213 108.46 213.12 ;
      RECT 108.98 213 109.18 213.12 ;
      RECT 107.18 214.02 107.38 214.14 ;
      RECT 108.62 214.02 108.82 214.14 ;
      RECT 110.06 214.02 110.26 214.14 ;
      RECT 107.9 214.26 108.1 214.38 ;
      RECT 109.34 214.26 109.54 214.38 ;
      RECT 108.98 215.28 109.18 215.4 ;
      RECT 107.54 215.28 107.74 215.4 ;
      RECT 109.7 215.28 109.9 215.4 ;
      RECT 110.42 215.52 110.62 215.64 ;
      RECT 108.26 215.52 108.46 215.64 ;
      RECT 106.82 215.52 107.02 215.64 ;
      RECT 107.9 216.54 108.1 216.66 ;
      RECT 108.62 216.54 108.82 216.66 ;
      RECT 110.06 216.54 110.26 216.66 ;
      RECT 107.18 216.78 107.38 216.9 ;
      RECT 109.34 216.78 109.54 216.9 ;
      RECT 110.06 219.3 110.26 219.42 ;
      RECT 108.62 219.3 108.82 219.42 ;
      RECT 107.18 219.06 107.38 219.18 ;
      RECT 109.34 219.06 109.54 219.18 ;
      RECT 107.9 219.06 108.1 219.18 ;
      RECT 109.34 223.798 109.54 223.918 ;
      RECT 107.18 223.558 107.38 223.678 ;
      RECT 107.9 223.558 108.1 223.678 ;
      RECT 108.62 223.558 108.82 223.678 ;
      RECT 110.06 223.558 110.26 223.678 ;
      RECT 106.82 223.08 107.02 223.2 ;
      RECT 108.98 223.08 109.18 223.2 ;
      RECT 107.54 222.84 107.74 222.96 ;
      RECT 108.26 222.84 108.46 222.96 ;
      RECT 109.7 222.84 109.9 222.96 ;
      RECT 110.42 222.84 110.62 222.96 ;
      RECT 107.9 229.14 108.1 229.26 ;
      RECT 108.62 229.14 108.82 229.26 ;
      RECT 107.18 229.38 107.38 229.5 ;
      RECT 109.34 229.38 109.54 229.5 ;
      RECT 110.06 229.38 110.26 229.5 ;
      RECT 110.06 231.9 110.26 232.02 ;
      RECT 108.62 231.9 108.82 232.02 ;
      RECT 109.34 231.66 109.54 231.78 ;
      RECT 107.9 231.66 108.1 231.78 ;
      RECT 107.18 231.66 107.38 231.78 ;
      RECT 110.06 234.42 110.26 234.54 ;
      RECT 108.62 234.42 108.82 234.54 ;
      RECT 107.18 234.18 107.38 234.3 ;
      RECT 107.9 234.18 108.1 234.3 ;
      RECT 109.34 234.18 109.54 234.3 ;
      RECT 107.9 236.94 108.1 237.06 ;
      RECT 110.06 236.94 110.26 237.06 ;
      RECT 107.18 236.7 107.38 236.82 ;
      RECT 108.62 236.7 108.82 236.82 ;
      RECT 109.34 236.7 109.54 236.82 ;
      RECT 109.34 239.46 109.54 239.58 ;
      RECT 107.9 239.46 108.1 239.58 ;
      RECT 107.18 239.46 107.38 239.58 ;
      RECT 110.06 239.22 110.26 239.34 ;
      RECT 108.62 239.22 108.82 239.34 ;
      RECT 108.62 241.98 108.82 242.1 ;
      RECT 107.18 241.74 107.38 241.86 ;
      RECT 107.9 241.74 108.1 241.86 ;
      RECT 109.34 241.74 109.54 241.86 ;
      RECT 110.06 241.74 110.26 241.86 ;
      RECT 110.06 244.26 110.26 244.38 ;
      RECT 108.62 244.26 108.82 244.38 ;
      RECT 107.18 244.26 107.38 244.38 ;
      RECT 107.9 244.5 108.1 244.62 ;
      RECT 109.34 244.5 109.54 244.62 ;
      RECT 109.34 247.02 109.54 247.14 ;
      RECT 107.9 247.02 108.1 247.14 ;
      RECT 110.06 246.78 110.26 246.9 ;
      RECT 108.62 246.78 108.82 246.9 ;
      RECT 107.18 246.78 107.38 246.9 ;
      RECT 109.34 249.54 109.54 249.66 ;
      RECT 107.9 249.54 108.1 249.66 ;
      RECT 110.06 249.3 110.26 249.42 ;
      RECT 108.62 249.3 108.82 249.42 ;
      RECT 107.18 249.3 107.38 249.42 ;
      RECT 109.34 252.06 109.54 252.18 ;
      RECT 107.9 252.06 108.1 252.18 ;
      RECT 110.06 251.82 110.26 251.94 ;
      RECT 108.62 251.82 108.82 251.94 ;
      RECT 107.18 251.82 107.38 251.94 ;
      RECT 108.62 254.58 108.82 254.7 ;
      RECT 107.18 254.58 107.38 254.7 ;
      RECT 110.06 254.34 110.26 254.46 ;
      RECT 109.34 254.34 109.54 254.46 ;
      RECT 107.9 254.34 108.1 254.46 ;
      RECT 110.06 257.1 110.26 257.22 ;
      RECT 108.62 257.1 108.82 257.22 ;
      RECT 107.18 257.1 107.38 257.22 ;
      RECT 109.34 256.86 109.54 256.98 ;
      RECT 107.9 256.86 108.1 256.98 ;
      RECT 109.7 258.99 109.9 259.11 ;
      RECT 108.98 258.99 109.18 259.11 ;
      RECT 107.54 258.99 107.74 259.11 ;
      RECT 110.42 258.75 110.62 258.87 ;
      RECT 108.26 258.75 108.46 258.87 ;
      RECT 106.82 258.75 107.02 258.87 ;
      RECT 108.26 260.25 108.46 260.37 ;
      RECT 106.82 260.25 107.02 260.37 ;
      RECT 108.26 190.32 108.46 190.44 ;
      RECT 106.82 190.08 107.02 190.2 ;
      RECT 107.54 190.08 107.74 190.2 ;
      RECT 108.98 190.08 109.18 190.2 ;
      RECT 110.42 190.08 110.62 190.2 ;
      RECT 108.62 191.58 108.82 191.7 ;
      RECT 107.9 191.58 108.1 191.7 ;
      RECT 107.18 191.58 107.38 191.7 ;
      RECT 110.06 191.34 110.26 191.46 ;
      RECT 109.34 191.34 109.54 191.46 ;
      RECT 110.42 192.84 110.62 192.96 ;
      RECT 108.98 192.84 109.18 192.96 ;
      RECT 106.82 192.84 107.02 192.96 ;
      RECT 107.54 192.6 107.74 192.72 ;
      RECT 108.26 192.6 108.46 192.72 ;
      RECT 109.7 192.6 109.9 192.72 ;
      RECT 110.06 194.1 110.26 194.22 ;
      RECT 108.62 194.1 108.82 194.22 ;
      RECT 109.34 193.86 109.54 193.98 ;
      RECT 107.9 193.86 108.1 193.98 ;
      RECT 107.18 193.86 107.38 193.98 ;
      RECT 110.42 195.12 110.62 195.24 ;
      RECT 109.7 195.12 109.9 195.24 ;
      RECT 108.98 195.12 109.18 195.24 ;
      RECT 106.82 195.12 107.02 195.24 ;
      RECT 107.54 195.36 107.74 195.48 ;
      RECT 108.26 195.36 108.46 195.48 ;
      RECT 108.62 196.38 108.82 196.5 ;
      RECT 107.9 196.38 108.1 196.5 ;
      RECT 107.18 196.62 107.38 196.74 ;
      RECT 109.34 196.62 109.54 196.74 ;
      RECT 110.06 196.62 110.26 196.74 ;
      RECT 106.82 197.64 107.02 197.76 ;
      RECT 108.98 197.64 109.18 197.76 ;
      RECT 110.42 197.64 110.62 197.76 ;
      RECT 109.7 197.88 109.9 198 ;
      RECT 108.26 197.88 108.46 198 ;
      RECT 107.54 197.88 107.74 198 ;
      RECT 107.9 198.9 108.1 199.02 ;
      RECT 110.06 198.9 110.26 199.02 ;
      RECT 108.62 198.9 108.82 199.02 ;
      RECT 107.18 199.14 107.38 199.26 ;
      RECT 109.34 199.14 109.54 199.26 ;
      RECT 106.82 200.16 107.02 200.28 ;
      RECT 107.54 200.16 107.74 200.28 ;
      RECT 108.98 200.16 109.18 200.28 ;
      RECT 108.26 200.4 108.46 200.52 ;
      RECT 109.7 200.4 109.9 200.52 ;
      RECT 110.42 200.4 110.62 200.52 ;
      RECT 109.34 201.42 109.54 201.54 ;
      RECT 108.62 201.42 108.82 201.54 ;
      RECT 107.9 201.42 108.1 201.54 ;
      RECT 110.06 201.66 110.26 201.78 ;
      RECT 107.18 201.66 107.38 201.78 ;
      RECT 108.98 202.68 109.18 202.8 ;
      RECT 108.26 202.68 108.46 202.8 ;
      RECT 106.82 202.68 107.02 202.8 ;
      RECT 107.54 202.92 107.74 203.04 ;
      RECT 109.7 202.92 109.9 203.04 ;
      RECT 110.42 202.92 110.62 203.04 ;
      RECT 107.18 203.94 107.38 204.06 ;
      RECT 109.34 203.94 109.54 204.06 ;
      RECT 110.06 204.18 110.26 204.3 ;
      RECT 108.62 204.18 108.82 204.3 ;
      RECT 107.9 204.18 108.1 204.3 ;
      RECT 106.82 205.2 107.02 205.32 ;
      RECT 108.98 205.2 109.18 205.32 ;
      RECT 109.7 205.2 109.9 205.32 ;
      RECT 110.42 205.44 110.62 205.56 ;
      RECT 108.26 205.44 108.46 205.56 ;
      RECT 107.54 205.44 107.74 205.56 ;
      RECT 108.62 206.46 108.82 206.58 ;
      RECT 110.06 206.7 110.26 206.82 ;
      RECT 109.34 206.7 109.54 206.82 ;
      RECT 107.9 206.7 108.1 206.82 ;
      RECT 107.18 206.7 107.38 206.82 ;
      RECT 110.42 207.72 110.62 207.84 ;
      RECT 108.26 207.72 108.46 207.84 ;
      RECT 109.7 207.96 109.9 208.08 ;
      RECT 108.98 207.96 109.18 208.08 ;
      RECT 107.54 207.96 107.74 208.08 ;
      RECT 106.82 207.96 107.02 208.08 ;
      RECT 110.06 208.98 110.26 209.1 ;
      RECT 109.34 208.98 109.54 209.1 ;
      RECT 108.62 208.98 108.82 209.1 ;
      RECT 107.18 208.98 107.38 209.1 ;
      RECT 107.9 209.22 108.1 209.34 ;
      RECT 109.7 210.48 109.9 210.6 ;
      RECT 108.98 210.48 109.18 210.6 ;
      RECT 108.26 210.48 108.46 210.6 ;
      RECT 107.18 211.5 107.38 211.62 ;
      RECT 110.06 211.5 110.26 211.62 ;
      RECT 110.42 210.24 110.62 210.36 ;
      RECT 107.54 210.24 107.74 210.36 ;
      RECT 106.82 210.24 107.02 210.36 ;
      RECT 107.9 211.74 108.1 211.86 ;
      RECT 108.62 211.74 108.82 211.86 ;
      RECT 109.34 211.74 109.54 211.86 ;
      RECT 110.42 212.76 110.62 212.88 ;
      RECT 109.7 212.76 109.9 212.88 ;
      RECT 107.54 212.76 107.74 212.88 ;
      RECT 106.82 213 107.02 213.12 ;
      RECT 110.06 166.14 110.26 166.26 ;
      RECT 107.18 166.14 107.38 166.26 ;
      RECT 110.42 167.64 110.62 167.76 ;
      RECT 109.7 167.64 109.9 167.76 ;
      RECT 108.26 167.64 108.46 167.76 ;
      RECT 106.82 167.64 107.02 167.76 ;
      RECT 108.98 167.4 109.18 167.52 ;
      RECT 107.54 167.4 107.74 167.52 ;
      RECT 110.06 168.9 110.26 169.02 ;
      RECT 107.9 168.9 108.1 169.02 ;
      RECT 107.18 168.9 107.38 169.02 ;
      RECT 108.62 168.66 108.82 168.78 ;
      RECT 109.34 168.66 109.54 168.78 ;
      RECT 109.7 170.16 109.9 170.28 ;
      RECT 108.98 170.16 109.18 170.28 ;
      RECT 107.54 170.16 107.74 170.28 ;
      RECT 110.42 169.92 110.62 170.04 ;
      RECT 108.26 169.92 108.46 170.04 ;
      RECT 106.82 169.92 107.02 170.04 ;
      RECT 109.34 171.42 109.54 171.54 ;
      RECT 107.9 171.42 108.1 171.54 ;
      RECT 110.06 171.18 110.26 171.3 ;
      RECT 108.62 171.18 108.82 171.3 ;
      RECT 107.18 171.18 107.38 171.3 ;
      RECT 106.82 172.68 107.02 172.8 ;
      RECT 110.42 172.68 110.62 172.8 ;
      RECT 109.7 172.68 109.9 172.8 ;
      RECT 108.98 172.68 109.18 172.8 ;
      RECT 107.54 172.68 107.74 172.8 ;
      RECT 108.26 172.44 108.46 172.56 ;
      RECT 109.34 173.94 109.54 174.06 ;
      RECT 107.18 173.94 107.38 174.06 ;
      RECT 110.06 173.7 110.26 173.82 ;
      RECT 108.62 173.7 108.82 173.82 ;
      RECT 107.9 173.7 108.1 173.82 ;
      RECT 109.7 175.2 109.9 175.32 ;
      RECT 107.54 175.2 107.74 175.32 ;
      RECT 106.82 175.2 107.02 175.32 ;
      RECT 108.26 174.96 108.46 175.08 ;
      RECT 108.98 174.96 109.18 175.08 ;
      RECT 110.42 174.96 110.62 175.08 ;
      RECT 110.06 176.46 110.26 176.58 ;
      RECT 108.62 176.46 108.82 176.58 ;
      RECT 109.34 176.22 109.54 176.34 ;
      RECT 107.9 176.22 108.1 176.34 ;
      RECT 107.18 176.22 107.38 176.34 ;
      RECT 108.62 178.74 108.82 178.86 ;
      RECT 109.34 178.74 109.54 178.86 ;
      RECT 106.82 177.72 107.02 177.84 ;
      RECT 107.54 177.72 107.74 177.84 ;
      RECT 109.7 177.72 109.9 177.84 ;
      RECT 108.26 177.72 108.46 177.84 ;
      RECT 110.42 177.48 110.62 177.6 ;
      RECT 108.98 177.48 109.18 177.6 ;
      RECT 109.7 180 109.9 180.12 ;
      RECT 107.54 180 107.74 180.12 ;
      RECT 106.82 180 107.02 180.12 ;
      RECT 110.06 178.98 110.26 179.1 ;
      RECT 107.9 178.98 108.1 179.1 ;
      RECT 107.18 178.98 107.38 179.1 ;
      RECT 109.34 181.5 109.54 181.62 ;
      RECT 107.18 181.26 107.38 181.38 ;
      RECT 107.9 181.26 108.1 181.38 ;
      RECT 108.62 181.26 108.82 181.38 ;
      RECT 110.06 181.26 110.26 181.38 ;
      RECT 110.42 180.24 110.62 180.36 ;
      RECT 108.98 180.24 109.18 180.36 ;
      RECT 108.26 180.24 108.46 180.36 ;
      RECT 108.26 182.76 108.46 182.88 ;
      RECT 106.82 182.76 107.02 182.88 ;
      RECT 110.42 182.52 110.62 182.64 ;
      RECT 109.7 182.52 109.9 182.64 ;
      RECT 108.98 182.52 109.18 182.64 ;
      RECT 107.54 182.52 107.74 182.64 ;
      RECT 109.34 184.02 109.54 184.14 ;
      RECT 108.62 184.02 108.82 184.14 ;
      RECT 110.06 183.78 110.26 183.9 ;
      RECT 107.9 183.78 108.1 183.9 ;
      RECT 107.18 183.78 107.38 183.9 ;
      RECT 106.82 185.28 107.02 185.4 ;
      RECT 108.26 185.28 108.46 185.4 ;
      RECT 110.42 185.28 110.62 185.4 ;
      RECT 109.7 185.04 109.9 185.16 ;
      RECT 108.98 185.04 109.18 185.16 ;
      RECT 107.54 185.04 107.74 185.16 ;
      RECT 108.62 186.54 108.82 186.66 ;
      RECT 109.34 186.54 109.54 186.66 ;
      RECT 110.06 186.3 110.26 186.42 ;
      RECT 107.9 186.3 108.1 186.42 ;
      RECT 107.18 186.3 107.38 186.42 ;
      RECT 109.7 187.8 109.9 187.92 ;
      RECT 108.26 187.8 108.46 187.92 ;
      RECT 106.82 187.8 107.02 187.92 ;
      RECT 107.54 187.56 107.74 187.68 ;
      RECT 110.42 187.56 110.62 187.68 ;
      RECT 108.98 187.56 109.18 187.68 ;
      RECT 107.9 189.06 108.1 189.18 ;
      RECT 110.06 188.82 110.26 188.94 ;
      RECT 109.34 188.82 109.54 188.94 ;
      RECT 108.62 188.82 108.82 188.94 ;
      RECT 107.18 188.82 107.38 188.94 ;
      RECT 109.7 190.32 109.9 190.44 ;
      RECT 108.98 142.44 109.18 142.56 ;
      RECT 108.26 142.44 108.46 142.56 ;
      RECT 110.42 142.2 110.62 142.32 ;
      RECT 109.7 142.2 109.9 142.32 ;
      RECT 107.54 142.2 107.74 142.32 ;
      RECT 106.82 142.2 107.02 142.32 ;
      RECT 107.18 143.46 107.38 143.58 ;
      RECT 107.9 143.46 108.1 143.58 ;
      RECT 108.62 143.46 108.82 143.58 ;
      RECT 109.34 143.46 109.54 143.58 ;
      RECT 110.06 143.46 110.26 143.58 ;
      RECT 107.18 145.98 107.38 146.1 ;
      RECT 107.9 145.98 108.1 146.1 ;
      RECT 108.62 145.98 108.82 146.1 ;
      RECT 109.34 145.98 109.54 146.1 ;
      RECT 110.06 145.98 110.26 146.1 ;
      RECT 107.54 144.96 107.74 145.08 ;
      RECT 108.98 144.96 109.18 145.08 ;
      RECT 110.42 144.96 110.62 145.08 ;
      RECT 106.82 144.72 107.02 144.84 ;
      RECT 108.26 144.72 108.46 144.84 ;
      RECT 109.7 144.72 109.9 144.84 ;
      RECT 110.06 148.74 110.26 148.86 ;
      RECT 108.62 148.74 108.82 148.86 ;
      RECT 107.9 148.74 108.1 148.86 ;
      RECT 107.18 148.5 107.38 148.62 ;
      RECT 109.34 148.5 109.54 148.62 ;
      RECT 109.7 150 109.9 150.12 ;
      RECT 110.42 149.76 110.62 149.88 ;
      RECT 108.98 149.76 109.18 149.88 ;
      RECT 108.26 149.76 108.46 149.88 ;
      RECT 107.54 149.76 107.74 149.88 ;
      RECT 106.82 149.76 107.02 149.88 ;
      RECT 110.06 151.26 110.26 151.38 ;
      RECT 109.34 151.26 109.54 151.38 ;
      RECT 107.9 151.26 108.1 151.38 ;
      RECT 107.18 151.26 107.38 151.38 ;
      RECT 108.62 151.02 108.82 151.14 ;
      RECT 110.42 152.52 110.62 152.64 ;
      RECT 108.98 152.52 109.18 152.64 ;
      RECT 106.82 152.52 107.02 152.64 ;
      RECT 109.7 152.28 109.9 152.4 ;
      RECT 108.26 152.28 108.46 152.4 ;
      RECT 107.54 152.28 107.74 152.4 ;
      RECT 109.34 153.78 109.54 153.9 ;
      RECT 107.18 153.54 107.38 153.66 ;
      RECT 107.9 153.54 108.1 153.66 ;
      RECT 108.62 153.54 108.82 153.66 ;
      RECT 110.06 153.54 110.26 153.66 ;
      RECT 109.7 155.04 109.9 155.16 ;
      RECT 108.98 155.04 109.18 155.16 ;
      RECT 107.54 155.04 107.74 155.16 ;
      RECT 106.82 154.8 107.02 154.92 ;
      RECT 108.26 154.8 108.46 154.92 ;
      RECT 110.42 154.8 110.62 154.92 ;
      RECT 108.62 156.3 108.82 156.42 ;
      RECT 107.9 156.3 108.1 156.42 ;
      RECT 110.06 156.06 110.26 156.18 ;
      RECT 109.34 156.06 109.54 156.18 ;
      RECT 107.18 156.06 107.38 156.18 ;
      RECT 110.42 157.56 110.62 157.68 ;
      RECT 107.54 157.56 107.74 157.68 ;
      RECT 109.7 157.32 109.9 157.44 ;
      RECT 108.98 157.32 109.18 157.44 ;
      RECT 108.26 157.32 108.46 157.44 ;
      RECT 106.82 157.32 107.02 157.44 ;
      RECT 109.34 158.82 109.54 158.94 ;
      RECT 107.18 158.82 107.38 158.94 ;
      RECT 107.9 158.58 108.1 158.7 ;
      RECT 108.62 158.58 108.82 158.7 ;
      RECT 110.06 158.58 110.26 158.7 ;
      RECT 110.42 160.08 110.62 160.2 ;
      RECT 108.26 160.08 108.46 160.2 ;
      RECT 109.7 159.84 109.9 159.96 ;
      RECT 108.98 159.84 109.18 159.96 ;
      RECT 107.54 159.84 107.74 159.96 ;
      RECT 106.82 159.84 107.02 159.96 ;
      RECT 110.42 162.34 110.62 162.46 ;
      RECT 108.98 162.34 109.18 162.46 ;
      RECT 108.26 162.34 108.46 162.46 ;
      RECT 107.54 162.34 107.74 162.46 ;
      RECT 107.18 161.1 107.38 161.22 ;
      RECT 107.9 161.1 108.1 161.22 ;
      RECT 108.62 161.1 108.82 161.22 ;
      RECT 109.34 161.1 109.54 161.22 ;
      RECT 110.06 161.1 110.26 161.22 ;
      RECT 110.06 163.62 110.26 163.74 ;
      RECT 108.62 163.62 108.82 163.74 ;
      RECT 107.18 163.62 107.38 163.74 ;
      RECT 106.82 162.6 107.02 162.72 ;
      RECT 109.7 162.6 109.9 162.72 ;
      RECT 109.7 165.12 109.9 165.24 ;
      RECT 108.26 165.12 108.46 165.24 ;
      RECT 106.82 165.12 107.02 165.24 ;
      RECT 110.42 164.88 110.62 165 ;
      RECT 108.98 164.88 109.18 165 ;
      RECT 107.54 164.88 107.74 165 ;
      RECT 109.34 163.86 109.54 163.98 ;
      RECT 107.9 163.86 108.1 163.98 ;
      RECT 107.9 166.38 108.1 166.5 ;
      RECT 108.62 166.38 108.82 166.5 ;
      RECT 109.34 166.38 109.54 166.5 ;
      RECT 103.22 271.35 103.42 271.47 ;
      RECT 103.94 271.35 104.14 271.47 ;
      RECT 104.66 270.33 104.86 270.45 ;
      RECT 103.94 270.33 104.14 270.45 ;
      RECT 103.22 270.33 103.42 270.45 ;
      RECT 106.46 272.22 106.66 272.34 ;
      RECT 105.02 272.22 105.22 272.34 ;
      RECT 104.3 272.22 104.5 272.34 ;
      RECT 103.58 272.22 103.78 272.34 ;
      RECT 105.74 271.98 105.94 272.1 ;
      RECT 102.86 271.98 103.06 272.1 ;
      RECT 106.46 274.74 106.66 274.86 ;
      RECT 104.3 274.74 104.5 274.86 ;
      RECT 102.86 274.74 103.06 274.86 ;
      RECT 105.74 274.5 105.94 274.62 ;
      RECT 105.02 274.5 105.22 274.62 ;
      RECT 103.58 274.5 103.78 274.62 ;
      RECT 106.46 277.02 106.66 277.14 ;
      RECT 105.74 277.02 105.94 277.14 ;
      RECT 105.02 277.02 105.22 277.14 ;
      RECT 103.58 277.02 103.78 277.14 ;
      RECT 104.3 277.26 104.5 277.38 ;
      RECT 102.86 277.26 103.06 277.38 ;
      RECT 102.86 308.496 103.06 308.616 ;
      RECT 103.58 308.496 103.78 308.616 ;
      RECT 104.3 308.496 104.5 308.616 ;
      RECT 105.02 308.496 105.22 308.616 ;
      RECT 105.74 308.496 105.94 308.616 ;
      RECT 106.46 308.496 106.66 308.616 ;
      RECT 106.1 323.3835 106.3 323.5035 ;
      RECT 105.38 323.3835 105.58 323.5035 ;
      RECT 104.66 323.3835 104.86 323.5035 ;
      RECT 102.5 323.3835 102.7 323.5035 ;
      RECT 103.22 323.3835 103.42 323.5035 ;
      RECT 103.94 323.3835 104.14 323.5035 ;
      RECT 102.86 325.9425 103.06 326.0625 ;
      RECT 103.58 325.9425 103.78 326.0625 ;
      RECT 104.3 325.9425 104.5 326.0625 ;
      RECT 105.02 325.9425 105.22 326.0625 ;
      RECT 105.74 325.9425 105.94 326.0625 ;
      RECT 106.46 325.9425 106.66 326.0625 ;
      RECT 102.5 348.339 102.7 348.459 ;
      RECT 103.22 348.339 103.42 348.459 ;
      RECT 103.94 348.339 104.14 348.459 ;
      RECT 104.66 348.339 104.86 348.459 ;
      RECT 105.38 348.339 105.58 348.459 ;
      RECT 106.1 348.339 106.3 348.459 ;
      RECT 109.7 127.32 109.9 127.44 ;
      RECT 108.26 127.32 108.46 127.44 ;
      RECT 107.54 127.32 107.74 127.44 ;
      RECT 110.42 127.08 110.62 127.2 ;
      RECT 108.98 127.08 109.18 127.2 ;
      RECT 106.82 127.08 107.02 127.2 ;
      RECT 110.42 129.6 110.62 129.72 ;
      RECT 108.98 129.6 109.18 129.72 ;
      RECT 107.54 129.6 107.74 129.72 ;
      RECT 107.9 128.58 108.1 128.7 ;
      RECT 109.34 128.58 109.54 128.7 ;
      RECT 110.06 128.34 110.26 128.46 ;
      RECT 108.62 128.34 108.82 128.46 ;
      RECT 107.18 128.34 107.38 128.46 ;
      RECT 109.34 130.86 109.54 130.98 ;
      RECT 108.62 130.86 108.82 130.98 ;
      RECT 106.82 129.84 107.02 129.96 ;
      RECT 108.26 129.84 108.46 129.96 ;
      RECT 109.7 129.84 109.9 129.96 ;
      RECT 110.42 132.36 110.62 132.48 ;
      RECT 108.26 132.36 108.46 132.48 ;
      RECT 106.82 132.36 107.02 132.48 ;
      RECT 109.7 132.12 109.9 132.24 ;
      RECT 108.98 132.12 109.18 132.24 ;
      RECT 107.54 132.12 107.74 132.24 ;
      RECT 110.06 131.1 110.26 131.22 ;
      RECT 107.18 131.1 107.38 131.22 ;
      RECT 107.9 131.1 108.1 131.22 ;
      RECT 110.06 133.62 110.26 133.74 ;
      RECT 108.62 133.62 108.82 133.74 ;
      RECT 107.18 133.62 107.38 133.74 ;
      RECT 107.9 133.38 108.1 133.5 ;
      RECT 109.34 133.38 109.54 133.5 ;
      RECT 110.42 134.88 110.62 135 ;
      RECT 108.98 134.88 109.18 135 ;
      RECT 108.26 134.88 108.46 135 ;
      RECT 106.82 134.88 107.02 135 ;
      RECT 109.7 134.64 109.9 134.76 ;
      RECT 107.54 134.64 107.74 134.76 ;
      RECT 107.9 134.338 108.1 134.458 ;
      RECT 110.06 134.098 110.26 134.218 ;
      RECT 109.34 134.098 109.54 134.218 ;
      RECT 108.62 134.098 108.82 134.218 ;
      RECT 107.18 134.098 107.38 134.218 ;
      RECT 110.42 135.598 110.62 135.718 ;
      RECT 109.7 135.598 109.9 135.718 ;
      RECT 108.26 135.598 108.46 135.718 ;
      RECT 106.82 135.598 107.02 135.718 ;
      RECT 108.98 135.358 109.18 135.478 ;
      RECT 107.54 135.358 107.74 135.478 ;
      RECT 109.34 141.18 109.54 141.3 ;
      RECT 107.18 141.18 107.38 141.3 ;
      RECT 107.9 140.94 108.1 141.06 ;
      RECT 108.62 140.94 108.82 141.06 ;
      RECT 110.06 140.94 110.26 141.06 ;
      RECT 105.02 249.54 105.22 249.66 ;
      RECT 102.86 249.54 103.06 249.66 ;
      RECT 104.3 249.54 104.5 249.66 ;
      RECT 105.74 249.3 105.94 249.42 ;
      RECT 103.58 249.3 103.78 249.42 ;
      RECT 106.46 252.06 106.66 252.18 ;
      RECT 104.3 252.06 104.5 252.18 ;
      RECT 102.86 252.06 103.06 252.18 ;
      RECT 105.74 251.82 105.94 251.94 ;
      RECT 105.02 251.82 105.22 251.94 ;
      RECT 103.58 251.82 103.78 251.94 ;
      RECT 105.74 254.58 105.94 254.7 ;
      RECT 105.02 254.58 105.22 254.7 ;
      RECT 103.58 254.58 103.78 254.7 ;
      RECT 106.46 254.34 106.66 254.46 ;
      RECT 104.3 254.34 104.5 254.46 ;
      RECT 102.86 254.34 103.06 254.46 ;
      RECT 106.46 257.1 106.66 257.22 ;
      RECT 105.74 257.1 105.94 257.22 ;
      RECT 102.86 257.1 103.06 257.22 ;
      RECT 105.02 256.86 105.22 256.98 ;
      RECT 104.3 256.86 104.5 256.98 ;
      RECT 103.58 256.86 103.78 256.98 ;
      RECT 106.1 258.99 106.3 259.11 ;
      RECT 104.66 258.99 104.86 259.11 ;
      RECT 102.5 258.99 102.7 259.11 ;
      RECT 105.38 258.75 105.58 258.87 ;
      RECT 103.94 258.75 104.14 258.87 ;
      RECT 103.22 258.75 103.42 258.87 ;
      RECT 105.38 260.25 105.58 260.37 ;
      RECT 103.94 260.25 104.14 260.37 ;
      RECT 103.22 260.25 103.42 260.37 ;
      RECT 106.1 260.01 106.3 260.13 ;
      RECT 104.66 260.01 104.86 260.13 ;
      RECT 102.5 260.01 102.7 260.13 ;
      RECT 106.46 259.62 106.66 259.74 ;
      RECT 104.3 259.62 104.5 259.74 ;
      RECT 103.58 259.38 103.78 259.5 ;
      RECT 102.86 259.38 103.06 259.5 ;
      RECT 105.02 259.38 105.22 259.5 ;
      RECT 105.74 259.38 105.94 259.5 ;
      RECT 105.02 261.9 105.22 262.02 ;
      RECT 106.1 261.51 106.3 261.63 ;
      RECT 105.38 261.51 105.58 261.63 ;
      RECT 103.94 261.51 104.14 261.63 ;
      RECT 102.5 261.51 102.7 261.63 ;
      RECT 104.66 261.27 104.86 261.39 ;
      RECT 103.22 261.27 103.42 261.39 ;
      RECT 106.1 262.77 106.3 262.89 ;
      RECT 105.38 262.77 105.58 262.89 ;
      RECT 104.66 262.77 104.86 262.89 ;
      RECT 103.94 262.77 104.14 262.89 ;
      RECT 102.5 262.77 102.7 262.89 ;
      RECT 103.22 262.53 103.42 262.65 ;
      RECT 106.46 262.14 106.66 262.26 ;
      RECT 105.74 262.14 105.94 262.26 ;
      RECT 104.3 262.14 104.5 262.26 ;
      RECT 103.58 262.14 103.78 262.26 ;
      RECT 102.86 262.14 103.06 262.26 ;
      RECT 104.3 264.66 104.5 264.78 ;
      RECT 103.58 264.66 103.78 264.78 ;
      RECT 105.02 264.42 105.22 264.54 ;
      RECT 106.46 264.42 106.66 264.54 ;
      RECT 105.74 264.42 105.94 264.54 ;
      RECT 102.86 264.42 103.06 264.54 ;
      RECT 106.1 264.03 106.3 264.15 ;
      RECT 104.66 264.03 104.86 264.15 ;
      RECT 103.94 264.03 104.14 264.15 ;
      RECT 102.5 264.03 102.7 264.15 ;
      RECT 105.38 263.79 105.58 263.91 ;
      RECT 103.22 263.79 103.42 263.91 ;
      RECT 105.74 267.18 105.94 267.3 ;
      RECT 102.86 267.18 103.06 267.3 ;
      RECT 106.46 266.94 106.66 267.06 ;
      RECT 105.02 266.94 105.22 267.06 ;
      RECT 103.58 266.94 103.78 267.06 ;
      RECT 104.3 266.94 104.5 267.06 ;
      RECT 106.1 266.2885 106.3 266.4085 ;
      RECT 105.38 266.2885 105.58 266.4085 ;
      RECT 104.66 266.2885 104.86 266.4085 ;
      RECT 103.94 266.2885 104.14 266.4085 ;
      RECT 103.22 266.2885 103.42 266.4085 ;
      RECT 102.5 266.2885 102.7 266.4085 ;
      RECT 106.1 267.81 106.3 267.93 ;
      RECT 105.38 267.81 105.58 267.93 ;
      RECT 104.66 267.81 104.86 267.93 ;
      RECT 103.94 267.81 104.14 267.93 ;
      RECT 103.22 267.81 103.42 267.93 ;
      RECT 102.5 267.81 102.7 267.93 ;
      RECT 106.1 270.09 106.3 270.21 ;
      RECT 105.38 270.09 105.58 270.21 ;
      RECT 102.5 270.09 102.7 270.21 ;
      RECT 105.74 269.7 105.94 269.82 ;
      RECT 104.3 269.7 104.5 269.82 ;
      RECT 102.86 269.7 103.06 269.82 ;
      RECT 106.46 269.46 106.66 269.58 ;
      RECT 105.02 269.46 105.22 269.58 ;
      RECT 103.58 269.46 103.78 269.58 ;
      RECT 106.1 271.59 106.3 271.71 ;
      RECT 105.38 271.59 105.58 271.71 ;
      RECT 104.66 271.59 104.86 271.71 ;
      RECT 102.5 271.59 102.7 271.71 ;
      RECT 105.02 211.5 105.22 211.62 ;
      RECT 103.58 211.5 103.78 211.62 ;
      RECT 103.94 210.48 104.14 210.6 ;
      RECT 104.66 210.48 104.86 210.6 ;
      RECT 105.38 210.48 105.58 210.6 ;
      RECT 102.5 210.24 102.7 210.36 ;
      RECT 103.22 210.24 103.42 210.36 ;
      RECT 106.1 210.24 106.3 210.36 ;
      RECT 103.22 212.76 103.42 212.88 ;
      RECT 104.66 212.76 104.86 212.88 ;
      RECT 106.46 211.74 106.66 211.86 ;
      RECT 104.3 211.74 104.5 211.86 ;
      RECT 102.86 211.74 103.06 211.86 ;
      RECT 105.74 214.26 105.94 214.38 ;
      RECT 104.3 214.26 104.5 214.38 ;
      RECT 103.58 214.26 103.78 214.38 ;
      RECT 106.46 214.02 106.66 214.14 ;
      RECT 105.02 214.02 105.22 214.14 ;
      RECT 102.86 214.02 103.06 214.14 ;
      RECT 102.5 213 102.7 213.12 ;
      RECT 103.94 213 104.14 213.12 ;
      RECT 106.1 213 106.3 213.12 ;
      RECT 105.38 213 105.58 213.12 ;
      RECT 103.94 215.52 104.14 215.64 ;
      RECT 104.66 215.52 104.86 215.64 ;
      RECT 102.5 215.52 102.7 215.64 ;
      RECT 103.22 215.28 103.42 215.4 ;
      RECT 105.38 215.28 105.58 215.4 ;
      RECT 106.1 215.28 106.3 215.4 ;
      RECT 106.46 216.78 106.66 216.9 ;
      RECT 104.3 216.78 104.5 216.9 ;
      RECT 102.86 216.78 103.06 216.9 ;
      RECT 105.74 216.54 105.94 216.66 ;
      RECT 105.02 216.54 105.22 216.66 ;
      RECT 103.58 216.54 103.78 216.66 ;
      RECT 106.46 219.3 106.66 219.42 ;
      RECT 105.74 219.3 105.94 219.42 ;
      RECT 104.3 219.3 104.5 219.42 ;
      RECT 102.86 219.06 103.06 219.18 ;
      RECT 103.58 219.06 103.78 219.18 ;
      RECT 105.02 219.06 105.22 219.18 ;
      RECT 102.86 223.798 103.06 223.918 ;
      RECT 105.02 223.798 105.22 223.918 ;
      RECT 105.74 223.798 105.94 223.918 ;
      RECT 103.58 223.558 103.78 223.678 ;
      RECT 104.3 223.558 104.5 223.678 ;
      RECT 106.46 223.558 106.66 223.678 ;
      RECT 103.22 223.08 103.42 223.2 ;
      RECT 104.66 223.08 104.86 223.2 ;
      RECT 106.1 223.08 106.3 223.2 ;
      RECT 102.5 222.84 102.7 222.96 ;
      RECT 103.94 222.84 104.14 222.96 ;
      RECT 105.38 222.84 105.58 222.96 ;
      RECT 102.86 229.14 103.06 229.26 ;
      RECT 105.02 229.14 105.22 229.26 ;
      RECT 103.58 229.38 103.78 229.5 ;
      RECT 104.3 229.38 104.5 229.5 ;
      RECT 105.74 229.38 105.94 229.5 ;
      RECT 106.46 229.38 106.66 229.5 ;
      RECT 106.46 231.9 106.66 232.02 ;
      RECT 103.58 231.9 103.78 232.02 ;
      RECT 102.86 231.9 103.06 232.02 ;
      RECT 105.74 231.66 105.94 231.78 ;
      RECT 105.02 231.66 105.22 231.78 ;
      RECT 104.3 231.66 104.5 231.78 ;
      RECT 106.46 234.42 106.66 234.54 ;
      RECT 103.58 234.42 103.78 234.54 ;
      RECT 102.86 234.18 103.06 234.3 ;
      RECT 104.3 234.18 104.5 234.3 ;
      RECT 105.02 234.18 105.22 234.3 ;
      RECT 105.74 234.18 105.94 234.3 ;
      RECT 104.3 236.94 104.5 237.06 ;
      RECT 106.46 236.94 106.66 237.06 ;
      RECT 102.86 236.7 103.06 236.82 ;
      RECT 103.58 236.7 103.78 236.82 ;
      RECT 105.02 236.7 105.22 236.82 ;
      RECT 105.74 236.7 105.94 236.82 ;
      RECT 106.46 239.46 106.66 239.58 ;
      RECT 103.58 239.46 103.78 239.58 ;
      RECT 102.86 239.46 103.06 239.58 ;
      RECT 105.74 239.22 105.94 239.34 ;
      RECT 105.02 239.22 105.22 239.34 ;
      RECT 104.3 239.22 104.5 239.34 ;
      RECT 103.58 241.98 103.78 242.1 ;
      RECT 104.3 241.98 104.5 242.1 ;
      RECT 105.02 241.98 105.22 242.1 ;
      RECT 106.46 241.98 106.66 242.1 ;
      RECT 102.86 241.74 103.06 241.86 ;
      RECT 105.74 241.74 105.94 241.86 ;
      RECT 105.02 244.26 105.22 244.38 ;
      RECT 104.3 244.26 104.5 244.38 ;
      RECT 103.58 244.26 103.78 244.38 ;
      RECT 102.86 244.5 103.06 244.62 ;
      RECT 105.74 244.5 105.94 244.62 ;
      RECT 106.46 244.5 106.66 244.62 ;
      RECT 106.46 247.02 106.66 247.14 ;
      RECT 105.74 247.02 105.94 247.14 ;
      RECT 104.3 247.02 104.5 247.14 ;
      RECT 102.86 247.02 103.06 247.14 ;
      RECT 105.02 246.78 105.22 246.9 ;
      RECT 103.58 246.78 103.78 246.9 ;
      RECT 106.46 249.54 106.66 249.66 ;
      RECT 106.46 189.06 106.66 189.18 ;
      RECT 105.74 188.82 105.94 188.94 ;
      RECT 105.02 188.82 105.22 188.94 ;
      RECT 103.58 188.82 103.78 188.94 ;
      RECT 102.86 188.82 103.06 188.94 ;
      RECT 106.1 190.32 106.3 190.44 ;
      RECT 105.38 190.32 105.58 190.44 ;
      RECT 103.94 190.32 104.14 190.44 ;
      RECT 102.5 190.32 102.7 190.44 ;
      RECT 103.22 190.08 103.42 190.2 ;
      RECT 104.66 190.08 104.86 190.2 ;
      RECT 105.02 191.58 105.22 191.7 ;
      RECT 102.86 191.58 103.06 191.7 ;
      RECT 106.46 191.34 106.66 191.46 ;
      RECT 105.74 191.34 105.94 191.46 ;
      RECT 104.3 191.34 104.5 191.46 ;
      RECT 103.58 191.34 103.78 191.46 ;
      RECT 103.94 192.84 104.14 192.96 ;
      RECT 103.22 192.84 103.42 192.96 ;
      RECT 102.5 192.84 102.7 192.96 ;
      RECT 104.66 192.6 104.86 192.72 ;
      RECT 105.38 192.6 105.58 192.72 ;
      RECT 106.1 192.6 106.3 192.72 ;
      RECT 105.74 194.1 105.94 194.22 ;
      RECT 104.3 194.1 104.5 194.22 ;
      RECT 102.86 194.1 103.06 194.22 ;
      RECT 106.46 193.86 106.66 193.98 ;
      RECT 105.02 193.86 105.22 193.98 ;
      RECT 103.58 193.86 103.78 193.98 ;
      RECT 105.38 195.12 105.58 195.24 ;
      RECT 104.66 195.12 104.86 195.24 ;
      RECT 102.5 195.12 102.7 195.24 ;
      RECT 103.22 195.36 103.42 195.48 ;
      RECT 103.94 195.36 104.14 195.48 ;
      RECT 106.1 195.36 106.3 195.48 ;
      RECT 105.74 196.38 105.94 196.5 ;
      RECT 105.02 196.38 105.22 196.5 ;
      RECT 103.58 196.38 103.78 196.5 ;
      RECT 102.86 196.38 103.06 196.5 ;
      RECT 106.46 196.62 106.66 196.74 ;
      RECT 104.3 196.62 104.5 196.74 ;
      RECT 103.22 197.64 103.42 197.76 ;
      RECT 103.94 197.64 104.14 197.76 ;
      RECT 105.38 197.64 105.58 197.76 ;
      RECT 106.1 197.88 106.3 198 ;
      RECT 104.66 197.88 104.86 198 ;
      RECT 102.5 197.88 102.7 198 ;
      RECT 103.58 198.9 103.78 199.02 ;
      RECT 104.3 198.9 104.5 199.02 ;
      RECT 105.02 198.9 105.22 199.02 ;
      RECT 106.46 198.9 106.66 199.02 ;
      RECT 102.86 199.14 103.06 199.26 ;
      RECT 105.74 199.14 105.94 199.26 ;
      RECT 106.1 200.4 106.3 200.52 ;
      RECT 104.66 200.4 104.86 200.52 ;
      RECT 103.94 200.4 104.14 200.52 ;
      RECT 102.5 200.4 102.7 200.52 ;
      RECT 105.38 200.16 105.58 200.28 ;
      RECT 103.22 200.16 103.42 200.28 ;
      RECT 102.86 201.66 103.06 201.78 ;
      RECT 106.46 201.66 106.66 201.78 ;
      RECT 103.58 201.42 103.78 201.54 ;
      RECT 104.3 201.42 104.5 201.54 ;
      RECT 105.02 201.42 105.22 201.54 ;
      RECT 105.74 201.42 105.94 201.54 ;
      RECT 106.1 202.92 106.3 203.04 ;
      RECT 105.38 202.92 105.58 203.04 ;
      RECT 104.66 202.92 104.86 203.04 ;
      RECT 103.94 202.92 104.14 203.04 ;
      RECT 103.22 202.68 103.42 202.8 ;
      RECT 102.5 202.68 102.7 202.8 ;
      RECT 104.3 204.18 104.5 204.3 ;
      RECT 105.74 204.18 105.94 204.3 ;
      RECT 106.46 204.18 106.66 204.3 ;
      RECT 105.02 203.94 105.22 204.06 ;
      RECT 103.58 203.94 103.78 204.06 ;
      RECT 102.86 203.94 103.06 204.06 ;
      RECT 102.5 205.44 102.7 205.56 ;
      RECT 103.94 205.44 104.14 205.56 ;
      RECT 106.1 205.2 106.3 205.32 ;
      RECT 105.38 205.2 105.58 205.32 ;
      RECT 104.66 205.2 104.86 205.32 ;
      RECT 103.22 205.2 103.42 205.32 ;
      RECT 104.3 206.7 104.5 206.82 ;
      RECT 106.46 206.46 106.66 206.58 ;
      RECT 105.74 206.46 105.94 206.58 ;
      RECT 105.02 206.46 105.22 206.58 ;
      RECT 103.58 206.46 103.78 206.58 ;
      RECT 102.86 206.46 103.06 206.58 ;
      RECT 103.94 207.96 104.14 208.08 ;
      RECT 106.1 207.96 106.3 208.08 ;
      RECT 103.22 207.96 103.42 208.08 ;
      RECT 102.5 207.72 102.7 207.84 ;
      RECT 104.66 207.72 104.86 207.84 ;
      RECT 105.38 207.72 105.58 207.84 ;
      RECT 105.02 209.22 105.22 209.34 ;
      RECT 103.58 209.22 103.78 209.34 ;
      RECT 102.86 209.22 103.06 209.34 ;
      RECT 104.3 208.98 104.5 209.1 ;
      RECT 105.74 208.98 105.94 209.1 ;
      RECT 106.46 208.98 106.66 209.1 ;
      RECT 105.74 211.5 105.94 211.62 ;
      RECT 102.5 167.64 102.7 167.76 ;
      RECT 103.22 167.4 103.42 167.52 ;
      RECT 103.94 167.4 104.14 167.52 ;
      RECT 105.38 167.4 105.58 167.52 ;
      RECT 106.1 167.4 106.3 167.52 ;
      RECT 105.02 168.9 105.22 169.02 ;
      RECT 104.3 168.9 104.5 169.02 ;
      RECT 102.86 168.9 103.06 169.02 ;
      RECT 103.58 168.66 103.78 168.78 ;
      RECT 105.74 168.66 105.94 168.78 ;
      RECT 106.46 168.66 106.66 168.78 ;
      RECT 106.1 170.16 106.3 170.28 ;
      RECT 104.66 170.16 104.86 170.28 ;
      RECT 103.94 170.16 104.14 170.28 ;
      RECT 105.38 169.92 105.58 170.04 ;
      RECT 103.22 169.92 103.42 170.04 ;
      RECT 102.5 169.92 102.7 170.04 ;
      RECT 105.74 171.42 105.94 171.54 ;
      RECT 105.02 171.42 105.22 171.54 ;
      RECT 104.3 171.42 104.5 171.54 ;
      RECT 102.86 171.42 103.06 171.54 ;
      RECT 106.46 171.18 106.66 171.3 ;
      RECT 103.58 171.18 103.78 171.3 ;
      RECT 104.66 172.68 104.86 172.8 ;
      RECT 103.22 172.68 103.42 172.8 ;
      RECT 102.5 172.44 102.7 172.56 ;
      RECT 103.94 172.44 104.14 172.56 ;
      RECT 105.38 172.44 105.58 172.56 ;
      RECT 106.1 172.44 106.3 172.56 ;
      RECT 105.74 173.94 105.94 174.06 ;
      RECT 104.3 173.94 104.5 174.06 ;
      RECT 106.46 173.7 106.66 173.82 ;
      RECT 105.02 173.7 105.22 173.82 ;
      RECT 103.58 173.7 103.78 173.82 ;
      RECT 102.86 173.7 103.06 173.82 ;
      RECT 106.1 175.2 106.3 175.32 ;
      RECT 104.66 175.2 104.86 175.32 ;
      RECT 103.22 175.2 103.42 175.32 ;
      RECT 102.5 174.96 102.7 175.08 ;
      RECT 103.94 174.96 104.14 175.08 ;
      RECT 105.38 174.96 105.58 175.08 ;
      RECT 106.46 176.46 106.66 176.58 ;
      RECT 104.3 176.46 104.5 176.58 ;
      RECT 102.86 176.46 103.06 176.58 ;
      RECT 105.74 176.22 105.94 176.34 ;
      RECT 105.02 176.22 105.22 176.34 ;
      RECT 103.58 176.22 103.78 176.34 ;
      RECT 105.02 178.74 105.22 178.86 ;
      RECT 103.58 178.74 103.78 178.86 ;
      RECT 102.86 178.74 103.06 178.86 ;
      RECT 105.74 178.74 105.94 178.86 ;
      RECT 106.46 178.74 106.66 178.86 ;
      RECT 106.1 177.72 106.3 177.84 ;
      RECT 104.66 177.72 104.86 177.84 ;
      RECT 103.22 177.72 103.42 177.84 ;
      RECT 105.38 177.48 105.58 177.6 ;
      RECT 103.94 177.48 104.14 177.6 ;
      RECT 102.5 177.48 102.7 177.6 ;
      RECT 106.1 180 106.3 180.12 ;
      RECT 104.66 180 104.86 180.12 ;
      RECT 104.3 178.98 104.5 179.1 ;
      RECT 105.74 181.5 105.94 181.62 ;
      RECT 104.3 181.5 104.5 181.62 ;
      RECT 102.86 181.5 103.06 181.62 ;
      RECT 103.58 181.26 103.78 181.38 ;
      RECT 105.02 181.26 105.22 181.38 ;
      RECT 106.46 181.26 106.66 181.38 ;
      RECT 105.38 180.24 105.58 180.36 ;
      RECT 103.94 180.24 104.14 180.36 ;
      RECT 103.22 180.24 103.42 180.36 ;
      RECT 102.5 180.24 102.7 180.36 ;
      RECT 106.1 182.76 106.3 182.88 ;
      RECT 103.94 182.76 104.14 182.88 ;
      RECT 103.22 182.76 103.42 182.88 ;
      RECT 102.5 182.76 102.7 182.88 ;
      RECT 105.38 182.52 105.58 182.64 ;
      RECT 104.66 182.52 104.86 182.64 ;
      RECT 106.46 184.02 106.66 184.14 ;
      RECT 103.58 184.02 103.78 184.14 ;
      RECT 102.86 184.02 103.06 184.14 ;
      RECT 104.3 183.78 104.5 183.9 ;
      RECT 105.02 183.78 105.22 183.9 ;
      RECT 105.74 183.78 105.94 183.9 ;
      RECT 103.22 185.28 103.42 185.4 ;
      RECT 104.66 185.28 104.86 185.4 ;
      RECT 106.1 185.28 106.3 185.4 ;
      RECT 105.38 185.04 105.58 185.16 ;
      RECT 103.94 185.04 104.14 185.16 ;
      RECT 102.5 185.04 102.7 185.16 ;
      RECT 102.86 186.54 103.06 186.66 ;
      RECT 105.02 186.54 105.22 186.66 ;
      RECT 106.46 186.54 106.66 186.66 ;
      RECT 105.74 186.3 105.94 186.42 ;
      RECT 104.3 186.3 104.5 186.42 ;
      RECT 103.58 186.3 103.78 186.42 ;
      RECT 103.94 187.8 104.14 187.92 ;
      RECT 103.22 187.8 103.42 187.92 ;
      RECT 102.5 187.56 102.7 187.68 ;
      RECT 104.66 187.56 104.86 187.68 ;
      RECT 105.38 187.56 105.58 187.68 ;
      RECT 106.1 187.56 106.3 187.68 ;
      RECT 104.3 189.06 104.5 189.18 ;
      RECT 103.58 145.98 103.78 146.1 ;
      RECT 104.3 145.98 104.5 146.1 ;
      RECT 105.02 145.98 105.22 146.1 ;
      RECT 105.74 145.98 105.94 146.1 ;
      RECT 106.46 145.98 106.66 146.1 ;
      RECT 102.5 144.96 102.7 145.08 ;
      RECT 103.94 144.96 104.14 145.08 ;
      RECT 103.22 144.72 103.42 144.84 ;
      RECT 104.66 144.72 104.86 144.84 ;
      RECT 105.38 144.72 105.58 144.84 ;
      RECT 106.1 144.72 106.3 144.84 ;
      RECT 106.46 148.74 106.66 148.86 ;
      RECT 104.3 148.74 104.5 148.86 ;
      RECT 102.86 148.74 103.06 148.86 ;
      RECT 103.58 148.5 103.78 148.62 ;
      RECT 105.02 148.5 105.22 148.62 ;
      RECT 105.74 148.5 105.94 148.62 ;
      RECT 103.94 150 104.14 150.12 ;
      RECT 103.22 150 103.42 150.12 ;
      RECT 102.5 150 102.7 150.12 ;
      RECT 106.1 149.76 106.3 149.88 ;
      RECT 105.38 149.76 105.58 149.88 ;
      RECT 104.66 149.76 104.86 149.88 ;
      RECT 104.3 151.26 104.5 151.38 ;
      RECT 102.86 151.26 103.06 151.38 ;
      RECT 106.46 151.02 106.66 151.14 ;
      RECT 105.74 151.02 105.94 151.14 ;
      RECT 105.02 151.02 105.22 151.14 ;
      RECT 103.58 151.02 103.78 151.14 ;
      RECT 105.38 152.52 105.58 152.64 ;
      RECT 103.22 152.52 103.42 152.64 ;
      RECT 102.5 152.52 102.7 152.64 ;
      RECT 106.1 152.28 106.3 152.4 ;
      RECT 104.66 152.28 104.86 152.4 ;
      RECT 103.94 152.28 104.14 152.4 ;
      RECT 106.46 153.78 106.66 153.9 ;
      RECT 104.3 153.78 104.5 153.9 ;
      RECT 102.86 153.78 103.06 153.9 ;
      RECT 103.58 153.54 103.78 153.66 ;
      RECT 105.02 153.54 105.22 153.66 ;
      RECT 105.74 153.54 105.94 153.66 ;
      RECT 105.38 155.04 105.58 155.16 ;
      RECT 104.66 155.04 104.86 155.16 ;
      RECT 103.22 155.04 103.42 155.16 ;
      RECT 102.5 154.8 102.7 154.92 ;
      RECT 103.94 154.8 104.14 154.92 ;
      RECT 106.1 154.8 106.3 154.92 ;
      RECT 106.46 156.3 106.66 156.42 ;
      RECT 105.74 156.3 105.94 156.42 ;
      RECT 104.3 156.3 104.5 156.42 ;
      RECT 102.86 156.3 103.06 156.42 ;
      RECT 105.02 156.06 105.22 156.18 ;
      RECT 103.58 156.06 103.78 156.18 ;
      RECT 105.38 157.56 105.58 157.68 ;
      RECT 104.66 157.56 104.86 157.68 ;
      RECT 103.94 157.56 104.14 157.68 ;
      RECT 102.5 157.56 102.7 157.68 ;
      RECT 106.1 157.32 106.3 157.44 ;
      RECT 103.22 157.32 103.42 157.44 ;
      RECT 106.46 158.82 106.66 158.94 ;
      RECT 105.02 158.82 105.22 158.94 ;
      RECT 103.58 158.82 103.78 158.94 ;
      RECT 102.86 158.58 103.06 158.7 ;
      RECT 104.3 158.58 104.5 158.7 ;
      RECT 105.74 158.58 105.94 158.7 ;
      RECT 105.38 160.08 105.58 160.2 ;
      RECT 104.66 160.08 104.86 160.2 ;
      RECT 102.5 160.08 102.7 160.2 ;
      RECT 106.1 159.84 106.3 159.96 ;
      RECT 103.94 159.84 104.14 159.96 ;
      RECT 103.22 159.84 103.42 159.96 ;
      RECT 102.86 161.1 103.06 161.22 ;
      RECT 103.58 161.1 103.78 161.22 ;
      RECT 104.3 161.1 104.5 161.22 ;
      RECT 105.02 161.1 105.22 161.22 ;
      RECT 105.74 161.1 105.94 161.22 ;
      RECT 106.46 161.1 106.66 161.22 ;
      RECT 102.86 163.62 103.06 163.74 ;
      RECT 104.3 163.62 104.5 163.74 ;
      RECT 105.02 163.62 105.22 163.74 ;
      RECT 105.74 163.62 105.94 163.74 ;
      RECT 103.94 162.6 104.14 162.72 ;
      RECT 103.22 162.6 103.42 162.72 ;
      RECT 102.5 162.6 102.7 162.72 ;
      RECT 104.66 162.6 104.86 162.72 ;
      RECT 105.38 162.6 105.58 162.72 ;
      RECT 106.1 162.6 106.3 162.72 ;
      RECT 103.94 165.12 104.14 165.24 ;
      RECT 102.5 165.12 102.7 165.24 ;
      RECT 105.38 164.88 105.58 165 ;
      RECT 104.66 164.88 104.86 165 ;
      RECT 103.22 164.88 103.42 165 ;
      RECT 106.1 164.88 106.3 165 ;
      RECT 106.46 163.86 106.66 163.98 ;
      RECT 103.58 163.86 103.78 163.98 ;
      RECT 102.86 166.38 103.06 166.5 ;
      RECT 104.3 166.38 104.5 166.5 ;
      RECT 105.02 166.38 105.22 166.5 ;
      RECT 106.46 166.38 106.66 166.5 ;
      RECT 105.74 166.14 105.94 166.26 ;
      RECT 103.58 166.14 103.78 166.26 ;
      RECT 104.66 167.64 104.86 167.76 ;
      RECT 99.98 269.7 100.18 269.82 ;
      RECT 102.14 269.46 102.34 269.58 ;
      RECT 99.26 269.46 99.46 269.58 ;
      RECT 98.54 269.46 98.74 269.58 ;
      RECT 101.78 271.59 101.98 271.71 ;
      RECT 101.06 271.59 101.26 271.71 ;
      RECT 98.9 271.59 99.1 271.71 ;
      RECT 100.34 271.35 100.54 271.47 ;
      RECT 99.62 271.35 99.82 271.47 ;
      RECT 101.78 270.33 101.98 270.45 ;
      RECT 99.62 270.33 99.82 270.45 ;
      RECT 98.9 270.33 99.1 270.45 ;
      RECT 102.14 272.22 102.34 272.34 ;
      RECT 101.42 272.22 101.62 272.34 ;
      RECT 99.26 272.22 99.46 272.34 ;
      RECT 98.54 272.22 98.74 272.34 ;
      RECT 100.7 271.98 100.9 272.1 ;
      RECT 99.98 271.98 100.18 272.1 ;
      RECT 101.42 274.74 101.62 274.86 ;
      RECT 102.14 274.5 102.34 274.62 ;
      RECT 100.7 274.5 100.9 274.62 ;
      RECT 99.98 274.5 100.18 274.62 ;
      RECT 99.26 274.5 99.46 274.62 ;
      RECT 98.54 274.5 98.74 274.62 ;
      RECT 101.42 277.02 101.62 277.14 ;
      RECT 99.98 277.02 100.18 277.14 ;
      RECT 102.14 277.26 102.34 277.38 ;
      RECT 100.7 277.26 100.9 277.38 ;
      RECT 99.26 277.26 99.46 277.38 ;
      RECT 98.54 277.26 98.74 277.38 ;
      RECT 98.54 308.496 98.74 308.616 ;
      RECT 99.26 308.496 99.46 308.616 ;
      RECT 99.98 308.496 100.18 308.616 ;
      RECT 100.7 308.496 100.9 308.616 ;
      RECT 101.42 308.496 101.62 308.616 ;
      RECT 102.14 308.496 102.34 308.616 ;
      RECT 98.9 323.3835 99.1 323.5035 ;
      RECT 99.62 323.3835 99.82 323.5035 ;
      RECT 100.34 323.3835 100.54 323.5035 ;
      RECT 101.06 323.3835 101.26 323.5035 ;
      RECT 101.78 323.3835 101.98 323.5035 ;
      RECT 98.54 325.9425 98.74 326.0625 ;
      RECT 99.26 325.9425 99.46 326.0625 ;
      RECT 99.98 325.9425 100.18 326.0625 ;
      RECT 100.7 325.9425 100.9 326.0625 ;
      RECT 101.42 325.9425 101.62 326.0625 ;
      RECT 102.14 325.9425 102.34 326.0625 ;
      RECT 98.9 348.339 99.1 348.459 ;
      RECT 99.62 348.339 99.82 348.459 ;
      RECT 100.34 348.339 100.54 348.459 ;
      RECT 101.06 348.339 101.26 348.459 ;
      RECT 101.78 348.339 101.98 348.459 ;
      RECT 106.1 127.32 106.3 127.44 ;
      RECT 106.46 128.58 106.66 128.7 ;
      RECT 105.74 128.34 105.94 128.46 ;
      RECT 106.46 130.86 106.66 130.98 ;
      RECT 105.74 130.86 105.94 130.98 ;
      RECT 106.1 129.84 106.3 129.96 ;
      RECT 106.1 132.36 106.3 132.48 ;
      RECT 106.46 133.62 106.66 133.74 ;
      RECT 105.74 133.62 105.94 133.74 ;
      RECT 104.3 133.62 104.5 133.74 ;
      RECT 102.86 133.62 103.06 133.74 ;
      RECT 103.58 133.38 103.78 133.5 ;
      RECT 105.02 133.38 105.22 133.5 ;
      RECT 103.94 134.88 104.14 135 ;
      RECT 103.22 134.88 103.42 135 ;
      RECT 102.5 134.88 102.7 135 ;
      RECT 106.1 134.64 106.3 134.76 ;
      RECT 105.38 134.64 105.58 134.76 ;
      RECT 104.66 134.64 104.86 134.76 ;
      RECT 106.46 134.338 106.66 134.458 ;
      RECT 105.74 134.338 105.94 134.458 ;
      RECT 104.3 134.338 104.5 134.458 ;
      RECT 102.86 134.338 103.06 134.458 ;
      RECT 105.02 134.098 105.22 134.218 ;
      RECT 103.58 134.098 103.78 134.218 ;
      RECT 106.1 135.598 106.3 135.718 ;
      RECT 104.66 135.598 104.86 135.718 ;
      RECT 102.5 135.598 102.7 135.718 ;
      RECT 105.38 135.358 105.58 135.478 ;
      RECT 103.94 135.358 104.14 135.478 ;
      RECT 103.22 135.358 103.42 135.478 ;
      RECT 104.3 141.18 104.5 141.3 ;
      RECT 103.58 141.18 103.78 141.3 ;
      RECT 102.86 140.94 103.06 141.06 ;
      RECT 105.02 140.94 105.22 141.06 ;
      RECT 105.74 140.94 105.94 141.06 ;
      RECT 106.46 140.94 106.66 141.06 ;
      RECT 106.1 142.44 106.3 142.56 ;
      RECT 105.38 142.44 105.58 142.56 ;
      RECT 103.94 142.44 104.14 142.56 ;
      RECT 104.66 142.2 104.86 142.32 ;
      RECT 103.22 142.2 103.42 142.32 ;
      RECT 102.5 142.2 102.7 142.32 ;
      RECT 102.86 143.46 103.06 143.58 ;
      RECT 103.58 143.46 103.78 143.58 ;
      RECT 104.3 143.46 104.5 143.58 ;
      RECT 105.02 143.46 105.22 143.58 ;
      RECT 105.74 143.46 105.94 143.58 ;
      RECT 106.46 143.46 106.66 143.58 ;
      RECT 102.86 145.98 103.06 146.1 ;
      RECT 99.98 241.74 100.18 241.86 ;
      RECT 100.7 241.74 100.9 241.86 ;
      RECT 102.14 241.74 102.34 241.86 ;
      RECT 101.42 244.26 101.62 244.38 ;
      RECT 99.98 244.26 100.18 244.38 ;
      RECT 102.14 244.5 102.34 244.62 ;
      RECT 100.7 244.5 100.9 244.62 ;
      RECT 99.26 244.5 99.46 244.62 ;
      RECT 98.54 244.5 98.74 244.62 ;
      RECT 101.42 247.02 101.62 247.14 ;
      RECT 102.14 246.78 102.34 246.9 ;
      RECT 100.7 246.78 100.9 246.9 ;
      RECT 99.98 246.78 100.18 246.9 ;
      RECT 99.26 246.78 99.46 246.9 ;
      RECT 98.54 246.78 98.74 246.9 ;
      RECT 99.26 249.54 99.46 249.66 ;
      RECT 101.42 249.54 101.62 249.66 ;
      RECT 98.54 249.54 98.74 249.66 ;
      RECT 102.14 249.3 102.34 249.42 ;
      RECT 100.7 249.3 100.9 249.42 ;
      RECT 99.98 249.3 100.18 249.42 ;
      RECT 101.42 252.06 101.62 252.18 ;
      RECT 100.7 252.06 100.9 252.18 ;
      RECT 99.98 252.06 100.18 252.18 ;
      RECT 99.26 252.06 99.46 252.18 ;
      RECT 102.14 251.82 102.34 251.94 ;
      RECT 98.54 251.82 98.74 251.94 ;
      RECT 101.42 254.58 101.62 254.7 ;
      RECT 99.98 254.58 100.18 254.7 ;
      RECT 99.26 254.58 99.46 254.7 ;
      RECT 102.14 254.34 102.34 254.46 ;
      RECT 100.7 254.34 100.9 254.46 ;
      RECT 98.54 254.34 98.74 254.46 ;
      RECT 102.14 257.1 102.34 257.22 ;
      RECT 100.7 257.1 100.9 257.22 ;
      RECT 98.54 257.1 98.74 257.22 ;
      RECT 101.42 256.86 101.62 256.98 ;
      RECT 99.98 256.86 100.18 256.98 ;
      RECT 99.26 256.86 99.46 256.98 ;
      RECT 101.06 258.99 101.26 259.11 ;
      RECT 98.9 258.99 99.1 259.11 ;
      RECT 101.78 258.75 101.98 258.87 ;
      RECT 100.34 258.75 100.54 258.87 ;
      RECT 99.62 258.75 99.82 258.87 ;
      RECT 101.06 260.25 101.26 260.37 ;
      RECT 99.62 260.25 99.82 260.37 ;
      RECT 98.9 260.01 99.1 260.13 ;
      RECT 101.78 260.01 101.98 260.13 ;
      RECT 100.34 260.01 100.54 260.13 ;
      RECT 102.14 259.62 102.34 259.74 ;
      RECT 101.42 259.62 101.62 259.74 ;
      RECT 99.98 259.62 100.18 259.74 ;
      RECT 99.26 259.62 99.46 259.74 ;
      RECT 100.7 259.38 100.9 259.5 ;
      RECT 98.54 259.38 98.74 259.5 ;
      RECT 102.14 261.9 102.34 262.02 ;
      RECT 100.7 261.9 100.9 262.02 ;
      RECT 99.98 261.9 100.18 262.02 ;
      RECT 98.54 261.9 98.74 262.02 ;
      RECT 100.34 261.51 100.54 261.63 ;
      RECT 99.62 261.51 99.82 261.63 ;
      RECT 101.78 261.51 101.98 261.63 ;
      RECT 101.06 261.27 101.26 261.39 ;
      RECT 98.9 261.27 99.1 261.39 ;
      RECT 101.06 262.77 101.26 262.89 ;
      RECT 100.34 262.77 100.54 262.89 ;
      RECT 98.9 262.77 99.1 262.89 ;
      RECT 101.78 262.53 101.98 262.65 ;
      RECT 99.62 262.53 99.82 262.65 ;
      RECT 99.26 262.14 99.46 262.26 ;
      RECT 101.42 262.14 101.62 262.26 ;
      RECT 101.42 264.66 101.62 264.78 ;
      RECT 99.26 264.66 99.46 264.78 ;
      RECT 102.14 264.42 102.34 264.54 ;
      RECT 100.7 264.42 100.9 264.54 ;
      RECT 99.98 264.42 100.18 264.54 ;
      RECT 98.54 264.42 98.74 264.54 ;
      RECT 101.06 264.03 101.26 264.15 ;
      RECT 98.9 264.03 99.1 264.15 ;
      RECT 101.78 263.79 101.98 263.91 ;
      RECT 100.34 263.79 100.54 263.91 ;
      RECT 99.62 263.79 99.82 263.91 ;
      RECT 101.42 267.18 101.62 267.3 ;
      RECT 100.7 267.18 100.9 267.3 ;
      RECT 98.54 267.18 98.74 267.3 ;
      RECT 99.98 266.94 100.18 267.06 ;
      RECT 99.26 266.94 99.46 267.06 ;
      RECT 102.14 266.94 102.34 267.06 ;
      RECT 101.78 266.2885 101.98 266.4085 ;
      RECT 101.06 266.2885 101.26 266.4085 ;
      RECT 100.34 266.2885 100.54 266.4085 ;
      RECT 99.62 266.2885 99.82 266.4085 ;
      RECT 98.9 266.2885 99.1 266.4085 ;
      RECT 99.62 267.81 99.82 267.93 ;
      RECT 100.34 267.81 100.54 267.93 ;
      RECT 101.06 267.81 101.26 267.93 ;
      RECT 98.9 267.81 99.1 267.93 ;
      RECT 101.78 267.81 101.98 267.93 ;
      RECT 101.06 270.09 101.26 270.21 ;
      RECT 100.34 270.09 100.54 270.21 ;
      RECT 101.42 269.7 101.62 269.82 ;
      RECT 100.7 269.7 100.9 269.82 ;
      RECT 101.78 205.2 101.98 205.32 ;
      RECT 100.34 205.2 100.54 205.32 ;
      RECT 99.26 206.7 99.46 206.82 ;
      RECT 99.98 206.7 100.18 206.82 ;
      RECT 100.7 206.7 100.9 206.82 ;
      RECT 102.14 206.7 102.34 206.82 ;
      RECT 101.42 206.46 101.62 206.58 ;
      RECT 98.54 206.46 98.74 206.58 ;
      RECT 101.78 207.96 101.98 208.08 ;
      RECT 99.62 207.96 99.82 208.08 ;
      RECT 98.9 207.72 99.1 207.84 ;
      RECT 100.34 207.72 100.54 207.84 ;
      RECT 101.06 207.72 101.26 207.84 ;
      RECT 101.42 209.22 101.62 209.34 ;
      RECT 99.98 209.22 100.18 209.34 ;
      RECT 99.26 209.22 99.46 209.34 ;
      RECT 98.54 208.98 98.74 209.1 ;
      RECT 100.7 208.98 100.9 209.1 ;
      RECT 102.14 208.98 102.34 209.1 ;
      RECT 101.42 211.5 101.62 211.62 ;
      RECT 100.7 211.5 100.9 211.62 ;
      RECT 99.98 211.5 100.18 211.62 ;
      RECT 98.54 211.5 98.74 211.62 ;
      RECT 101.06 210.48 101.26 210.6 ;
      RECT 101.78 210.48 101.98 210.6 ;
      RECT 98.9 210.48 99.1 210.6 ;
      RECT 99.62 210.48 99.82 210.6 ;
      RECT 100.34 210.24 100.54 210.36 ;
      RECT 100.34 212.76 100.54 212.88 ;
      RECT 101.78 212.76 101.98 212.88 ;
      RECT 102.14 211.74 102.34 211.86 ;
      RECT 99.26 211.74 99.46 211.86 ;
      RECT 101.42 214.26 101.62 214.38 ;
      RECT 102.14 214.02 102.34 214.14 ;
      RECT 100.7 214.02 100.9 214.14 ;
      RECT 99.98 214.02 100.18 214.14 ;
      RECT 99.26 214.02 99.46 214.14 ;
      RECT 98.54 214.02 98.74 214.14 ;
      RECT 98.9 213 99.1 213.12 ;
      RECT 99.62 213 99.82 213.12 ;
      RECT 101.06 213 101.26 213.12 ;
      RECT 101.06 215.52 101.26 215.64 ;
      RECT 100.34 215.52 100.54 215.64 ;
      RECT 98.9 215.52 99.1 215.64 ;
      RECT 99.62 215.28 99.82 215.4 ;
      RECT 101.78 215.28 101.98 215.4 ;
      RECT 101.42 216.78 101.62 216.9 ;
      RECT 100.7 216.78 100.9 216.9 ;
      RECT 99.98 216.78 100.18 216.9 ;
      RECT 102.14 216.54 102.34 216.66 ;
      RECT 99.26 216.54 99.46 216.66 ;
      RECT 98.54 216.54 98.74 216.66 ;
      RECT 101.42 219.3 101.62 219.42 ;
      RECT 100.7 219.3 100.9 219.42 ;
      RECT 99.26 219.3 99.46 219.42 ;
      RECT 98.54 219.3 98.74 219.42 ;
      RECT 99.98 219.06 100.18 219.18 ;
      RECT 102.14 219.06 102.34 219.18 ;
      RECT 99.98 223.798 100.18 223.918 ;
      RECT 101.42 223.798 101.62 223.918 ;
      RECT 98.54 223.558 98.74 223.678 ;
      RECT 99.26 223.558 99.46 223.678 ;
      RECT 100.7 223.558 100.9 223.678 ;
      RECT 102.14 223.558 102.34 223.678 ;
      RECT 99.62 223.08 99.82 223.2 ;
      RECT 100.34 223.08 100.54 223.2 ;
      RECT 101.06 223.08 101.26 223.2 ;
      RECT 98.9 222.84 99.1 222.96 ;
      RECT 101.78 222.84 101.98 222.96 ;
      RECT 99.26 229.14 99.46 229.26 ;
      RECT 99.98 229.14 100.18 229.26 ;
      RECT 102.14 229.14 102.34 229.26 ;
      RECT 98.54 229.38 98.74 229.5 ;
      RECT 100.7 229.38 100.9 229.5 ;
      RECT 101.42 229.38 101.62 229.5 ;
      RECT 102.14 231.9 102.34 232.02 ;
      RECT 98.54 231.9 98.74 232.02 ;
      RECT 101.42 231.66 101.62 231.78 ;
      RECT 100.7 231.66 100.9 231.78 ;
      RECT 99.98 231.66 100.18 231.78 ;
      RECT 99.26 231.66 99.46 231.78 ;
      RECT 99.98 234.42 100.18 234.54 ;
      RECT 100.7 234.42 100.9 234.54 ;
      RECT 98.54 234.18 98.74 234.3 ;
      RECT 99.26 234.18 99.46 234.3 ;
      RECT 101.42 234.18 101.62 234.3 ;
      RECT 102.14 234.18 102.34 234.3 ;
      RECT 99.26 236.94 99.46 237.06 ;
      RECT 101.42 236.94 101.62 237.06 ;
      RECT 102.14 236.94 102.34 237.06 ;
      RECT 98.54 236.7 98.74 236.82 ;
      RECT 99.98 236.7 100.18 236.82 ;
      RECT 100.7 236.7 100.9 236.82 ;
      RECT 101.42 239.46 101.62 239.58 ;
      RECT 99.26 239.46 99.46 239.58 ;
      RECT 98.54 239.46 98.74 239.58 ;
      RECT 102.14 239.22 102.34 239.34 ;
      RECT 100.7 239.22 100.9 239.34 ;
      RECT 99.98 239.22 100.18 239.34 ;
      RECT 99.26 241.98 99.46 242.1 ;
      RECT 101.42 241.98 101.62 242.1 ;
      RECT 98.54 241.74 98.74 241.86 ;
      RECT 101.78 182.76 101.98 182.88 ;
      RECT 101.06 182.76 101.26 182.88 ;
      RECT 98.9 182.76 99.1 182.88 ;
      RECT 100.34 182.52 100.54 182.64 ;
      RECT 99.62 182.52 99.82 182.64 ;
      RECT 98.54 184.02 98.74 184.14 ;
      RECT 99.98 184.02 100.18 184.14 ;
      RECT 99.26 183.78 99.46 183.9 ;
      RECT 100.7 183.78 100.9 183.9 ;
      RECT 101.42 183.78 101.62 183.9 ;
      RECT 102.14 183.78 102.34 183.9 ;
      RECT 98.9 185.28 99.1 185.4 ;
      RECT 100.34 185.28 100.54 185.4 ;
      RECT 101.78 185.04 101.98 185.16 ;
      RECT 101.06 185.04 101.26 185.16 ;
      RECT 99.62 185.04 99.82 185.16 ;
      RECT 99.98 186.54 100.18 186.66 ;
      RECT 101.42 186.54 101.62 186.66 ;
      RECT 102.14 186.3 102.34 186.42 ;
      RECT 100.7 186.3 100.9 186.42 ;
      RECT 99.26 186.3 99.46 186.42 ;
      RECT 98.54 186.3 98.74 186.42 ;
      RECT 101.78 187.8 101.98 187.92 ;
      RECT 99.62 187.8 99.82 187.92 ;
      RECT 98.9 187.56 99.1 187.68 ;
      RECT 100.34 187.56 100.54 187.68 ;
      RECT 101.06 187.56 101.26 187.68 ;
      RECT 98.54 189.06 98.74 189.18 ;
      RECT 99.26 189.06 99.46 189.18 ;
      RECT 101.42 189.06 101.62 189.18 ;
      RECT 102.14 188.82 102.34 188.94 ;
      RECT 100.7 188.82 100.9 188.94 ;
      RECT 99.98 188.82 100.18 188.94 ;
      RECT 101.78 190.32 101.98 190.44 ;
      RECT 98.9 190.08 99.1 190.2 ;
      RECT 99.62 190.08 99.82 190.2 ;
      RECT 100.34 190.08 100.54 190.2 ;
      RECT 101.06 190.08 101.26 190.2 ;
      RECT 101.42 191.58 101.62 191.7 ;
      RECT 100.7 191.58 100.9 191.7 ;
      RECT 98.54 191.58 98.74 191.7 ;
      RECT 102.14 191.34 102.34 191.46 ;
      RECT 99.98 191.34 100.18 191.46 ;
      RECT 99.26 191.34 99.46 191.46 ;
      RECT 101.78 192.84 101.98 192.96 ;
      RECT 101.06 192.84 101.26 192.96 ;
      RECT 99.62 192.84 99.82 192.96 ;
      RECT 98.9 192.84 99.1 192.96 ;
      RECT 100.34 192.6 100.54 192.72 ;
      RECT 99.98 194.1 100.18 194.22 ;
      RECT 98.54 194.1 98.74 194.22 ;
      RECT 102.14 193.86 102.34 193.98 ;
      RECT 101.42 193.86 101.62 193.98 ;
      RECT 100.7 193.86 100.9 193.98 ;
      RECT 99.26 193.86 99.46 193.98 ;
      RECT 101.06 195.12 101.26 195.24 ;
      RECT 99.62 195.12 99.82 195.24 ;
      RECT 101.78 195.36 101.98 195.48 ;
      RECT 100.34 195.36 100.54 195.48 ;
      RECT 98.9 195.36 99.1 195.48 ;
      RECT 99.26 196.38 99.46 196.5 ;
      RECT 98.54 196.38 98.74 196.5 ;
      RECT 99.98 196.62 100.18 196.74 ;
      RECT 100.7 196.62 100.9 196.74 ;
      RECT 101.42 196.62 101.62 196.74 ;
      RECT 102.14 196.62 102.34 196.74 ;
      RECT 99.62 197.64 99.82 197.76 ;
      RECT 100.34 197.64 100.54 197.76 ;
      RECT 101.78 197.64 101.98 197.76 ;
      RECT 101.06 197.88 101.26 198 ;
      RECT 98.9 197.88 99.1 198 ;
      RECT 98.54 198.9 98.74 199.02 ;
      RECT 99.26 198.9 99.46 199.02 ;
      RECT 100.7 198.9 100.9 199.02 ;
      RECT 101.42 198.9 101.62 199.02 ;
      RECT 99.98 199.14 100.18 199.26 ;
      RECT 102.14 199.14 102.34 199.26 ;
      RECT 101.06 200.4 101.26 200.52 ;
      RECT 98.9 200.4 99.1 200.52 ;
      RECT 101.78 200.16 101.98 200.28 ;
      RECT 100.34 200.16 100.54 200.28 ;
      RECT 99.62 200.16 99.82 200.28 ;
      RECT 99.26 201.66 99.46 201.78 ;
      RECT 101.42 201.66 101.62 201.78 ;
      RECT 98.54 201.42 98.74 201.54 ;
      RECT 99.98 201.42 100.18 201.54 ;
      RECT 100.7 201.42 100.9 201.54 ;
      RECT 102.14 201.42 102.34 201.54 ;
      RECT 101.06 202.92 101.26 203.04 ;
      RECT 100.34 202.92 100.54 203.04 ;
      RECT 98.9 202.92 99.1 203.04 ;
      RECT 99.62 202.68 99.82 202.8 ;
      RECT 101.78 202.68 101.98 202.8 ;
      RECT 100.7 204.18 100.9 204.3 ;
      RECT 102.14 204.18 102.34 204.3 ;
      RECT 101.42 203.94 101.62 204.06 ;
      RECT 99.98 203.94 100.18 204.06 ;
      RECT 99.26 203.94 99.46 204.06 ;
      RECT 98.54 203.94 98.74 204.06 ;
      RECT 98.9 205.44 99.1 205.56 ;
      RECT 99.62 205.44 99.82 205.56 ;
      RECT 101.06 205.44 101.26 205.56 ;
      RECT 99.26 158.58 99.46 158.7 ;
      RECT 100.7 158.58 100.9 158.7 ;
      RECT 102.14 158.58 102.34 158.7 ;
      RECT 99.62 160.08 99.82 160.2 ;
      RECT 100.34 160.08 100.54 160.2 ;
      RECT 101.78 159.84 101.98 159.96 ;
      RECT 101.06 159.84 101.26 159.96 ;
      RECT 98.9 159.84 99.1 159.96 ;
      RECT 98.54 161.1 98.74 161.22 ;
      RECT 99.26 161.1 99.46 161.22 ;
      RECT 99.98 161.1 100.18 161.22 ;
      RECT 100.7 161.1 100.9 161.22 ;
      RECT 101.42 161.1 101.62 161.22 ;
      RECT 102.14 161.1 102.34 161.22 ;
      RECT 99.26 163.62 99.46 163.74 ;
      RECT 100.7 163.62 100.9 163.74 ;
      RECT 101.42 163.62 101.62 163.74 ;
      RECT 101.78 162.6 101.98 162.72 ;
      RECT 101.06 162.6 101.26 162.72 ;
      RECT 100.34 162.6 100.54 162.72 ;
      RECT 99.62 162.6 99.82 162.72 ;
      RECT 98.9 162.6 99.1 162.72 ;
      RECT 101.78 165.12 101.98 165.24 ;
      RECT 101.06 165.12 101.26 165.24 ;
      RECT 99.62 165.12 99.82 165.24 ;
      RECT 98.9 165.12 99.1 165.24 ;
      RECT 100.34 164.88 100.54 165 ;
      RECT 102.14 163.86 102.34 163.98 ;
      RECT 99.98 163.86 100.18 163.98 ;
      RECT 98.54 163.86 98.74 163.98 ;
      RECT 100.7 166.38 100.9 166.5 ;
      RECT 101.42 166.38 101.62 166.5 ;
      RECT 102.14 166.38 102.34 166.5 ;
      RECT 99.98 166.14 100.18 166.26 ;
      RECT 99.26 166.14 99.46 166.26 ;
      RECT 98.54 166.14 98.74 166.26 ;
      RECT 101.78 167.64 101.98 167.76 ;
      RECT 98.9 167.64 99.1 167.76 ;
      RECT 99.62 167.4 99.82 167.52 ;
      RECT 100.34 167.4 100.54 167.52 ;
      RECT 101.06 167.4 101.26 167.52 ;
      RECT 102.14 168.9 102.34 169.02 ;
      RECT 99.26 168.9 99.46 169.02 ;
      RECT 98.54 168.66 98.74 168.78 ;
      RECT 99.98 168.66 100.18 168.78 ;
      RECT 100.7 168.66 100.9 168.78 ;
      RECT 101.42 168.66 101.62 168.78 ;
      RECT 101.78 170.16 101.98 170.28 ;
      RECT 101.06 170.16 101.26 170.28 ;
      RECT 98.9 170.16 99.1 170.28 ;
      RECT 100.34 169.92 100.54 170.04 ;
      RECT 99.62 169.92 99.82 170.04 ;
      RECT 102.14 171.42 102.34 171.54 ;
      RECT 100.7 171.42 100.9 171.54 ;
      RECT 99.26 171.42 99.46 171.54 ;
      RECT 101.42 171.18 101.62 171.3 ;
      RECT 99.98 171.18 100.18 171.3 ;
      RECT 98.54 171.18 98.74 171.3 ;
      RECT 101.78 172.68 101.98 172.8 ;
      RECT 100.34 172.68 100.54 172.8 ;
      RECT 99.62 172.68 99.82 172.8 ;
      RECT 101.06 172.44 101.26 172.56 ;
      RECT 98.9 172.44 99.1 172.56 ;
      RECT 102.14 173.94 102.34 174.06 ;
      RECT 100.7 173.94 100.9 174.06 ;
      RECT 99.26 173.94 99.46 174.06 ;
      RECT 101.42 173.7 101.62 173.82 ;
      RECT 99.98 173.7 100.18 173.82 ;
      RECT 98.54 173.7 98.74 173.82 ;
      RECT 101.78 175.2 101.98 175.32 ;
      RECT 100.34 175.2 100.54 175.32 ;
      RECT 98.9 175.2 99.1 175.32 ;
      RECT 99.62 174.96 99.82 175.08 ;
      RECT 101.06 174.96 101.26 175.08 ;
      RECT 99.26 176.46 99.46 176.58 ;
      RECT 98.54 176.46 98.74 176.58 ;
      RECT 102.14 176.22 102.34 176.34 ;
      RECT 101.42 176.22 101.62 176.34 ;
      RECT 100.7 176.22 100.9 176.34 ;
      RECT 99.98 176.22 100.18 176.34 ;
      RECT 100.7 178.74 100.9 178.86 ;
      RECT 99.98 178.74 100.18 178.86 ;
      RECT 98.54 178.74 98.74 178.86 ;
      RECT 101.78 177.72 101.98 177.84 ;
      RECT 100.34 177.72 100.54 177.84 ;
      RECT 98.9 177.72 99.1 177.84 ;
      RECT 101.06 177.48 101.26 177.6 ;
      RECT 99.62 177.48 99.82 177.6 ;
      RECT 101.78 180 101.98 180.12 ;
      RECT 100.34 180 100.54 180.12 ;
      RECT 102.14 178.98 102.34 179.1 ;
      RECT 101.42 178.98 101.62 179.1 ;
      RECT 99.26 178.98 99.46 179.1 ;
      RECT 100.7 181.5 100.9 181.62 ;
      RECT 99.26 181.5 99.46 181.62 ;
      RECT 98.54 181.5 98.74 181.62 ;
      RECT 99.98 181.26 100.18 181.38 ;
      RECT 101.42 181.26 101.62 181.38 ;
      RECT 102.14 181.26 102.34 181.38 ;
      RECT 98.9 180.24 99.1 180.36 ;
      RECT 99.62 180.24 99.82 180.36 ;
      RECT 101.06 180.24 101.26 180.36 ;
      RECT 98.9 132.12 99.1 132.24 ;
      RECT 98.54 131.578 98.74 131.698 ;
      RECT 99.26 131.578 99.46 131.698 ;
      RECT 99.98 131.578 100.18 131.698 ;
      RECT 99.26 131.1 99.46 131.22 ;
      RECT 101.42 133.62 101.62 133.74 ;
      RECT 99.98 133.62 100.18 133.74 ;
      RECT 98.54 133.38 98.74 133.5 ;
      RECT 99.26 133.38 99.46 133.5 ;
      RECT 100.7 133.38 100.9 133.5 ;
      RECT 102.14 133.38 102.34 133.5 ;
      RECT 99.62 134.88 99.82 135 ;
      RECT 101.06 134.88 101.26 135 ;
      RECT 100.34 134.88 100.54 135 ;
      RECT 101.78 134.64 101.98 134.76 ;
      RECT 98.9 134.64 99.1 134.76 ;
      RECT 101.42 134.338 101.62 134.458 ;
      RECT 99.98 134.338 100.18 134.458 ;
      RECT 99.26 134.338 99.46 134.458 ;
      RECT 102.14 134.098 102.34 134.218 ;
      RECT 100.7 134.098 100.9 134.218 ;
      RECT 98.54 134.098 98.74 134.218 ;
      RECT 101.06 135.598 101.26 135.718 ;
      RECT 98.9 135.598 99.1 135.718 ;
      RECT 101.78 135.358 101.98 135.478 ;
      RECT 100.34 135.358 100.54 135.478 ;
      RECT 99.62 135.358 99.82 135.478 ;
      RECT 101.42 141.18 101.62 141.3 ;
      RECT 100.7 141.18 100.9 141.3 ;
      RECT 99.98 141.18 100.18 141.3 ;
      RECT 99.26 141.18 99.46 141.3 ;
      RECT 98.54 140.94 98.74 141.06 ;
      RECT 102.14 140.94 102.34 141.06 ;
      RECT 101.06 142.44 101.26 142.56 ;
      RECT 100.34 142.44 100.54 142.56 ;
      RECT 99.62 142.44 99.82 142.56 ;
      RECT 98.9 142.44 99.1 142.56 ;
      RECT 101.78 142.2 101.98 142.32 ;
      RECT 98.54 143.46 98.74 143.58 ;
      RECT 99.26 143.46 99.46 143.58 ;
      RECT 99.98 143.46 100.18 143.58 ;
      RECT 100.7 143.46 100.9 143.58 ;
      RECT 101.42 143.46 101.62 143.58 ;
      RECT 102.14 143.46 102.34 143.58 ;
      RECT 98.54 145.98 98.74 146.1 ;
      RECT 99.26 145.98 99.46 146.1 ;
      RECT 99.98 145.98 100.18 146.1 ;
      RECT 100.7 145.98 100.9 146.1 ;
      RECT 101.42 145.98 101.62 146.1 ;
      RECT 102.14 145.98 102.34 146.1 ;
      RECT 101.06 144.96 101.26 145.08 ;
      RECT 101.78 144.96 101.98 145.08 ;
      RECT 98.9 144.72 99.1 144.84 ;
      RECT 99.62 144.72 99.82 144.84 ;
      RECT 100.34 144.72 100.54 144.84 ;
      RECT 101.42 148.74 101.62 148.86 ;
      RECT 98.54 148.74 98.74 148.86 ;
      RECT 99.26 148.5 99.46 148.62 ;
      RECT 99.98 148.5 100.18 148.62 ;
      RECT 100.7 148.5 100.9 148.62 ;
      RECT 102.14 148.5 102.34 148.62 ;
      RECT 101.06 150 101.26 150.12 ;
      RECT 99.62 150 99.82 150.12 ;
      RECT 98.9 150 99.1 150.12 ;
      RECT 101.78 149.76 101.98 149.88 ;
      RECT 100.34 149.76 100.54 149.88 ;
      RECT 101.42 151.26 101.62 151.38 ;
      RECT 100.7 151.26 100.9 151.38 ;
      RECT 98.54 151.26 98.74 151.38 ;
      RECT 102.14 151.02 102.34 151.14 ;
      RECT 99.98 151.02 100.18 151.14 ;
      RECT 99.26 151.02 99.46 151.14 ;
      RECT 101.06 152.52 101.26 152.64 ;
      RECT 98.9 152.52 99.1 152.64 ;
      RECT 101.78 152.28 101.98 152.4 ;
      RECT 100.34 152.28 100.54 152.4 ;
      RECT 99.62 152.28 99.82 152.4 ;
      RECT 101.42 153.78 101.62 153.9 ;
      RECT 99.98 153.78 100.18 153.9 ;
      RECT 98.54 153.78 98.74 153.9 ;
      RECT 99.26 153.54 99.46 153.66 ;
      RECT 100.7 153.54 100.9 153.66 ;
      RECT 102.14 153.54 102.34 153.66 ;
      RECT 101.06 155.04 101.26 155.16 ;
      RECT 99.62 155.04 99.82 155.16 ;
      RECT 98.9 155.04 99.1 155.16 ;
      RECT 100.34 154.8 100.54 154.92 ;
      RECT 101.78 154.8 101.98 154.92 ;
      RECT 101.42 156.3 101.62 156.42 ;
      RECT 99.98 156.3 100.18 156.42 ;
      RECT 98.54 156.3 98.74 156.42 ;
      RECT 102.14 156.06 102.34 156.18 ;
      RECT 100.7 156.06 100.9 156.18 ;
      RECT 99.26 156.06 99.46 156.18 ;
      RECT 100.34 157.56 100.54 157.68 ;
      RECT 98.9 157.56 99.1 157.68 ;
      RECT 101.06 157.32 101.26 157.44 ;
      RECT 99.62 157.32 99.82 157.44 ;
      RECT 101.78 157.32 101.98 157.44 ;
      RECT 101.42 158.82 101.62 158.94 ;
      RECT 99.98 158.82 100.18 158.94 ;
      RECT 98.54 158.82 98.74 158.94 ;
      RECT 96.74 264.03 96.94 264.15 ;
      RECT 96.02 264.03 96.22 264.15 ;
      RECT 98.18 263.79 98.38 263.91 ;
      RECT 95.3 263.79 95.5 263.91 ;
      RECT 94.58 263.79 94.78 263.91 ;
      RECT 97.1 267.18 97.3 267.3 ;
      RECT 95.66 267.18 95.86 267.3 ;
      RECT 94.22 267.18 94.42 267.3 ;
      RECT 97.82 266.94 98.02 267.06 ;
      RECT 96.38 266.94 96.58 267.06 ;
      RECT 94.94 266.94 95.14 267.06 ;
      RECT 98.18 266.2885 98.38 266.4085 ;
      RECT 97.46 266.2885 97.66 266.4085 ;
      RECT 96.74 266.2885 96.94 266.4085 ;
      RECT 96.02 266.2885 96.22 266.4085 ;
      RECT 95.3 266.2885 95.5 266.4085 ;
      RECT 94.58 266.2885 94.78 266.4085 ;
      RECT 98.18 267.81 98.38 267.93 ;
      RECT 97.46 267.81 97.66 267.93 ;
      RECT 96.74 267.81 96.94 267.93 ;
      RECT 96.02 267.81 96.22 267.93 ;
      RECT 95.3 267.81 95.5 267.93 ;
      RECT 94.58 267.81 94.78 267.93 ;
      RECT 98.18 270.09 98.38 270.21 ;
      RECT 96.74 270.09 96.94 270.21 ;
      RECT 95.3 270.09 95.5 270.21 ;
      RECT 94.58 270.09 94.78 270.21 ;
      RECT 97.1 269.7 97.3 269.82 ;
      RECT 96.38 269.7 96.58 269.82 ;
      RECT 97.82 269.46 98.02 269.58 ;
      RECT 95.66 269.46 95.86 269.58 ;
      RECT 94.94 269.46 95.14 269.58 ;
      RECT 94.22 269.46 94.42 269.58 ;
      RECT 98.18 271.59 98.38 271.71 ;
      RECT 97.46 271.59 97.66 271.71 ;
      RECT 96.02 271.59 96.22 271.71 ;
      RECT 94.58 271.59 94.78 271.71 ;
      RECT 96.74 271.35 96.94 271.47 ;
      RECT 95.3 271.35 95.5 271.47 ;
      RECT 97.46 270.33 97.66 270.45 ;
      RECT 96.02 270.33 96.22 270.45 ;
      RECT 94.22 272.22 94.42 272.34 ;
      RECT 96.38 272.22 96.58 272.34 ;
      RECT 97.82 271.98 98.02 272.1 ;
      RECT 97.1 271.98 97.3 272.1 ;
      RECT 95.66 271.98 95.86 272.1 ;
      RECT 94.94 271.98 95.14 272.1 ;
      RECT 97.82 274.74 98.02 274.86 ;
      RECT 95.66 274.74 95.86 274.86 ;
      RECT 94.94 274.74 95.14 274.86 ;
      RECT 94.22 274.74 94.42 274.86 ;
      RECT 97.1 274.5 97.3 274.62 ;
      RECT 96.38 274.5 96.58 274.62 ;
      RECT 97.82 277.02 98.02 277.14 ;
      RECT 96.38 277.02 96.58 277.14 ;
      RECT 94.94 277.02 95.14 277.14 ;
      RECT 94.22 277.02 94.42 277.14 ;
      RECT 97.1 277.26 97.3 277.38 ;
      RECT 95.66 277.26 95.86 277.38 ;
      RECT 94.22 308.496 94.42 308.616 ;
      RECT 94.94 308.496 95.14 308.616 ;
      RECT 95.66 308.496 95.86 308.616 ;
      RECT 96.38 308.496 96.58 308.616 ;
      RECT 97.1 308.496 97.3 308.616 ;
      RECT 97.82 308.496 98.02 308.616 ;
      RECT 94.58 323.3835 94.78 323.5035 ;
      RECT 95.3 323.3835 95.5 323.5035 ;
      RECT 96.02 323.3835 96.22 323.5035 ;
      RECT 96.74 323.3835 96.94 323.5035 ;
      RECT 97.46 323.3835 97.66 323.5035 ;
      RECT 98.18 323.3835 98.38 323.5035 ;
      RECT 96.38 325.9425 96.58 326.0625 ;
      RECT 95.66 325.9425 95.86 326.0625 ;
      RECT 94.94 325.9425 95.14 326.0625 ;
      RECT 94.22 325.9425 94.42 326.0625 ;
      RECT 97.1 325.9425 97.3 326.0625 ;
      RECT 97.82 325.9425 98.02 326.0625 ;
      RECT 94.58 348.339 94.78 348.459 ;
      RECT 95.3 348.339 95.5 348.459 ;
      RECT 96.02 348.339 96.22 348.459 ;
      RECT 96.74 348.339 96.94 348.459 ;
      RECT 97.46 348.339 97.66 348.459 ;
      RECT 98.18 348.339 98.38 348.459 ;
      RECT 98.54 126.538 98.74 126.658 ;
      RECT 99.26 126.538 99.46 126.658 ;
      RECT 99.98 126.538 100.18 126.658 ;
      RECT 100.7 126.538 100.9 126.658 ;
      RECT 101.42 126.538 101.62 126.658 ;
      RECT 102.14 126.538 102.34 126.658 ;
      RECT 99.62 127.32 99.82 127.44 ;
      RECT 98.9 127.08 99.1 127.2 ;
      RECT 98.54 129.058 98.74 129.178 ;
      RECT 99.26 129.058 99.46 129.178 ;
      RECT 99.98 129.058 100.18 129.178 ;
      RECT 99.26 128.58 99.46 128.7 ;
      RECT 99.98 128.34 100.18 128.46 ;
      RECT 98.54 128.34 98.74 128.46 ;
      RECT 99.98 130.86 100.18 130.98 ;
      RECT 98.54 130.86 98.74 130.98 ;
      RECT 98.9 129.84 99.1 129.96 ;
      RECT 99.62 129.84 99.82 129.96 ;
      RECT 99.62 132.36 99.82 132.48 ;
      RECT 95.66 234.42 95.86 234.54 ;
      RECT 94.22 234.42 94.42 234.54 ;
      RECT 94.94 234.18 95.14 234.3 ;
      RECT 96.38 234.18 96.58 234.3 ;
      RECT 97.1 234.18 97.3 234.3 ;
      RECT 94.94 236.94 95.14 237.06 ;
      RECT 96.38 236.94 96.58 237.06 ;
      RECT 97.1 236.94 97.3 237.06 ;
      RECT 94.22 236.7 94.42 236.82 ;
      RECT 95.66 236.7 95.86 236.82 ;
      RECT 97.82 236.7 98.02 236.82 ;
      RECT 96.38 239.46 96.58 239.58 ;
      RECT 95.66 239.46 95.86 239.58 ;
      RECT 94.94 239.46 95.14 239.58 ;
      RECT 97.82 239.22 98.02 239.34 ;
      RECT 97.1 239.22 97.3 239.34 ;
      RECT 94.22 239.22 94.42 239.34 ;
      RECT 94.22 241.98 94.42 242.1 ;
      RECT 94.94 241.98 95.14 242.1 ;
      RECT 95.66 241.98 95.86 242.1 ;
      RECT 96.38 241.98 96.58 242.1 ;
      RECT 97.82 241.98 98.02 242.1 ;
      RECT 97.1 241.74 97.3 241.86 ;
      RECT 97.82 244.26 98.02 244.38 ;
      RECT 97.1 244.26 97.3 244.38 ;
      RECT 96.38 244.26 96.58 244.38 ;
      RECT 95.66 244.26 95.86 244.38 ;
      RECT 94.22 244.26 94.42 244.38 ;
      RECT 94.94 244.5 95.14 244.62 ;
      RECT 97.82 247.02 98.02 247.14 ;
      RECT 97.1 247.02 97.3 247.14 ;
      RECT 96.38 247.02 96.58 247.14 ;
      RECT 95.66 247.02 95.86 247.14 ;
      RECT 94.94 247.02 95.14 247.14 ;
      RECT 94.22 246.78 94.42 246.9 ;
      RECT 95.66 249.54 95.86 249.66 ;
      RECT 94.94 249.54 95.14 249.66 ;
      RECT 97.82 249.3 98.02 249.42 ;
      RECT 97.1 249.3 97.3 249.42 ;
      RECT 96.38 249.3 96.58 249.42 ;
      RECT 94.22 249.3 94.42 249.42 ;
      RECT 97.1 252.06 97.3 252.18 ;
      RECT 95.66 252.06 95.86 252.18 ;
      RECT 94.22 252.06 94.42 252.18 ;
      RECT 97.82 251.82 98.02 251.94 ;
      RECT 96.38 251.82 96.58 251.94 ;
      RECT 94.94 251.82 95.14 251.94 ;
      RECT 97.1 254.58 97.3 254.7 ;
      RECT 95.66 254.58 95.86 254.7 ;
      RECT 94.94 254.58 95.14 254.7 ;
      RECT 94.22 254.58 94.42 254.7 ;
      RECT 97.82 254.34 98.02 254.46 ;
      RECT 96.38 254.34 96.58 254.46 ;
      RECT 97.82 257.1 98.02 257.22 ;
      RECT 96.38 257.1 96.58 257.22 ;
      RECT 94.22 257.1 94.42 257.22 ;
      RECT 97.1 256.86 97.3 256.98 ;
      RECT 95.66 256.86 95.86 256.98 ;
      RECT 94.94 256.86 95.14 256.98 ;
      RECT 97.46 258.99 97.66 259.11 ;
      RECT 96.74 258.99 96.94 259.11 ;
      RECT 96.02 258.99 96.22 259.11 ;
      RECT 94.58 258.99 94.78 259.11 ;
      RECT 98.18 258.75 98.38 258.87 ;
      RECT 95.3 258.75 95.5 258.87 ;
      RECT 98.18 260.25 98.38 260.37 ;
      RECT 94.58 260.25 94.78 260.37 ;
      RECT 97.46 260.01 97.66 260.13 ;
      RECT 96.74 260.01 96.94 260.13 ;
      RECT 96.02 260.01 96.22 260.13 ;
      RECT 95.3 260.01 95.5 260.13 ;
      RECT 97.1 259.62 97.3 259.74 ;
      RECT 95.66 259.62 95.86 259.74 ;
      RECT 97.82 259.38 98.02 259.5 ;
      RECT 96.38 259.38 96.58 259.5 ;
      RECT 94.94 259.38 95.14 259.5 ;
      RECT 94.22 259.38 94.42 259.5 ;
      RECT 97.1 261.9 97.3 262.02 ;
      RECT 96.38 261.9 96.58 262.02 ;
      RECT 94.94 261.9 95.14 262.02 ;
      RECT 98.18 261.51 98.38 261.63 ;
      RECT 96.02 261.51 96.22 261.63 ;
      RECT 95.3 261.51 95.5 261.63 ;
      RECT 97.46 261.27 97.66 261.39 ;
      RECT 96.74 261.27 96.94 261.39 ;
      RECT 94.58 261.27 94.78 261.39 ;
      RECT 97.46 262.77 97.66 262.89 ;
      RECT 96.02 262.77 96.22 262.89 ;
      RECT 95.3 262.77 95.5 262.89 ;
      RECT 94.58 262.77 94.78 262.89 ;
      RECT 98.18 262.53 98.38 262.65 ;
      RECT 96.74 262.53 96.94 262.65 ;
      RECT 97.82 262.14 98.02 262.26 ;
      RECT 95.66 262.14 95.86 262.26 ;
      RECT 94.22 262.14 94.42 262.26 ;
      RECT 97.1 264.66 97.3 264.78 ;
      RECT 96.38 264.66 96.58 264.78 ;
      RECT 94.94 264.66 95.14 264.78 ;
      RECT 94.22 264.66 94.42 264.78 ;
      RECT 97.82 264.42 98.02 264.54 ;
      RECT 95.66 264.42 95.86 264.54 ;
      RECT 97.46 264.03 97.66 264.15 ;
      RECT 96.74 202.68 96.94 202.8 ;
      RECT 96.02 202.68 96.22 202.8 ;
      RECT 94.58 202.68 94.78 202.8 ;
      RECT 95.3 202.92 95.5 203.04 ;
      RECT 98.18 202.92 98.38 203.04 ;
      RECT 94.94 203.94 95.14 204.06 ;
      RECT 97.82 204.18 98.02 204.3 ;
      RECT 97.1 204.18 97.3 204.3 ;
      RECT 96.38 204.18 96.58 204.3 ;
      RECT 95.66 204.18 95.86 204.3 ;
      RECT 94.22 204.18 94.42 204.3 ;
      RECT 94.58 205.2 94.78 205.32 ;
      RECT 97.46 205.2 97.66 205.32 ;
      RECT 98.18 205.44 98.38 205.56 ;
      RECT 96.74 205.44 96.94 205.56 ;
      RECT 96.02 205.44 96.22 205.56 ;
      RECT 95.3 205.44 95.5 205.56 ;
      RECT 94.22 206.46 94.42 206.58 ;
      RECT 94.94 206.46 95.14 206.58 ;
      RECT 95.66 206.46 95.86 206.58 ;
      RECT 96.38 206.46 96.58 206.58 ;
      RECT 97.1 206.46 97.3 206.58 ;
      RECT 97.82 206.7 98.02 206.82 ;
      RECT 98.18 207.72 98.38 207.84 ;
      RECT 97.46 207.72 97.66 207.84 ;
      RECT 94.58 207.72 94.78 207.84 ;
      RECT 95.3 207.96 95.5 208.08 ;
      RECT 96.02 207.96 96.22 208.08 ;
      RECT 96.74 207.96 96.94 208.08 ;
      RECT 97.1 208.98 97.3 209.1 ;
      RECT 95.66 208.98 95.86 209.1 ;
      RECT 94.94 208.98 95.14 209.1 ;
      RECT 94.22 209.22 94.42 209.34 ;
      RECT 96.38 209.22 96.58 209.34 ;
      RECT 97.82 209.22 98.02 209.34 ;
      RECT 97.1 211.5 97.3 211.62 ;
      RECT 96.38 211.5 96.58 211.62 ;
      RECT 94.94 211.5 95.14 211.62 ;
      RECT 95.3 210.48 95.5 210.6 ;
      RECT 96.02 210.48 96.22 210.6 ;
      RECT 98.18 210.48 98.38 210.6 ;
      RECT 94.58 210.24 94.78 210.36 ;
      RECT 96.74 210.24 96.94 210.36 ;
      RECT 97.46 210.24 97.66 210.36 ;
      RECT 96.02 212.76 96.22 212.88 ;
      RECT 96.74 212.76 96.94 212.88 ;
      RECT 97.46 212.76 97.66 212.88 ;
      RECT 97.82 211.74 98.02 211.86 ;
      RECT 95.66 211.74 95.86 211.86 ;
      RECT 94.22 211.74 94.42 211.86 ;
      RECT 97.82 214.26 98.02 214.38 ;
      RECT 95.66 214.26 95.86 214.38 ;
      RECT 94.22 214.26 94.42 214.38 ;
      RECT 97.1 214.02 97.3 214.14 ;
      RECT 96.38 214.02 96.58 214.14 ;
      RECT 94.94 214.02 95.14 214.14 ;
      RECT 98.18 213 98.38 213.12 ;
      RECT 95.3 213 95.5 213.12 ;
      RECT 94.58 213 94.78 213.12 ;
      RECT 97.46 215.52 97.66 215.64 ;
      RECT 95.3 215.52 95.5 215.64 ;
      RECT 94.58 215.52 94.78 215.64 ;
      RECT 96.02 215.28 96.22 215.4 ;
      RECT 96.74 215.28 96.94 215.4 ;
      RECT 98.18 215.28 98.38 215.4 ;
      RECT 97.82 216.78 98.02 216.9 ;
      RECT 97.1 216.78 97.3 216.9 ;
      RECT 95.66 216.78 95.86 216.9 ;
      RECT 94.22 216.78 94.42 216.9 ;
      RECT 96.38 216.54 96.58 216.66 ;
      RECT 94.94 216.54 95.14 216.66 ;
      RECT 97.1 219.3 97.3 219.42 ;
      RECT 95.66 219.3 95.86 219.42 ;
      RECT 94.22 219.06 94.42 219.18 ;
      RECT 94.94 219.06 95.14 219.18 ;
      RECT 96.38 219.06 96.58 219.18 ;
      RECT 97.82 219.06 98.02 219.18 ;
      RECT 95.66 223.798 95.86 223.918 ;
      RECT 96.38 223.798 96.58 223.918 ;
      RECT 97.1 223.798 97.3 223.918 ;
      RECT 94.22 223.558 94.42 223.678 ;
      RECT 94.94 223.558 95.14 223.678 ;
      RECT 97.82 223.558 98.02 223.678 ;
      RECT 94.58 223.08 94.78 223.2 ;
      RECT 96.02 223.08 96.22 223.2 ;
      RECT 96.74 223.08 96.94 223.2 ;
      RECT 97.46 223.08 97.66 223.2 ;
      RECT 95.3 222.84 95.5 222.96 ;
      RECT 98.18 222.84 98.38 222.96 ;
      RECT 94.22 229.14 94.42 229.26 ;
      RECT 95.66 229.14 95.86 229.26 ;
      RECT 96.38 229.14 96.58 229.26 ;
      RECT 97.1 229.14 97.3 229.26 ;
      RECT 94.94 229.38 95.14 229.5 ;
      RECT 97.82 229.38 98.02 229.5 ;
      RECT 97.82 231.9 98.02 232.02 ;
      RECT 96.38 231.9 96.58 232.02 ;
      RECT 97.1 231.66 97.3 231.78 ;
      RECT 95.66 231.66 95.86 231.78 ;
      RECT 94.94 231.66 95.14 231.78 ;
      RECT 94.22 231.66 94.42 231.78 ;
      RECT 97.82 234.42 98.02 234.54 ;
      RECT 96.38 181.26 96.58 181.38 ;
      RECT 95.66 181.26 95.86 181.38 ;
      RECT 94.94 181.26 95.14 181.38 ;
      RECT 96.02 180.24 96.22 180.36 ;
      RECT 95.3 180.24 95.5 180.36 ;
      RECT 96.74 182.76 96.94 182.88 ;
      RECT 96.02 182.76 96.22 182.88 ;
      RECT 95.3 182.76 95.5 182.88 ;
      RECT 98.18 182.52 98.38 182.64 ;
      RECT 97.46 182.52 97.66 182.64 ;
      RECT 94.58 182.52 94.78 182.64 ;
      RECT 96.38 184.02 96.58 184.14 ;
      RECT 94.94 184.02 95.14 184.14 ;
      RECT 94.22 184.02 94.42 184.14 ;
      RECT 95.66 183.78 95.86 183.9 ;
      RECT 97.1 183.78 97.3 183.9 ;
      RECT 97.82 183.78 98.02 183.9 ;
      RECT 95.3 185.28 95.5 185.4 ;
      RECT 96.74 185.28 96.94 185.4 ;
      RECT 97.46 185.28 97.66 185.4 ;
      RECT 98.18 185.04 98.38 185.16 ;
      RECT 96.02 185.04 96.22 185.16 ;
      RECT 94.58 185.04 94.78 185.16 ;
      RECT 94.22 186.54 94.42 186.66 ;
      RECT 95.66 186.54 95.86 186.66 ;
      RECT 97.1 186.54 97.3 186.66 ;
      RECT 97.82 186.3 98.02 186.42 ;
      RECT 96.38 186.3 96.58 186.42 ;
      RECT 94.94 186.3 95.14 186.42 ;
      RECT 96.74 187.8 96.94 187.92 ;
      RECT 96.02 187.8 96.22 187.92 ;
      RECT 94.58 187.8 94.78 187.92 ;
      RECT 95.3 187.56 95.5 187.68 ;
      RECT 97.46 187.56 97.66 187.68 ;
      RECT 98.18 187.56 98.38 187.68 ;
      RECT 94.22 189.06 94.42 189.18 ;
      RECT 95.66 189.06 95.86 189.18 ;
      RECT 97.82 189.06 98.02 189.18 ;
      RECT 97.1 188.82 97.3 188.94 ;
      RECT 96.38 188.82 96.58 188.94 ;
      RECT 94.94 188.82 95.14 188.94 ;
      RECT 98.18 190.32 98.38 190.44 ;
      RECT 96.74 190.32 96.94 190.44 ;
      RECT 96.02 190.32 96.22 190.44 ;
      RECT 95.3 190.32 95.5 190.44 ;
      RECT 94.58 190.32 94.78 190.44 ;
      RECT 97.46 190.08 97.66 190.2 ;
      RECT 97.1 191.58 97.3 191.7 ;
      RECT 96.38 191.58 96.58 191.7 ;
      RECT 95.66 191.58 95.86 191.7 ;
      RECT 94.94 191.58 95.14 191.7 ;
      RECT 97.82 191.34 98.02 191.46 ;
      RECT 94.22 191.34 94.42 191.46 ;
      RECT 96.02 192.84 96.22 192.96 ;
      RECT 94.58 192.6 94.78 192.72 ;
      RECT 95.3 192.6 95.5 192.72 ;
      RECT 96.74 192.6 96.94 192.72 ;
      RECT 97.46 192.6 97.66 192.72 ;
      RECT 98.18 192.6 98.38 192.72 ;
      RECT 97.1 194.1 97.3 194.22 ;
      RECT 95.66 194.1 95.86 194.22 ;
      RECT 94.94 194.1 95.14 194.22 ;
      RECT 97.82 193.86 98.02 193.98 ;
      RECT 96.38 193.86 96.58 193.98 ;
      RECT 94.22 193.86 94.42 193.98 ;
      RECT 98.18 195.12 98.38 195.24 ;
      RECT 96.74 195.12 96.94 195.24 ;
      RECT 95.3 195.12 95.5 195.24 ;
      RECT 97.46 195.36 97.66 195.48 ;
      RECT 96.02 195.36 96.22 195.48 ;
      RECT 94.58 195.36 94.78 195.48 ;
      RECT 97.1 196.38 97.3 196.5 ;
      RECT 94.94 196.38 95.14 196.5 ;
      RECT 94.22 196.62 94.42 196.74 ;
      RECT 95.66 196.62 95.86 196.74 ;
      RECT 96.38 196.62 96.58 196.74 ;
      RECT 97.82 196.62 98.02 196.74 ;
      RECT 96.74 197.64 96.94 197.76 ;
      RECT 98.18 197.64 98.38 197.76 ;
      RECT 97.46 197.88 97.66 198 ;
      RECT 96.02 197.88 96.22 198 ;
      RECT 95.3 197.88 95.5 198 ;
      RECT 94.58 197.88 94.78 198 ;
      RECT 94.22 198.9 94.42 199.02 ;
      RECT 94.94 198.9 95.14 199.02 ;
      RECT 95.66 198.9 95.86 199.02 ;
      RECT 96.38 199.14 96.58 199.26 ;
      RECT 97.1 199.14 97.3 199.26 ;
      RECT 97.82 199.14 98.02 199.26 ;
      RECT 95.3 200.16 95.5 200.28 ;
      RECT 96.74 200.16 96.94 200.28 ;
      RECT 94.58 200.4 94.78 200.52 ;
      RECT 96.02 200.4 96.22 200.52 ;
      RECT 97.46 200.4 97.66 200.52 ;
      RECT 98.18 200.4 98.38 200.52 ;
      RECT 96.38 201.42 96.58 201.54 ;
      RECT 94.22 201.42 94.42 201.54 ;
      RECT 97.82 201.66 98.02 201.78 ;
      RECT 97.1 201.66 97.3 201.78 ;
      RECT 95.66 201.66 95.86 201.78 ;
      RECT 94.94 201.66 95.14 201.78 ;
      RECT 97.46 202.68 97.66 202.8 ;
      RECT 96.02 160.08 96.22 160.2 ;
      RECT 97.46 160.08 97.66 160.2 ;
      RECT 98.18 160.08 98.38 160.2 ;
      RECT 96.74 159.84 96.94 159.96 ;
      RECT 95.3 159.84 95.5 159.96 ;
      RECT 94.22 161.1 94.42 161.22 ;
      RECT 94.94 161.1 95.14 161.22 ;
      RECT 95.66 161.1 95.86 161.22 ;
      RECT 96.38 161.1 96.58 161.22 ;
      RECT 97.1 161.1 97.3 161.22 ;
      RECT 97.82 161.1 98.02 161.22 ;
      RECT 94.22 163.62 94.42 163.74 ;
      RECT 94.94 163.62 95.14 163.74 ;
      RECT 95.66 163.62 95.86 163.74 ;
      RECT 96.38 163.62 96.58 163.74 ;
      RECT 97.82 163.62 98.02 163.74 ;
      RECT 98.18 162.6 98.38 162.72 ;
      RECT 97.46 162.6 97.66 162.72 ;
      RECT 96.02 162.6 96.22 162.72 ;
      RECT 94.58 162.6 94.78 162.72 ;
      RECT 96.74 162.6 96.94 162.72 ;
      RECT 95.3 162.6 95.5 162.72 ;
      RECT 97.46 165.12 97.66 165.24 ;
      RECT 95.3 165.12 95.5 165.24 ;
      RECT 98.18 164.88 98.38 165 ;
      RECT 96.74 164.88 96.94 165 ;
      RECT 96.02 164.88 96.22 165 ;
      RECT 94.58 164.88 94.78 165 ;
      RECT 97.1 163.86 97.3 163.98 ;
      RECT 94.22 166.38 94.42 166.5 ;
      RECT 96.38 166.38 96.58 166.5 ;
      RECT 97.82 166.38 98.02 166.5 ;
      RECT 97.1 166.14 97.3 166.26 ;
      RECT 95.66 166.14 95.86 166.26 ;
      RECT 94.94 166.14 95.14 166.26 ;
      RECT 97.46 167.64 97.66 167.76 ;
      RECT 96.74 167.64 96.94 167.76 ;
      RECT 96.02 167.64 96.22 167.76 ;
      RECT 95.3 167.64 95.5 167.76 ;
      RECT 94.58 167.64 94.78 167.76 ;
      RECT 98.18 167.4 98.38 167.52 ;
      RECT 97.82 168.9 98.02 169.02 ;
      RECT 97.1 168.9 97.3 169.02 ;
      RECT 96.38 168.9 96.58 169.02 ;
      RECT 94.22 168.66 94.42 168.78 ;
      RECT 94.94 168.66 95.14 168.78 ;
      RECT 95.66 168.66 95.86 168.78 ;
      RECT 97.46 170.16 97.66 170.28 ;
      RECT 96.02 170.16 96.22 170.28 ;
      RECT 95.3 170.16 95.5 170.28 ;
      RECT 98.18 169.92 98.38 170.04 ;
      RECT 96.74 169.92 96.94 170.04 ;
      RECT 94.58 169.92 94.78 170.04 ;
      RECT 95.66 171.42 95.86 171.54 ;
      RECT 97.82 171.42 98.02 171.54 ;
      RECT 97.1 171.18 97.3 171.3 ;
      RECT 96.38 171.18 96.58 171.3 ;
      RECT 94.94 171.18 95.14 171.3 ;
      RECT 94.22 171.18 94.42 171.3 ;
      RECT 97.46 172.68 97.66 172.8 ;
      RECT 96.74 172.68 96.94 172.8 ;
      RECT 95.3 172.68 95.5 172.8 ;
      RECT 94.58 172.44 94.78 172.56 ;
      RECT 96.02 172.44 96.22 172.56 ;
      RECT 98.18 172.44 98.38 172.56 ;
      RECT 97.1 173.94 97.3 174.06 ;
      RECT 95.66 173.94 95.86 174.06 ;
      RECT 94.22 173.94 94.42 174.06 ;
      RECT 97.82 173.7 98.02 173.82 ;
      RECT 96.38 173.7 96.58 173.82 ;
      RECT 94.94 173.7 95.14 173.82 ;
      RECT 97.46 175.2 97.66 175.32 ;
      RECT 95.3 175.2 95.5 175.32 ;
      RECT 94.58 174.96 94.78 175.08 ;
      RECT 96.02 174.96 96.22 175.08 ;
      RECT 96.74 174.96 96.94 175.08 ;
      RECT 98.18 174.96 98.38 175.08 ;
      RECT 97.82 176.46 98.02 176.58 ;
      RECT 97.1 176.46 97.3 176.58 ;
      RECT 94.22 176.46 94.42 176.58 ;
      RECT 96.38 176.22 96.58 176.34 ;
      RECT 95.66 176.22 95.86 176.34 ;
      RECT 94.94 176.22 95.14 176.34 ;
      RECT 94.94 178.74 95.14 178.86 ;
      RECT 94.22 178.74 94.42 178.86 ;
      RECT 97.46 177.72 97.66 177.84 ;
      RECT 94.58 177.72 94.78 177.84 ;
      RECT 98.18 177.48 98.38 177.6 ;
      RECT 96.74 177.48 96.94 177.6 ;
      RECT 96.02 177.48 96.22 177.6 ;
      RECT 95.3 177.48 95.5 177.6 ;
      RECT 98.18 180 98.38 180.12 ;
      RECT 97.46 180 97.66 180.12 ;
      RECT 96.74 180 96.94 180.12 ;
      RECT 94.58 180 94.78 180.12 ;
      RECT 97.82 178.98 98.02 179.1 ;
      RECT 97.1 178.98 97.3 179.1 ;
      RECT 96.38 178.98 96.58 179.1 ;
      RECT 95.66 178.98 95.86 179.1 ;
      RECT 97.82 181.5 98.02 181.62 ;
      RECT 94.22 181.5 94.42 181.62 ;
      RECT 97.1 181.26 97.3 181.38 ;
      RECT 98.18 134.64 98.38 134.76 ;
      RECT 96.02 134.64 96.22 134.76 ;
      RECT 97.82 134.338 98.02 134.458 ;
      RECT 97.1 134.338 97.3 134.458 ;
      RECT 94.22 134.098 94.42 134.218 ;
      RECT 96.38 134.098 96.58 134.218 ;
      RECT 95.66 134.098 95.86 134.218 ;
      RECT 94.94 136.14 95.14 136.26 ;
      RECT 94.22 136.14 94.42 136.26 ;
      RECT 96.02 135.598 96.22 135.718 ;
      RECT 95.3 135.598 95.5 135.718 ;
      RECT 98.18 135.358 98.38 135.478 ;
      RECT 97.46 135.358 97.66 135.478 ;
      RECT 96.74 135.358 96.94 135.478 ;
      RECT 94.22 136.858 94.42 136.978 ;
      RECT 94.94 139.138 95.14 139.258 ;
      RECT 94.22 138.42 94.42 138.54 ;
      RECT 94.22 139.378 94.42 139.498 ;
      RECT 94.22 141.18 94.42 141.3 ;
      RECT 97.82 141.18 98.02 141.3 ;
      RECT 95.66 141.18 95.86 141.3 ;
      RECT 96.38 140.94 96.58 141.06 ;
      RECT 97.1 140.94 97.3 141.06 ;
      RECT 96.74 142.44 96.94 142.56 ;
      RECT 96.02 142.44 96.22 142.56 ;
      RECT 98.18 142.2 98.38 142.32 ;
      RECT 97.46 142.2 97.66 142.32 ;
      RECT 95.3 142.2 95.5 142.32 ;
      RECT 94.58 142.2 94.78 142.32 ;
      RECT 94.22 143.46 94.42 143.58 ;
      RECT 94.94 143.46 95.14 143.58 ;
      RECT 95.66 143.46 95.86 143.58 ;
      RECT 96.38 143.46 96.58 143.58 ;
      RECT 97.1 143.46 97.3 143.58 ;
      RECT 97.82 143.46 98.02 143.58 ;
      RECT 94.22 145.98 94.42 146.1 ;
      RECT 94.94 145.98 95.14 146.1 ;
      RECT 95.66 145.98 95.86 146.1 ;
      RECT 96.38 145.98 96.58 146.1 ;
      RECT 97.1 145.98 97.3 146.1 ;
      RECT 97.82 145.98 98.02 146.1 ;
      RECT 96.74 144.96 96.94 145.08 ;
      RECT 97.46 144.96 97.66 145.08 ;
      RECT 98.18 144.96 98.38 145.08 ;
      RECT 94.58 144.72 94.78 144.84 ;
      RECT 95.3 144.72 95.5 144.84 ;
      RECT 96.02 144.72 96.22 144.84 ;
      RECT 97.82 148.74 98.02 148.86 ;
      RECT 94.94 148.74 95.14 148.86 ;
      RECT 94.22 148.74 94.42 148.86 ;
      RECT 95.66 148.5 95.86 148.62 ;
      RECT 96.38 148.5 96.58 148.62 ;
      RECT 97.1 148.5 97.3 148.62 ;
      RECT 98.18 150 98.38 150.12 ;
      RECT 96.02 150 96.22 150.12 ;
      RECT 94.58 150 94.78 150.12 ;
      RECT 97.46 149.76 97.66 149.88 ;
      RECT 96.74 149.76 96.94 149.88 ;
      RECT 95.3 149.76 95.5 149.88 ;
      RECT 95.66 151.26 95.86 151.38 ;
      RECT 96.38 151.26 96.58 151.38 ;
      RECT 97.82 151.02 98.02 151.14 ;
      RECT 97.1 151.02 97.3 151.14 ;
      RECT 94.94 151.02 95.14 151.14 ;
      RECT 94.22 151.02 94.42 151.14 ;
      RECT 97.46 152.52 97.66 152.64 ;
      RECT 96.02 152.52 96.22 152.64 ;
      RECT 94.58 152.52 94.78 152.64 ;
      RECT 98.18 152.28 98.38 152.4 ;
      RECT 96.74 152.28 96.94 152.4 ;
      RECT 95.3 152.28 95.5 152.4 ;
      RECT 96.38 153.78 96.58 153.9 ;
      RECT 94.94 153.78 95.14 153.9 ;
      RECT 94.22 153.54 94.42 153.66 ;
      RECT 95.66 153.54 95.86 153.66 ;
      RECT 97.1 153.54 97.3 153.66 ;
      RECT 97.82 153.54 98.02 153.66 ;
      RECT 97.46 155.04 97.66 155.16 ;
      RECT 96.02 155.04 96.22 155.16 ;
      RECT 95.3 154.8 95.5 154.92 ;
      RECT 96.74 154.8 96.94 154.92 ;
      RECT 98.18 154.8 98.38 154.92 ;
      RECT 94.58 154.8 94.78 154.92 ;
      RECT 97.1 156.3 97.3 156.42 ;
      RECT 95.66 156.3 95.86 156.42 ;
      RECT 97.82 156.06 98.02 156.18 ;
      RECT 96.38 156.06 96.58 156.18 ;
      RECT 94.94 156.06 95.14 156.18 ;
      RECT 94.22 156.06 94.42 156.18 ;
      RECT 96.74 157.56 96.94 157.68 ;
      RECT 96.02 157.56 96.22 157.68 ;
      RECT 95.3 157.56 95.5 157.68 ;
      RECT 98.18 157.32 98.38 157.44 ;
      RECT 97.46 157.32 97.66 157.44 ;
      RECT 94.58 157.32 94.78 157.44 ;
      RECT 97.1 158.82 97.3 158.94 ;
      RECT 95.66 158.82 95.86 158.94 ;
      RECT 94.94 158.58 95.14 158.7 ;
      RECT 96.38 158.58 96.58 158.7 ;
      RECT 97.82 158.58 98.02 158.7 ;
      RECT 94.22 158.58 94.42 158.7 ;
      RECT 94.58 160.08 94.78 160.2 ;
      RECT 92.06 266.94 92.26 267.06 ;
      RECT 93.86 266.2885 94.06 266.4085 ;
      RECT 93.14 266.2885 93.34 266.4085 ;
      RECT 92.42 266.2885 92.62 266.4085 ;
      RECT 91.7 266.2885 91.9 266.4085 ;
      RECT 92.42 267.81 92.62 267.93 ;
      RECT 91.7 267.81 91.9 267.93 ;
      RECT 93.86 267.81 94.06 267.93 ;
      RECT 93.14 267.81 93.34 267.93 ;
      RECT 93.14 270.09 93.34 270.21 ;
      RECT 91.7 270.09 91.9 270.21 ;
      RECT 93.5 269.7 93.7 269.82 ;
      RECT 92.78 269.46 92.98 269.58 ;
      RECT 92.06 269.46 92.26 269.58 ;
      RECT 91.34 269.46 91.54 269.58 ;
      RECT 92.42 271.59 92.62 271.71 ;
      RECT 91.7 271.59 91.9 271.71 ;
      RECT 93.86 271.35 94.06 271.47 ;
      RECT 93.14 271.35 93.34 271.47 ;
      RECT 93.86 270.33 94.06 270.45 ;
      RECT 92.42 270.33 92.62 270.45 ;
      RECT 93.5 272.22 93.7 272.34 ;
      RECT 91.34 272.22 91.54 272.34 ;
      RECT 92.78 271.98 92.98 272.1 ;
      RECT 92.06 271.98 92.26 272.1 ;
      RECT 92.78 274.74 92.98 274.86 ;
      RECT 91.34 274.74 91.54 274.86 ;
      RECT 92.06 274.5 92.26 274.62 ;
      RECT 93.5 274.5 93.7 274.62 ;
      RECT 92.78 277.02 92.98 277.14 ;
      RECT 92.06 277.02 92.26 277.14 ;
      RECT 93.5 277.26 93.7 277.38 ;
      RECT 91.34 277.26 91.54 277.38 ;
      RECT 91.34 308.496 91.54 308.616 ;
      RECT 92.06 308.496 92.26 308.616 ;
      RECT 92.78 308.496 92.98 308.616 ;
      RECT 93.5 308.496 93.7 308.616 ;
      RECT 91.7 323.3835 91.9 323.5035 ;
      RECT 92.42 323.3835 92.62 323.5035 ;
      RECT 93.14 323.3835 93.34 323.5035 ;
      RECT 93.86 323.3835 94.06 323.5035 ;
      RECT 93.5 325.9425 93.7 326.0625 ;
      RECT 92.78 325.9425 92.98 326.0625 ;
      RECT 91.34 325.9425 91.54 326.0625 ;
      RECT 92.06 325.9425 92.26 326.0625 ;
      RECT 91.7 348.339 91.9 348.459 ;
      RECT 92.42 348.339 92.62 348.459 ;
      RECT 93.14 348.339 93.34 348.459 ;
      RECT 93.86 348.339 94.06 348.459 ;
      RECT 94.22 118.5 94.42 118.62 ;
      RECT 94.94 118.26 95.14 118.38 ;
      RECT 94.22 126.538 94.42 126.658 ;
      RECT 94.94 126.538 95.14 126.658 ;
      RECT 95.66 126.538 95.86 126.658 ;
      RECT 96.38 126.538 96.58 126.658 ;
      RECT 97.1 126.538 97.3 126.658 ;
      RECT 97.82 126.538 98.02 126.658 ;
      RECT 98.18 127.32 98.38 127.44 ;
      RECT 96.74 127.32 96.94 127.44 ;
      RECT 95.3 127.08 95.5 127.2 ;
      RECT 96.02 127.08 96.22 127.2 ;
      RECT 97.46 127.08 97.66 127.2 ;
      RECT 97.46 129.6 97.66 129.72 ;
      RECT 96.74 129.6 96.94 129.72 ;
      RECT 96.02 129.6 96.22 129.72 ;
      RECT 95.3 129.6 95.5 129.72 ;
      RECT 94.22 129.058 94.42 129.178 ;
      RECT 94.94 129.058 95.14 129.178 ;
      RECT 95.66 129.058 95.86 129.178 ;
      RECT 96.38 129.058 96.58 129.178 ;
      RECT 97.1 129.058 97.3 129.178 ;
      RECT 97.82 129.058 98.02 129.178 ;
      RECT 97.82 128.58 98.02 128.7 ;
      RECT 97.1 128.58 97.3 128.7 ;
      RECT 94.22 128.34 94.42 128.46 ;
      RECT 96.38 128.34 96.58 128.46 ;
      RECT 95.66 128.34 95.86 128.46 ;
      RECT 94.22 130.86 94.42 130.98 ;
      RECT 97.1 130.86 97.3 130.98 ;
      RECT 95.66 130.86 95.86 130.98 ;
      RECT 98.18 129.84 98.38 129.96 ;
      RECT 97.46 132.36 97.66 132.48 ;
      RECT 96.74 132.36 96.94 132.48 ;
      RECT 96.02 132.12 96.22 132.24 ;
      RECT 98.18 132.12 98.38 132.24 ;
      RECT 95.3 132.12 95.5 132.24 ;
      RECT 94.22 131.578 94.42 131.698 ;
      RECT 94.94 131.578 95.14 131.698 ;
      RECT 95.66 131.578 95.86 131.698 ;
      RECT 96.38 131.578 96.58 131.698 ;
      RECT 97.1 131.578 97.3 131.698 ;
      RECT 97.82 131.578 98.02 131.698 ;
      RECT 96.38 131.1 96.58 131.22 ;
      RECT 97.82 131.1 98.02 131.22 ;
      RECT 97.82 133.62 98.02 133.74 ;
      RECT 96.38 133.62 96.58 133.74 ;
      RECT 95.66 133.38 95.86 133.5 ;
      RECT 97.1 133.38 97.3 133.5 ;
      RECT 94.22 133.38 94.42 133.5 ;
      RECT 97.46 134.88 97.66 135 ;
      RECT 96.74 134.88 96.94 135 ;
      RECT 95.3 134.88 95.5 135 ;
      RECT 91.7 215.28 91.9 215.4 ;
      RECT 92.42 215.28 92.62 215.4 ;
      RECT 93.14 215.28 93.34 215.4 ;
      RECT 92.78 216.78 92.98 216.9 ;
      RECT 91.34 216.78 91.54 216.9 ;
      RECT 93.5 216.54 93.7 216.66 ;
      RECT 92.06 216.54 92.26 216.66 ;
      RECT 93.5 219.3 93.7 219.42 ;
      RECT 92.78 219.3 92.98 219.42 ;
      RECT 91.34 219.3 91.54 219.42 ;
      RECT 92.06 219.06 92.26 219.18 ;
      RECT 92.06 223.798 92.26 223.918 ;
      RECT 93.5 223.798 93.7 223.918 ;
      RECT 91.34 223.558 91.54 223.678 ;
      RECT 92.78 223.558 92.98 223.678 ;
      RECT 92.42 223.08 92.62 223.2 ;
      RECT 93.86 223.08 94.06 223.2 ;
      RECT 91.7 222.84 91.9 222.96 ;
      RECT 93.14 222.84 93.34 222.96 ;
      RECT 93.5 229.14 93.7 229.26 ;
      RECT 91.34 229.38 91.54 229.5 ;
      RECT 92.06 229.38 92.26 229.5 ;
      RECT 92.78 229.38 92.98 229.5 ;
      RECT 93.5 231.9 93.7 232.02 ;
      RECT 92.06 231.9 92.26 232.02 ;
      RECT 91.34 231.9 91.54 232.02 ;
      RECT 92.78 231.66 92.98 231.78 ;
      RECT 93.5 234.42 93.7 234.54 ;
      RECT 91.34 234.18 91.54 234.3 ;
      RECT 92.06 234.18 92.26 234.3 ;
      RECT 92.78 234.18 92.98 234.3 ;
      RECT 91.34 236.94 91.54 237.06 ;
      RECT 92.06 236.94 92.26 237.06 ;
      RECT 93.5 236.94 93.7 237.06 ;
      RECT 92.78 236.7 92.98 236.82 ;
      RECT 93.5 239.46 93.7 239.58 ;
      RECT 92.06 239.46 92.26 239.58 ;
      RECT 91.34 239.46 91.54 239.58 ;
      RECT 92.78 239.22 92.98 239.34 ;
      RECT 91.34 241.98 91.54 242.1 ;
      RECT 92.06 241.98 92.26 242.1 ;
      RECT 93.5 241.98 93.7 242.1 ;
      RECT 92.78 241.74 92.98 241.86 ;
      RECT 91.34 244.26 91.54 244.38 ;
      RECT 92.06 244.5 92.26 244.62 ;
      RECT 92.78 244.5 92.98 244.62 ;
      RECT 93.5 244.5 93.7 244.62 ;
      RECT 92.78 247.02 92.98 247.14 ;
      RECT 92.06 247.02 92.26 247.14 ;
      RECT 93.5 246.78 93.7 246.9 ;
      RECT 91.34 246.78 91.54 246.9 ;
      RECT 93.5 249.54 93.7 249.66 ;
      RECT 92.78 249.54 92.98 249.66 ;
      RECT 92.06 249.54 92.26 249.66 ;
      RECT 91.34 249.3 91.54 249.42 ;
      RECT 92.78 252.06 92.98 252.18 ;
      RECT 91.34 252.06 91.54 252.18 ;
      RECT 93.5 251.82 93.7 251.94 ;
      RECT 92.06 251.82 92.26 251.94 ;
      RECT 92.78 254.58 92.98 254.7 ;
      RECT 93.5 254.34 93.7 254.46 ;
      RECT 92.06 254.34 92.26 254.46 ;
      RECT 91.34 254.34 91.54 254.46 ;
      RECT 92.78 257.1 92.98 257.22 ;
      RECT 91.34 257.1 91.54 257.22 ;
      RECT 93.5 256.86 93.7 256.98 ;
      RECT 92.06 256.86 92.26 256.98 ;
      RECT 93.86 258.99 94.06 259.11 ;
      RECT 92.42 258.99 92.62 259.11 ;
      RECT 93.14 258.75 93.34 258.87 ;
      RECT 91.7 258.75 91.9 258.87 ;
      RECT 93.86 260.25 94.06 260.37 ;
      RECT 92.42 260.25 92.62 260.37 ;
      RECT 93.14 260.01 93.34 260.13 ;
      RECT 91.7 260.01 91.9 260.13 ;
      RECT 93.5 259.62 93.7 259.74 ;
      RECT 91.34 259.62 91.54 259.74 ;
      RECT 92.78 259.38 92.98 259.5 ;
      RECT 92.06 259.38 92.26 259.5 ;
      RECT 92.78 261.9 92.98 262.02 ;
      RECT 92.06 261.9 92.26 262.02 ;
      RECT 91.34 261.9 91.54 262.02 ;
      RECT 93.86 261.51 94.06 261.63 ;
      RECT 91.7 261.51 91.9 261.63 ;
      RECT 93.14 261.27 93.34 261.39 ;
      RECT 92.42 261.27 92.62 261.39 ;
      RECT 92.42 262.77 92.62 262.89 ;
      RECT 93.86 262.53 94.06 262.65 ;
      RECT 93.14 262.53 93.34 262.65 ;
      RECT 91.7 262.53 91.9 262.65 ;
      RECT 93.5 262.14 93.7 262.26 ;
      RECT 93.5 264.66 93.7 264.78 ;
      RECT 92.06 264.66 92.26 264.78 ;
      RECT 91.34 264.66 91.54 264.78 ;
      RECT 92.78 264.42 92.98 264.54 ;
      RECT 93.86 264.03 94.06 264.15 ;
      RECT 92.42 264.03 92.62 264.15 ;
      RECT 91.7 264.03 91.9 264.15 ;
      RECT 93.14 264.03 93.34 264.15 ;
      RECT 93.5 267.18 93.7 267.3 ;
      RECT 91.34 267.18 91.54 267.3 ;
      RECT 92.78 266.94 92.98 267.06 ;
      RECT 91.7 182.52 91.9 182.64 ;
      RECT 93.5 184.02 93.7 184.14 ;
      RECT 92.06 184.02 92.26 184.14 ;
      RECT 91.34 184.02 91.54 184.14 ;
      RECT 92.78 183.78 92.98 183.9 ;
      RECT 93.86 185.28 94.06 185.4 ;
      RECT 91.7 185.28 91.9 185.4 ;
      RECT 93.14 185.04 93.34 185.16 ;
      RECT 92.42 185.04 92.62 185.16 ;
      RECT 92.06 186.54 92.26 186.66 ;
      RECT 93.5 186.54 93.7 186.66 ;
      RECT 91.34 186.3 91.54 186.42 ;
      RECT 92.78 186.3 92.98 186.42 ;
      RECT 93.14 187.8 93.34 187.92 ;
      RECT 92.42 187.8 92.62 187.92 ;
      RECT 91.7 187.8 91.9 187.92 ;
      RECT 93.86 187.56 94.06 187.68 ;
      RECT 91.34 189.06 91.54 189.18 ;
      RECT 93.5 188.82 93.7 188.94 ;
      RECT 92.78 188.82 92.98 188.94 ;
      RECT 92.06 188.82 92.26 188.94 ;
      RECT 93.14 190.32 93.34 190.44 ;
      RECT 91.7 190.32 91.9 190.44 ;
      RECT 92.42 190.08 92.62 190.2 ;
      RECT 93.86 190.08 94.06 190.2 ;
      RECT 91.34 191.58 91.54 191.7 ;
      RECT 93.5 191.34 93.7 191.46 ;
      RECT 92.78 191.34 92.98 191.46 ;
      RECT 92.06 191.34 92.26 191.46 ;
      RECT 92.42 192.84 92.62 192.96 ;
      RECT 91.7 192.84 91.9 192.96 ;
      RECT 93.86 192.84 94.06 192.96 ;
      RECT 93.14 192.6 93.34 192.72 ;
      RECT 93.5 194.1 93.7 194.22 ;
      RECT 92.78 193.86 92.98 193.98 ;
      RECT 92.06 193.86 92.26 193.98 ;
      RECT 91.34 193.86 91.54 193.98 ;
      RECT 92.42 195.12 92.62 195.24 ;
      RECT 91.7 195.12 91.9 195.24 ;
      RECT 93.86 195.36 94.06 195.48 ;
      RECT 93.14 195.36 93.34 195.48 ;
      RECT 93.5 196.38 93.7 196.5 ;
      RECT 92.78 196.38 92.98 196.5 ;
      RECT 91.34 196.38 91.54 196.5 ;
      RECT 92.06 196.62 92.26 196.74 ;
      RECT 91.7 197.64 91.9 197.76 ;
      RECT 93.86 197.64 94.06 197.76 ;
      RECT 93.14 197.88 93.34 198 ;
      RECT 92.42 197.88 92.62 198 ;
      RECT 91.34 198.9 91.54 199.02 ;
      RECT 93.5 199.14 93.7 199.26 ;
      RECT 92.78 199.14 92.98 199.26 ;
      RECT 92.06 199.14 92.26 199.26 ;
      RECT 92.42 200.16 92.62 200.28 ;
      RECT 93.86 200.16 94.06 200.28 ;
      RECT 91.7 200.4 91.9 200.52 ;
      RECT 93.14 200.4 93.34 200.52 ;
      RECT 93.5 201.66 93.7 201.78 ;
      RECT 92.78 201.66 92.98 201.78 ;
      RECT 92.06 201.66 92.26 201.78 ;
      RECT 91.34 201.66 91.54 201.78 ;
      RECT 93.86 202.68 94.06 202.8 ;
      RECT 93.14 202.68 93.34 202.8 ;
      RECT 92.42 202.68 92.62 202.8 ;
      RECT 91.7 202.68 91.9 202.8 ;
      RECT 91.34 203.94 91.54 204.06 ;
      RECT 92.06 203.94 92.26 204.06 ;
      RECT 92.78 203.94 92.98 204.06 ;
      RECT 93.5 203.94 93.7 204.06 ;
      RECT 93.14 205.2 93.34 205.32 ;
      RECT 93.86 205.44 94.06 205.56 ;
      RECT 92.42 205.44 92.62 205.56 ;
      RECT 91.7 205.44 91.9 205.56 ;
      RECT 91.34 206.46 91.54 206.58 ;
      RECT 92.06 206.46 92.26 206.58 ;
      RECT 92.78 206.7 92.98 206.82 ;
      RECT 93.5 206.7 93.7 206.82 ;
      RECT 92.42 207.72 92.62 207.84 ;
      RECT 93.14 207.96 93.34 208.08 ;
      RECT 93.86 207.96 94.06 208.08 ;
      RECT 91.7 207.96 91.9 208.08 ;
      RECT 93.5 208.98 93.7 209.1 ;
      RECT 91.34 209.22 91.54 209.34 ;
      RECT 92.06 209.22 92.26 209.34 ;
      RECT 92.78 209.22 92.98 209.34 ;
      RECT 93.5 211.5 93.7 211.62 ;
      RECT 91.34 211.5 91.54 211.62 ;
      RECT 93.14 210.48 93.34 210.6 ;
      RECT 91.7 210.24 91.9 210.36 ;
      RECT 92.42 210.24 92.62 210.36 ;
      RECT 93.86 210.24 94.06 210.36 ;
      RECT 91.7 212.76 91.9 212.88 ;
      RECT 93.14 212.76 93.34 212.88 ;
      RECT 93.86 212.76 94.06 212.88 ;
      RECT 92.78 211.74 92.98 211.86 ;
      RECT 92.06 211.74 92.26 211.86 ;
      RECT 92.78 214.26 92.98 214.38 ;
      RECT 92.06 214.26 92.26 214.38 ;
      RECT 91.34 214.26 91.54 214.38 ;
      RECT 93.5 214.02 93.7 214.14 ;
      RECT 92.42 213 92.62 213.12 ;
      RECT 93.86 215.52 94.06 215.64 ;
      RECT 93.5 151.26 93.7 151.38 ;
      RECT 92.78 151.02 92.98 151.14 ;
      RECT 92.06 151.02 92.26 151.14 ;
      RECT 93.14 152.52 93.34 152.64 ;
      RECT 91.7 152.52 91.9 152.64 ;
      RECT 93.86 152.28 94.06 152.4 ;
      RECT 92.42 152.28 92.62 152.4 ;
      RECT 92.06 153.78 92.26 153.9 ;
      RECT 92.78 153.78 92.98 153.9 ;
      RECT 91.34 153.54 91.54 153.66 ;
      RECT 93.5 153.54 93.7 153.66 ;
      RECT 92.42 155.04 92.62 155.16 ;
      RECT 91.7 154.8 91.9 154.92 ;
      RECT 93.14 154.8 93.34 154.92 ;
      RECT 93.86 154.8 94.06 154.92 ;
      RECT 93.5 156.3 93.7 156.42 ;
      RECT 91.34 156.3 91.54 156.42 ;
      RECT 92.78 156.06 92.98 156.18 ;
      RECT 92.06 156.06 92.26 156.18 ;
      RECT 93.14 157.56 93.34 157.68 ;
      RECT 92.42 157.56 92.62 157.68 ;
      RECT 93.86 157.32 94.06 157.44 ;
      RECT 91.7 157.32 91.9 157.44 ;
      RECT 93.5 158.82 93.7 158.94 ;
      RECT 91.34 158.82 91.54 158.94 ;
      RECT 92.78 158.58 92.98 158.7 ;
      RECT 92.06 158.58 92.26 158.7 ;
      RECT 92.42 160.08 92.62 160.2 ;
      RECT 93.14 160.08 93.34 160.2 ;
      RECT 93.86 159.84 94.06 159.96 ;
      RECT 91.7 159.84 91.9 159.96 ;
      RECT 91.34 161.1 91.54 161.22 ;
      RECT 92.06 161.1 92.26 161.22 ;
      RECT 92.78 161.1 92.98 161.22 ;
      RECT 93.5 161.1 93.7 161.22 ;
      RECT 92.78 163.62 92.98 163.74 ;
      RECT 93.86 162.6 94.06 162.72 ;
      RECT 93.14 162.6 93.34 162.72 ;
      RECT 92.42 162.6 92.62 162.72 ;
      RECT 91.7 162.6 91.9 162.72 ;
      RECT 92.42 165.12 92.62 165.24 ;
      RECT 91.7 165.12 91.9 165.24 ;
      RECT 93.86 164.88 94.06 165 ;
      RECT 93.14 164.88 93.34 165 ;
      RECT 93.5 163.86 93.7 163.98 ;
      RECT 92.06 163.86 92.26 163.98 ;
      RECT 91.34 163.86 91.54 163.98 ;
      RECT 92.06 166.38 92.26 166.5 ;
      RECT 92.78 166.38 92.98 166.5 ;
      RECT 93.5 166.14 93.7 166.26 ;
      RECT 91.34 166.14 91.54 166.26 ;
      RECT 93.14 167.64 93.34 167.76 ;
      RECT 91.7 167.64 91.9 167.76 ;
      RECT 92.42 167.4 92.62 167.52 ;
      RECT 93.86 167.4 94.06 167.52 ;
      RECT 92.78 168.9 92.98 169.02 ;
      RECT 92.06 168.9 92.26 169.02 ;
      RECT 91.34 168.66 91.54 168.78 ;
      RECT 93.5 168.66 93.7 168.78 ;
      RECT 93.86 170.16 94.06 170.28 ;
      RECT 92.42 170.16 92.62 170.28 ;
      RECT 93.14 169.92 93.34 170.04 ;
      RECT 91.7 169.92 91.9 170.04 ;
      RECT 92.06 171.42 92.26 171.54 ;
      RECT 93.5 171.18 93.7 171.3 ;
      RECT 92.78 171.18 92.98 171.3 ;
      RECT 91.34 171.18 91.54 171.3 ;
      RECT 91.7 172.68 91.9 172.8 ;
      RECT 92.42 172.44 92.62 172.56 ;
      RECT 93.14 172.44 93.34 172.56 ;
      RECT 93.86 172.44 94.06 172.56 ;
      RECT 92.78 173.94 92.98 174.06 ;
      RECT 92.06 173.94 92.26 174.06 ;
      RECT 91.34 173.94 91.54 174.06 ;
      RECT 93.5 173.7 93.7 173.82 ;
      RECT 93.14 175.2 93.34 175.32 ;
      RECT 92.42 175.2 92.62 175.32 ;
      RECT 91.7 175.2 91.9 175.32 ;
      RECT 93.86 174.96 94.06 175.08 ;
      RECT 93.5 176.46 93.7 176.58 ;
      RECT 92.06 176.46 92.26 176.58 ;
      RECT 92.78 176.22 92.98 176.34 ;
      RECT 91.34 176.22 91.54 176.34 ;
      RECT 93.5 178.74 93.7 178.86 ;
      RECT 91.34 178.74 91.54 178.86 ;
      RECT 93.86 177.72 94.06 177.84 ;
      RECT 91.7 177.72 91.9 177.84 ;
      RECT 93.14 177.48 93.34 177.6 ;
      RECT 92.42 177.48 92.62 177.6 ;
      RECT 93.86 180 94.06 180.12 ;
      RECT 92.42 180 92.62 180.12 ;
      RECT 92.78 178.98 92.98 179.1 ;
      RECT 92.06 178.98 92.26 179.1 ;
      RECT 92.78 181.5 92.98 181.62 ;
      RECT 91.34 181.5 91.54 181.62 ;
      RECT 93.5 181.26 93.7 181.38 ;
      RECT 92.06 181.26 92.26 181.38 ;
      RECT 93.14 180.24 93.34 180.36 ;
      RECT 91.7 180.24 91.9 180.36 ;
      RECT 93.86 182.76 94.06 182.88 ;
      RECT 92.42 182.76 92.62 182.88 ;
      RECT 93.14 182.52 93.34 182.64 ;
      RECT 86.66 270.33 86.86 270.45 ;
      RECT 85.94 270.33 86.14 270.45 ;
      RECT 85.22 270.33 85.42 270.45 ;
      RECT 84.5 270.33 84.7 270.45 ;
      RECT 83.06 270.33 83.26 270.45 ;
      RECT 83.78 275.76 83.98 275.88 ;
      RECT 83.42 274.74 83.62 274.86 ;
      RECT 82.7 274.74 82.9 274.86 ;
      RECT 81.98 274.74 82.18 274.86 ;
      RECT 84.14 274.5 84.34 274.62 ;
      RECT 83.78 273.48 83.98 273.6 ;
      RECT 82.34 273.24 82.54 273.36 ;
      RECT 83.78 278.28 83.98 278.4 ;
      RECT 82.34 278.28 82.54 278.4 ;
      RECT 84.14 277.26 84.34 277.38 ;
      RECT 82.7 277.26 82.9 277.38 ;
      RECT 83.42 277.02 83.62 277.14 ;
      RECT 81.98 277.02 82.18 277.14 ;
      RECT 82.34 276 82.54 276.12 ;
      RECT 82.7 308.496 82.9 308.616 ;
      RECT 81.98 308.496 82.18 308.616 ;
      RECT 84.14 308.496 84.34 308.616 ;
      RECT 83.42 308.496 83.62 308.616 ;
      RECT 87.38 323.3835 87.58 323.5035 ;
      RECT 86.66 323.3835 86.86 323.5035 ;
      RECT 85.94 323.3835 86.14 323.5035 ;
      RECT 85.22 323.3835 85.42 323.5035 ;
      RECT 84.5 323.3835 84.7 323.5035 ;
      RECT 83.06 323.3835 83.26 323.5035 ;
      RECT 84.14 325.9425 84.34 326.0625 ;
      RECT 83.42 325.9425 83.62 326.0625 ;
      RECT 82.7 325.9425 82.9 326.0625 ;
      RECT 81.98 325.9425 82.18 326.0625 ;
      RECT 85.22 348.339 85.42 348.459 ;
      RECT 84.5 348.339 84.7 348.459 ;
      RECT 83.06 348.339 83.26 348.459 ;
      RECT 87.38 348.339 87.58 348.459 ;
      RECT 86.66 348.339 86.86 348.459 ;
      RECT 85.94 348.339 86.14 348.459 ;
      RECT 92.78 118.5 92.98 118.62 ;
      RECT 91.34 118.5 91.54 118.62 ;
      RECT 93.5 118.26 93.7 118.38 ;
      RECT 92.06 118.26 92.26 118.38 ;
      RECT 93.5 126.538 93.7 126.658 ;
      RECT 93.5 129.058 93.7 129.178 ;
      RECT 93.5 128.34 93.7 128.46 ;
      RECT 93.5 130.86 93.7 130.98 ;
      RECT 93.5 131.578 93.7 131.698 ;
      RECT 91.34 133.62 91.54 133.74 ;
      RECT 92.06 133.38 92.26 133.5 ;
      RECT 93.5 133.38 93.7 133.5 ;
      RECT 91.7 134.88 91.9 135 ;
      RECT 92.42 134.64 92.62 134.76 ;
      RECT 91.34 134.098 91.54 134.218 ;
      RECT 92.06 134.098 92.26 134.218 ;
      RECT 92.78 134.098 92.98 134.218 ;
      RECT 93.5 134.098 93.7 134.218 ;
      RECT 91.34 136.14 91.54 136.26 ;
      RECT 92.06 135.9 92.26 136.02 ;
      RECT 93.5 135.9 93.7 136.02 ;
      RECT 91.7 137.4 91.9 137.52 ;
      RECT 92.42 137.16 92.62 137.28 ;
      RECT 91.34 136.858 91.54 136.978 ;
      RECT 92.78 136.858 92.98 136.978 ;
      RECT 92.06 136.618 92.26 136.738 ;
      RECT 93.5 136.618 93.7 136.738 ;
      RECT 92.06 139.138 92.26 139.258 ;
      RECT 93.5 139.138 93.7 139.258 ;
      RECT 93.5 138.66 93.7 138.78 ;
      RECT 91.34 138.66 91.54 138.78 ;
      RECT 92.06 138.42 92.26 138.54 ;
      RECT 91.7 139.92 91.9 140.04 ;
      RECT 92.42 139.68 92.62 139.8 ;
      RECT 91.34 139.378 91.54 139.498 ;
      RECT 92.78 139.378 92.98 139.498 ;
      RECT 91.34 141.18 91.54 141.3 ;
      RECT 92.06 140.94 92.26 141.06 ;
      RECT 93.5 140.94 93.7 141.06 ;
      RECT 93.86 142.44 94.06 142.56 ;
      RECT 92.42 142.44 92.62 142.56 ;
      RECT 93.14 142.2 93.34 142.32 ;
      RECT 91.7 142.2 91.9 142.32 ;
      RECT 93.5 143.46 93.7 143.58 ;
      RECT 92.06 143.46 92.26 143.58 ;
      RECT 91.34 143.7 91.54 143.82 ;
      RECT 91.34 145.98 91.54 146.1 ;
      RECT 92.06 145.98 92.26 146.1 ;
      RECT 92.78 145.98 92.98 146.1 ;
      RECT 93.5 145.98 93.7 146.1 ;
      RECT 91.7 144.96 91.9 145.08 ;
      RECT 93.86 144.96 94.06 145.08 ;
      RECT 92.42 144.72 92.62 144.84 ;
      RECT 93.14 144.72 93.34 144.84 ;
      RECT 92.78 148.74 92.98 148.86 ;
      RECT 91.34 148.74 91.54 148.86 ;
      RECT 92.06 148.5 92.26 148.62 ;
      RECT 93.5 148.5 93.7 148.62 ;
      RECT 92.42 150 92.62 150.12 ;
      RECT 91.7 150 91.9 150.12 ;
      RECT 93.86 150 94.06 150.12 ;
      RECT 93.14 149.76 93.34 149.88 ;
      RECT 91.34 151.26 91.54 151.38 ;
      RECT 81.98 249.3 82.18 249.42 ;
      RECT 83.78 253.32 83.98 253.44 ;
      RECT 82.34 253.32 82.54 253.44 ;
      RECT 81.98 252.06 82.18 252.18 ;
      RECT 83.42 252.06 83.62 252.18 ;
      RECT 84.14 251.82 84.34 251.94 ;
      RECT 82.7 251.82 82.9 251.94 ;
      RECT 82.34 255.84 82.54 255.96 ;
      RECT 83.78 255.6 83.98 255.72 ;
      RECT 82.7 254.58 82.9 254.7 ;
      RECT 81.98 254.58 82.18 254.7 ;
      RECT 84.14 254.34 84.34 254.46 ;
      RECT 83.42 254.34 83.62 254.46 ;
      RECT 84.14 259.38 84.34 259.5 ;
      RECT 87.38 258.99 87.58 259.11 ;
      RECT 85.94 258.99 86.14 259.11 ;
      RECT 83.06 258.99 83.26 259.11 ;
      RECT 86.66 258.75 86.86 258.87 ;
      RECT 85.22 258.75 85.42 258.87 ;
      RECT 84.5 258.75 84.7 258.87 ;
      RECT 82.34 258.36 82.54 258.48 ;
      RECT 83.78 258.12 83.98 258.24 ;
      RECT 84.14 257.1 84.34 257.22 ;
      RECT 81.98 257.1 82.18 257.22 ;
      RECT 83.42 256.86 83.62 256.98 ;
      RECT 82.7 256.86 82.9 256.98 ;
      RECT 84.14 261.9 84.34 262.02 ;
      RECT 83.42 261.9 83.62 262.02 ;
      RECT 87.38 261.51 87.58 261.63 ;
      RECT 85.22 261.51 85.42 261.63 ;
      RECT 83.06 261.51 83.26 261.63 ;
      RECT 86.66 261.27 86.86 261.39 ;
      RECT 85.94 261.27 86.14 261.39 ;
      RECT 84.5 261.27 84.7 261.39 ;
      RECT 82.34 260.88 82.54 261 ;
      RECT 83.78 260.64 83.98 260.76 ;
      RECT 85.22 260.25 85.42 260.37 ;
      RECT 85.94 260.25 86.14 260.37 ;
      RECT 87.38 260.25 87.58 260.37 ;
      RECT 84.5 260.25 84.7 260.37 ;
      RECT 86.66 260.01 86.86 260.13 ;
      RECT 83.06 260.01 83.26 260.13 ;
      RECT 83.42 259.62 83.62 259.74 ;
      RECT 82.7 259.62 82.9 259.74 ;
      RECT 81.98 259.62 82.18 259.74 ;
      RECT 82.7 264.66 82.9 264.78 ;
      RECT 83.42 264.66 83.62 264.78 ;
      RECT 84.14 264.42 84.34 264.54 ;
      RECT 81.98 264.42 82.18 264.54 ;
      RECT 85.22 264.03 85.42 264.15 ;
      RECT 83.06 264.03 83.26 264.15 ;
      RECT 86.66 264.03 86.86 264.15 ;
      RECT 87.38 263.79 87.58 263.91 ;
      RECT 85.94 263.79 86.14 263.91 ;
      RECT 84.5 263.79 84.7 263.91 ;
      RECT 83.78 263.4 83.98 263.52 ;
      RECT 82.34 263.16 82.54 263.28 ;
      RECT 87.38 262.77 87.58 262.89 ;
      RECT 85.22 262.77 85.42 262.89 ;
      RECT 84.5 262.77 84.7 262.89 ;
      RECT 83.06 262.77 83.26 262.89 ;
      RECT 86.66 262.53 86.86 262.65 ;
      RECT 85.94 262.53 86.14 262.65 ;
      RECT 82.7 262.14 82.9 262.26 ;
      RECT 81.98 262.14 82.18 262.26 ;
      RECT 84.14 267.18 84.34 267.3 ;
      RECT 83.42 267.18 83.62 267.3 ;
      RECT 81.98 267.18 82.18 267.3 ;
      RECT 82.7 266.94 82.9 267.06 ;
      RECT 87.38 266.2885 87.58 266.4085 ;
      RECT 86.66 266.2885 86.86 266.4085 ;
      RECT 85.94 266.2885 86.14 266.4085 ;
      RECT 85.22 266.2885 85.42 266.4085 ;
      RECT 84.5 266.2885 84.7 266.4085 ;
      RECT 83.06 266.2885 83.26 266.4085 ;
      RECT 82.34 265.92 82.54 266.04 ;
      RECT 83.78 265.92 83.98 266.04 ;
      RECT 87.38 270.09 87.58 270.21 ;
      RECT 84.14 269.7 84.34 269.82 ;
      RECT 83.42 269.7 83.62 269.82 ;
      RECT 81.98 269.7 82.18 269.82 ;
      RECT 82.7 269.46 82.9 269.58 ;
      RECT 82.34 268.44 82.54 268.56 ;
      RECT 83.78 268.2 83.98 268.32 ;
      RECT 87.38 267.81 87.58 267.93 ;
      RECT 86.66 267.81 86.86 267.93 ;
      RECT 85.94 267.81 86.14 267.93 ;
      RECT 85.22 267.81 85.42 267.93 ;
      RECT 84.5 267.81 84.7 267.93 ;
      RECT 83.06 267.81 83.26 267.93 ;
      RECT 82.7 272.22 82.9 272.34 ;
      RECT 81.98 272.22 82.18 272.34 ;
      RECT 84.14 271.98 84.34 272.1 ;
      RECT 83.42 271.98 83.62 272.1 ;
      RECT 87.38 271.59 87.58 271.71 ;
      RECT 86.66 271.59 86.86 271.71 ;
      RECT 85.22 271.59 85.42 271.71 ;
      RECT 83.06 271.59 83.26 271.71 ;
      RECT 85.94 271.35 86.14 271.47 ;
      RECT 84.5 271.35 84.7 271.47 ;
      RECT 83.78 270.96 83.98 271.08 ;
      RECT 82.34 270.96 82.54 271.08 ;
      RECT 85.94 205.2 86.14 205.32 ;
      RECT 84.5 210.24 84.7 210.36 ;
      RECT 83.42 209.22 83.62 209.34 ;
      RECT 82.7 209.22 82.9 209.34 ;
      RECT 81.98 208.98 82.18 209.1 ;
      RECT 84.14 208.98 84.34 209.1 ;
      RECT 82.34 208.502 82.54 208.622 ;
      RECT 83.78 208.262 83.98 208.382 ;
      RECT 87.38 207.96 87.58 208.08 ;
      RECT 85.94 207.96 86.14 208.08 ;
      RECT 84.5 207.96 84.7 208.08 ;
      RECT 83.06 207.72 83.26 207.84 ;
      RECT 85.22 207.72 85.42 207.84 ;
      RECT 86.66 207.72 86.86 207.84 ;
      RECT 84.5 212.76 84.7 212.88 ;
      RECT 86.66 212.76 86.86 212.88 ;
      RECT 82.7 211.74 82.9 211.86 ;
      RECT 81.98 211.74 82.18 211.86 ;
      RECT 84.14 211.5 84.34 211.62 ;
      RECT 83.42 211.5 83.62 211.62 ;
      RECT 82.34 211.198 82.54 211.318 ;
      RECT 83.78 210.958 83.98 211.078 ;
      RECT 83.06 210.48 83.26 210.6 ;
      RECT 85.22 210.48 85.42 210.6 ;
      RECT 85.94 210.48 86.14 210.6 ;
      RECT 86.66 210.48 86.86 210.6 ;
      RECT 87.38 210.48 87.58 210.6 ;
      RECT 87.38 215.52 87.58 215.64 ;
      RECT 86.66 215.52 86.86 215.64 ;
      RECT 85.94 215.52 86.14 215.64 ;
      RECT 84.5 215.52 84.7 215.64 ;
      RECT 83.06 215.28 83.26 215.4 ;
      RECT 85.22 215.28 85.42 215.4 ;
      RECT 82.7 214.26 82.9 214.38 ;
      RECT 81.98 214.26 82.18 214.38 ;
      RECT 84.14 214.26 84.34 214.38 ;
      RECT 83.42 214.02 83.62 214.14 ;
      RECT 83.06 213 83.26 213.12 ;
      RECT 85.22 213 85.42 213.12 ;
      RECT 85.94 213 86.14 213.12 ;
      RECT 87.38 213 87.58 213.12 ;
      RECT 82.7 216.78 82.9 216.9 ;
      RECT 84.14 216.54 84.34 216.66 ;
      RECT 83.42 216.54 83.62 216.66 ;
      RECT 81.98 216.54 82.18 216.66 ;
      RECT 84.14 219.3 84.34 219.42 ;
      RECT 82.7 219.3 82.9 219.42 ;
      RECT 81.98 219.06 82.18 219.18 ;
      RECT 83.42 219.06 83.62 219.18 ;
      RECT 81.98 223.798 82.18 223.918 ;
      RECT 83.42 223.798 83.62 223.918 ;
      RECT 82.7 223.558 82.9 223.678 ;
      RECT 84.14 223.558 84.34 223.678 ;
      RECT 83.06 223.08 83.26 223.2 ;
      RECT 84.5 223.08 84.7 223.2 ;
      RECT 87.38 223.08 87.58 223.2 ;
      RECT 85.22 222.84 85.42 222.96 ;
      RECT 85.94 222.84 86.14 222.96 ;
      RECT 86.66 222.84 86.86 222.96 ;
      RECT 83.78 222.362 83.98 222.482 ;
      RECT 82.34 222.122 82.54 222.242 ;
      RECT 85.58 224.8315 85.78 224.9515 ;
      RECT 87.02 224.8315 87.22 224.9515 ;
      RECT 86.3 224.5915 86.5 224.7115 ;
      RECT 87.74 224.5915 87.94 224.7115 ;
      RECT 81.98 229.14 82.18 229.26 ;
      RECT 84.14 229.14 84.34 229.26 ;
      RECT 83.42 231.9 83.62 232.02 ;
      RECT 82.7 231.9 82.9 232.02 ;
      RECT 84.14 231.66 84.34 231.78 ;
      RECT 81.98 231.66 82.18 231.78 ;
      RECT 82.7 229.38 82.9 229.5 ;
      RECT 83.42 229.38 83.62 229.5 ;
      RECT 84.14 234.42 84.34 234.54 ;
      RECT 81.98 234.42 82.18 234.54 ;
      RECT 82.7 234.18 82.9 234.3 ;
      RECT 83.42 234.18 83.62 234.3 ;
      RECT 82.7 236.94 82.9 237.06 ;
      RECT 83.42 236.94 83.62 237.06 ;
      RECT 81.98 236.7 82.18 236.82 ;
      RECT 84.14 236.7 84.34 236.82 ;
      RECT 84.14 239.46 84.34 239.58 ;
      RECT 82.7 239.46 82.9 239.58 ;
      RECT 83.42 239.22 83.62 239.34 ;
      RECT 81.98 239.22 82.18 239.34 ;
      RECT 82.7 241.98 82.9 242.1 ;
      RECT 81.98 241.74 82.18 241.86 ;
      RECT 83.42 241.74 83.62 241.86 ;
      RECT 84.14 241.74 84.34 241.86 ;
      RECT 81.98 244.5 82.18 244.62 ;
      RECT 84.14 244.5 84.34 244.62 ;
      RECT 83.42 244.26 83.62 244.38 ;
      RECT 82.7 244.26 82.9 244.38 ;
      RECT 83.42 247.02 83.62 247.14 ;
      RECT 82.7 247.02 82.9 247.14 ;
      RECT 84.14 246.78 84.34 246.9 ;
      RECT 81.98 246.78 82.18 246.9 ;
      RECT 83.78 250.56 83.98 250.68 ;
      RECT 82.34 250.56 82.54 250.68 ;
      RECT 83.42 249.54 83.62 249.66 ;
      RECT 82.7 249.54 82.9 249.66 ;
      RECT 84.14 249.3 84.34 249.42 ;
      RECT 85.58 187.082 85.78 187.202 ;
      RECT 87.02 187.082 87.22 187.202 ;
      RECT 84.86 186.842 85.06 186.962 ;
      RECT 86.3 186.842 86.5 186.962 ;
      RECT 87.74 186.842 87.94 186.962 ;
      RECT 83.42 186.54 83.62 186.66 ;
      RECT 81.98 186.3 82.18 186.42 ;
      RECT 82.7 186.3 82.9 186.42 ;
      RECT 84.14 186.3 84.34 186.42 ;
      RECT 85.58 185.822 85.78 185.942 ;
      RECT 87.74 185.822 87.94 185.942 ;
      RECT 82.34 190.862 82.54 190.982 ;
      RECT 83.78 190.622 83.98 190.742 ;
      RECT 86.66 190.32 86.86 190.44 ;
      RECT 85.94 190.32 86.14 190.44 ;
      RECT 83.06 190.32 83.26 190.44 ;
      RECT 84.5 190.08 84.7 190.2 ;
      RECT 85.22 190.08 85.42 190.2 ;
      RECT 87.38 190.08 87.58 190.2 ;
      RECT 83.42 189.06 83.62 189.18 ;
      RECT 84.14 188.82 84.34 188.94 ;
      RECT 82.7 188.82 82.9 188.94 ;
      RECT 81.98 188.82 82.18 188.94 ;
      RECT 84.14 193.86 84.34 193.98 ;
      RECT 83.42 193.86 83.62 193.98 ;
      RECT 82.34 193.382 82.54 193.502 ;
      RECT 83.78 193.142 83.98 193.262 ;
      RECT 86.66 192.84 86.86 192.96 ;
      RECT 85.94 192.84 86.14 192.96 ;
      RECT 83.06 192.84 83.26 192.96 ;
      RECT 84.5 192.6 84.7 192.72 ;
      RECT 85.22 192.6 85.42 192.72 ;
      RECT 87.38 192.6 87.58 192.72 ;
      RECT 82.34 191.882 82.54 192.002 ;
      RECT 83.78 191.882 83.98 192.002 ;
      RECT 84.14 191.58 84.34 191.7 ;
      RECT 83.42 191.58 83.62 191.7 ;
      RECT 81.98 191.58 82.18 191.7 ;
      RECT 82.7 191.34 82.9 191.46 ;
      RECT 83.78 194.402 83.98 194.522 ;
      RECT 82.34 194.402 82.54 194.522 ;
      RECT 82.7 194.1 82.9 194.22 ;
      RECT 81.98 194.1 82.18 194.22 ;
      RECT 83.42 196.38 83.62 196.5 ;
      RECT 84.14 196.38 84.34 196.5 ;
      RECT 83.78 195.662 83.98 195.782 ;
      RECT 82.34 195.662 82.54 195.782 ;
      RECT 83.06 195.36 83.26 195.48 ;
      RECT 84.5 195.36 84.7 195.48 ;
      RECT 87.38 195.36 87.58 195.48 ;
      RECT 85.22 195.12 85.42 195.24 ;
      RECT 85.94 195.12 86.14 195.24 ;
      RECT 86.66 195.12 86.86 195.24 ;
      RECT 81.98 199.14 82.18 199.26 ;
      RECT 84.14 198.9 84.34 199.02 ;
      RECT 83.42 198.9 83.62 199.02 ;
      RECT 82.7 198.9 82.9 199.02 ;
      RECT 82.34 198.422 82.54 198.542 ;
      RECT 83.78 198.182 83.98 198.302 ;
      RECT 84.5 197.88 84.7 198 ;
      RECT 85.94 197.88 86.14 198 ;
      RECT 87.38 197.64 87.58 197.76 ;
      RECT 86.66 197.64 86.86 197.76 ;
      RECT 85.22 197.64 85.42 197.76 ;
      RECT 83.06 197.64 83.26 197.76 ;
      RECT 82.7 196.62 82.9 196.74 ;
      RECT 81.98 196.62 82.18 196.74 ;
      RECT 82.7 201.66 82.9 201.78 ;
      RECT 81.98 201.42 82.18 201.54 ;
      RECT 83.42 201.42 83.62 201.54 ;
      RECT 84.14 201.42 84.34 201.54 ;
      RECT 83.78 200.702 83.98 200.822 ;
      RECT 82.34 200.702 82.54 200.822 ;
      RECT 87.38 200.4 87.58 200.52 ;
      RECT 85.94 200.4 86.14 200.52 ;
      RECT 84.5 200.4 84.7 200.52 ;
      RECT 86.66 200.16 86.86 200.28 ;
      RECT 85.22 200.16 85.42 200.28 ;
      RECT 83.06 200.16 83.26 200.28 ;
      RECT 84.14 204.18 84.34 204.3 ;
      RECT 83.42 203.94 83.62 204.06 ;
      RECT 82.7 203.94 82.9 204.06 ;
      RECT 81.98 203.94 82.18 204.06 ;
      RECT 83.78 203.222 83.98 203.342 ;
      RECT 82.34 203.222 82.54 203.342 ;
      RECT 87.38 202.92 87.58 203.04 ;
      RECT 86.66 202.92 86.86 203.04 ;
      RECT 85.94 202.92 86.14 203.04 ;
      RECT 85.22 202.92 85.42 203.04 ;
      RECT 84.5 202.92 84.7 203.04 ;
      RECT 83.06 202.68 83.26 202.8 ;
      RECT 83.42 206.7 83.62 206.82 ;
      RECT 82.7 206.7 82.9 206.82 ;
      RECT 81.98 206.7 82.18 206.82 ;
      RECT 84.14 206.46 84.34 206.58 ;
      RECT 82.34 205.742 82.54 205.862 ;
      RECT 83.78 205.742 83.98 205.862 ;
      RECT 83.06 205.44 83.26 205.56 ;
      RECT 84.5 205.44 84.7 205.56 ;
      RECT 85.22 205.44 85.42 205.56 ;
      RECT 87.38 205.44 87.58 205.56 ;
      RECT 86.66 205.2 86.86 205.32 ;
      RECT 83.06 162.6 83.26 162.72 ;
      RECT 81.98 161.1 82.18 161.22 ;
      RECT 82.7 161.1 82.9 161.22 ;
      RECT 83.42 161.1 83.62 161.22 ;
      RECT 84.14 161.1 84.34 161.22 ;
      RECT 84.14 166.38 84.34 166.5 ;
      RECT 83.42 166.14 83.62 166.26 ;
      RECT 82.7 166.14 82.9 166.26 ;
      RECT 81.98 166.14 82.18 166.26 ;
      RECT 87.38 165.12 87.58 165.24 ;
      RECT 85.94 165.12 86.14 165.24 ;
      RECT 84.5 165.12 84.7 165.24 ;
      RECT 86.66 164.88 86.86 165 ;
      RECT 85.22 164.88 85.42 165 ;
      RECT 83.06 164.88 83.26 165 ;
      RECT 84.14 163.86 84.34 163.98 ;
      RECT 82.7 163.86 82.9 163.98 ;
      RECT 82.7 168.9 82.9 169.02 ;
      RECT 81.98 168.9 82.18 169.02 ;
      RECT 83.42 168.66 83.62 168.78 ;
      RECT 84.14 168.66 84.34 168.78 ;
      RECT 87.38 167.64 87.58 167.76 ;
      RECT 86.66 167.64 86.86 167.76 ;
      RECT 83.06 167.64 83.26 167.76 ;
      RECT 84.5 167.4 84.7 167.52 ;
      RECT 85.22 167.4 85.42 167.52 ;
      RECT 85.94 167.4 86.14 167.52 ;
      RECT 84.14 171.42 84.34 171.54 ;
      RECT 83.42 171.42 83.62 171.54 ;
      RECT 82.7 171.42 82.9 171.54 ;
      RECT 81.98 171.18 82.18 171.3 ;
      RECT 87.38 170.16 87.58 170.28 ;
      RECT 85.22 170.16 85.42 170.28 ;
      RECT 84.5 170.16 84.7 170.28 ;
      RECT 83.06 170.16 83.26 170.28 ;
      RECT 86.66 169.92 86.86 170.04 ;
      RECT 85.94 169.92 86.14 170.04 ;
      RECT 84.14 173.94 84.34 174.06 ;
      RECT 81.98 173.94 82.18 174.06 ;
      RECT 83.42 173.7 83.62 173.82 ;
      RECT 82.7 173.7 82.9 173.82 ;
      RECT 86.66 172.68 86.86 172.8 ;
      RECT 85.94 172.68 86.14 172.8 ;
      RECT 85.22 172.68 85.42 172.8 ;
      RECT 84.5 172.68 84.7 172.8 ;
      RECT 83.06 172.44 83.26 172.56 ;
      RECT 87.38 172.44 87.58 172.56 ;
      RECT 86.66 177.48 86.86 177.6 ;
      RECT 84.5 177.48 84.7 177.6 ;
      RECT 81.98 176.46 82.18 176.58 ;
      RECT 84.14 176.22 84.34 176.34 ;
      RECT 83.42 176.22 83.62 176.34 ;
      RECT 82.7 176.22 82.9 176.34 ;
      RECT 87.38 175.2 87.58 175.32 ;
      RECT 85.94 175.2 86.14 175.32 ;
      RECT 85.22 175.2 85.42 175.32 ;
      RECT 83.06 175.2 83.26 175.32 ;
      RECT 84.5 174.96 84.7 175.08 ;
      RECT 86.66 174.96 86.86 175.08 ;
      RECT 86.66 180 86.86 180.12 ;
      RECT 84.5 180 84.7 180.12 ;
      RECT 83.42 178.98 83.62 179.1 ;
      RECT 82.7 178.74 82.9 178.86 ;
      RECT 84.14 178.74 84.34 178.86 ;
      RECT 81.98 178.74 82.18 178.86 ;
      RECT 87.38 177.72 87.58 177.84 ;
      RECT 85.22 177.72 85.42 177.84 ;
      RECT 85.94 177.72 86.14 177.84 ;
      RECT 83.06 177.72 83.26 177.84 ;
      RECT 87.38 182.76 87.58 182.88 ;
      RECT 86.66 182.76 86.86 182.88 ;
      RECT 85.94 182.76 86.14 182.88 ;
      RECT 84.5 182.76 84.7 182.88 ;
      RECT 85.22 182.52 85.42 182.64 ;
      RECT 83.06 182.52 83.26 182.64 ;
      RECT 84.14 181.26 84.34 181.38 ;
      RECT 83.42 181.26 83.62 181.38 ;
      RECT 82.7 181.26 82.9 181.38 ;
      RECT 81.98 181.26 82.18 181.38 ;
      RECT 87.38 180.24 87.58 180.36 ;
      RECT 85.94 180.24 86.14 180.36 ;
      RECT 85.22 180.24 85.42 180.36 ;
      RECT 83.06 180.24 83.26 180.36 ;
      RECT 84.86 185.582 85.06 185.702 ;
      RECT 86.3 185.582 86.5 185.702 ;
      RECT 87.02 185.582 87.22 185.702 ;
      RECT 87.38 185.28 87.58 185.4 ;
      RECT 86.66 185.28 86.86 185.4 ;
      RECT 85.94 185.28 86.14 185.4 ;
      RECT 84.5 185.28 84.7 185.4 ;
      RECT 85.22 185.04 85.42 185.16 ;
      RECT 83.06 185.04 83.26 185.16 ;
      RECT 83.42 184.02 83.62 184.14 ;
      RECT 81.98 184.02 82.18 184.14 ;
      RECT 82.7 183.78 82.9 183.9 ;
      RECT 84.14 183.78 84.34 183.9 ;
      RECT 86.66 187.8 86.86 187.92 ;
      RECT 85.22 187.8 85.42 187.92 ;
      RECT 83.06 187.8 83.26 187.92 ;
      RECT 84.5 187.56 84.7 187.68 ;
      RECT 85.94 187.56 86.14 187.68 ;
      RECT 87.38 187.56 87.58 187.68 ;
      RECT 76.94 325.9425 77.14 326.0625 ;
      RECT 77.66 325.9425 77.86 326.0625 ;
      RECT 75.86 348.339 76.06 348.459 ;
      RECT 77.3 348.339 77.5 348.459 ;
      RECT 81.62 348.339 81.82 348.459 ;
      RECT 83.42 118.5 83.62 118.62 ;
      RECT 84.14 118.26 84.34 118.38 ;
      RECT 82.7 118.26 82.9 118.38 ;
      RECT 81.98 118.26 82.18 118.38 ;
      RECT 83.42 133.62 83.62 133.74 ;
      RECT 81.98 133.62 82.18 133.74 ;
      RECT 82.7 133.38 82.9 133.5 ;
      RECT 84.14 133.38 84.34 133.5 ;
      RECT 81.98 135.9 82.18 136.02 ;
      RECT 81.98 134.098 82.18 134.218 ;
      RECT 82.7 134.098 82.9 134.218 ;
      RECT 83.42 134.098 83.62 134.218 ;
      RECT 84.14 134.098 84.34 134.218 ;
      RECT 81.98 139.138 82.18 139.258 ;
      RECT 81.98 138.42 82.18 138.54 ;
      RECT 81.98 136.618 82.18 136.738 ;
      RECT 83.42 141.18 83.62 141.3 ;
      RECT 81.98 140.94 82.18 141.06 ;
      RECT 82.7 140.94 82.9 141.06 ;
      RECT 84.14 140.94 84.34 141.06 ;
      RECT 83.42 143.7 83.62 143.82 ;
      RECT 84.14 143.46 84.34 143.58 ;
      RECT 82.7 143.46 82.9 143.58 ;
      RECT 81.98 143.46 82.18 143.58 ;
      RECT 85.22 142.44 85.42 142.56 ;
      RECT 85.94 142.44 86.14 142.56 ;
      RECT 86.66 142.44 86.86 142.56 ;
      RECT 87.38 142.2 87.58 142.32 ;
      RECT 84.5 142.2 84.7 142.32 ;
      RECT 83.06 142.2 83.26 142.32 ;
      RECT 81.98 145.98 82.18 146.1 ;
      RECT 82.7 145.98 82.9 146.1 ;
      RECT 83.42 145.98 83.62 146.1 ;
      RECT 84.14 145.98 84.34 146.1 ;
      RECT 83.06 144.96 83.26 145.08 ;
      RECT 84.5 144.96 84.7 145.08 ;
      RECT 86.66 144.96 86.86 145.08 ;
      RECT 87.38 144.96 87.58 145.08 ;
      RECT 85.22 144.72 85.42 144.84 ;
      RECT 85.94 144.72 86.14 144.84 ;
      RECT 86.66 150 86.86 150.12 ;
      RECT 85.22 150 85.42 150.12 ;
      RECT 84.5 150 84.7 150.12 ;
      RECT 87.38 149.76 87.58 149.88 ;
      RECT 85.94 149.76 86.14 149.88 ;
      RECT 83.06 149.76 83.26 149.88 ;
      RECT 82.7 148.74 82.9 148.86 ;
      RECT 81.98 148.5 82.18 148.62 ;
      RECT 83.42 148.5 83.62 148.62 ;
      RECT 84.14 148.5 84.34 148.62 ;
      RECT 87.38 152.52 87.58 152.64 ;
      RECT 85.94 152.52 86.14 152.64 ;
      RECT 84.5 152.52 84.7 152.64 ;
      RECT 83.06 152.52 83.26 152.64 ;
      RECT 86.66 152.28 86.86 152.4 ;
      RECT 85.22 152.28 85.42 152.4 ;
      RECT 81.98 151.26 82.18 151.38 ;
      RECT 82.7 151.26 82.9 151.38 ;
      RECT 84.14 151.02 84.34 151.14 ;
      RECT 83.42 151.02 83.62 151.14 ;
      RECT 87.38 155.04 87.58 155.16 ;
      RECT 86.66 155.04 86.86 155.16 ;
      RECT 85.94 155.04 86.14 155.16 ;
      RECT 84.5 155.04 84.7 155.16 ;
      RECT 83.06 155.04 83.26 155.16 ;
      RECT 85.22 154.8 85.42 154.92 ;
      RECT 84.14 153.78 84.34 153.9 ;
      RECT 82.7 153.78 82.9 153.9 ;
      RECT 81.98 153.54 82.18 153.66 ;
      RECT 83.42 153.54 83.62 153.66 ;
      RECT 87.38 157.56 87.58 157.68 ;
      RECT 85.94 157.56 86.14 157.68 ;
      RECT 83.06 157.56 83.26 157.68 ;
      RECT 86.66 157.32 86.86 157.44 ;
      RECT 85.22 157.32 85.42 157.44 ;
      RECT 84.5 157.32 84.7 157.44 ;
      RECT 82.7 156.3 82.9 156.42 ;
      RECT 84.14 156.06 84.34 156.18 ;
      RECT 83.42 156.06 83.62 156.18 ;
      RECT 81.98 156.06 82.18 156.18 ;
      RECT 84.5 160.08 84.7 160.2 ;
      RECT 85.22 160.08 85.42 160.2 ;
      RECT 85.94 160.08 86.14 160.2 ;
      RECT 87.38 160.08 87.58 160.2 ;
      RECT 86.66 159.84 86.86 159.96 ;
      RECT 83.06 159.84 83.26 159.96 ;
      RECT 84.14 158.82 84.34 158.94 ;
      RECT 83.42 158.58 83.62 158.7 ;
      RECT 82.7 158.58 82.9 158.7 ;
      RECT 81.98 158.58 82.18 158.7 ;
      RECT 81.98 163.62 82.18 163.74 ;
      RECT 83.42 163.62 83.62 163.74 ;
      RECT 87.38 162.6 87.58 162.72 ;
      RECT 86.66 162.6 86.86 162.72 ;
      RECT 85.94 162.6 86.14 162.72 ;
      RECT 85.22 162.6 85.42 162.72 ;
      RECT 84.5 162.6 84.7 162.72 ;
      RECT 80.9 263.16 81.1 263.28 ;
      RECT 81.62 262.53 81.82 262.65 ;
      RECT 77.3 262.53 77.5 262.65 ;
      RECT 75.86 262.53 76.06 262.65 ;
      RECT 81.26 262.14 81.46 262.26 ;
      RECT 80.54 262.14 80.74 262.26 ;
      RECT 76.94 262.14 77.14 262.26 ;
      RECT 76.22 262.14 76.42 262.26 ;
      RECT 74.78 262.14 74.98 262.26 ;
      RECT 80.54 267.18 80.74 267.3 ;
      RECT 76.94 267.18 77.14 267.3 ;
      RECT 75.5 267.18 75.7 267.3 ;
      RECT 74.78 267.18 74.98 267.3 ;
      RECT 81.26 266.94 81.46 267.06 ;
      RECT 78.38 266.94 78.58 267.06 ;
      RECT 77.66 266.94 77.86 267.06 ;
      RECT 76.22 266.94 76.42 267.06 ;
      RECT 77.3 266.2885 77.5 266.4085 ;
      RECT 81.62 266.2885 81.82 266.4085 ;
      RECT 75.86 266.2885 76.06 266.4085 ;
      RECT 78.02 265.92 78.22 266.04 ;
      RECT 80.9 265.68 81.1 265.8 ;
      RECT 76.58 265.68 76.78 265.8 ;
      RECT 75.14 265.68 75.34 265.8 ;
      RECT 81.62 270.09 81.82 270.21 ;
      RECT 75.86 270.09 76.06 270.21 ;
      RECT 80.54 269.7 80.74 269.82 ;
      RECT 78.38 269.7 78.58 269.82 ;
      RECT 76.94 269.7 77.14 269.82 ;
      RECT 76.22 269.7 76.42 269.82 ;
      RECT 74.78 269.7 74.98 269.82 ;
      RECT 81.26 269.46 81.46 269.58 ;
      RECT 77.66 269.46 77.86 269.58 ;
      RECT 75.5 269.46 75.7 269.58 ;
      RECT 78.02 268.44 78.22 268.56 ;
      RECT 80.9 268.2 81.1 268.32 ;
      RECT 76.58 268.2 76.78 268.32 ;
      RECT 75.14 268.2 75.34 268.32 ;
      RECT 77.3 267.81 77.5 267.93 ;
      RECT 75.86 267.81 76.06 267.93 ;
      RECT 81.62 267.81 81.82 267.93 ;
      RECT 80.54 272.22 80.74 272.34 ;
      RECT 78.38 272.22 78.58 272.34 ;
      RECT 76.94 272.22 77.14 272.34 ;
      RECT 76.22 272.22 76.42 272.34 ;
      RECT 74.78 271.98 74.98 272.1 ;
      RECT 75.5 271.98 75.7 272.1 ;
      RECT 81.26 271.98 81.46 272.1 ;
      RECT 77.66 271.98 77.86 272.1 ;
      RECT 75.86 271.59 76.06 271.71 ;
      RECT 81.62 271.35 81.82 271.47 ;
      RECT 77.3 271.35 77.5 271.47 ;
      RECT 80.9 270.96 81.1 271.08 ;
      RECT 76.58 270.96 76.78 271.08 ;
      RECT 78.02 270.72 78.22 270.84 ;
      RECT 75.14 270.72 75.34 270.84 ;
      RECT 77.3 270.33 77.5 270.45 ;
      RECT 78.02 275.76 78.22 275.88 ;
      RECT 75.14 275.76 75.34 275.88 ;
      RECT 81.26 274.74 81.46 274.86 ;
      RECT 77.66 274.74 77.86 274.86 ;
      RECT 76.94 274.74 77.14 274.86 ;
      RECT 76.22 274.74 76.42 274.86 ;
      RECT 75.5 274.74 75.7 274.86 ;
      RECT 80.54 274.5 80.74 274.62 ;
      RECT 78.38 274.5 78.58 274.62 ;
      RECT 74.78 274.5 74.98 274.62 ;
      RECT 80.9 273.48 81.1 273.6 ;
      RECT 76.58 273.48 76.78 273.6 ;
      RECT 78.02 273.24 78.22 273.36 ;
      RECT 75.14 273.24 75.34 273.36 ;
      RECT 78.02 278.28 78.22 278.4 ;
      RECT 75.14 278.28 75.34 278.4 ;
      RECT 81.26 277.26 81.46 277.38 ;
      RECT 80.54 277.26 80.74 277.38 ;
      RECT 77.66 277.26 77.86 277.38 ;
      RECT 76.22 277.26 76.42 277.38 ;
      RECT 78.38 277.02 78.58 277.14 ;
      RECT 76.94 277.02 77.14 277.14 ;
      RECT 75.5 277.02 75.7 277.14 ;
      RECT 74.78 277.02 74.98 277.14 ;
      RECT 80.9 276 81.1 276.12 ;
      RECT 76.58 276 76.78 276.12 ;
      RECT 80.9 278.52 81.1 278.64 ;
      RECT 76.58 278.52 76.78 278.64 ;
      RECT 81.26 308.496 81.46 308.616 ;
      RECT 80.54 308.496 80.74 308.616 ;
      RECT 78.38 308.496 78.58 308.616 ;
      RECT 77.66 308.496 77.86 308.616 ;
      RECT 76.94 308.496 77.14 308.616 ;
      RECT 76.22 308.496 76.42 308.616 ;
      RECT 75.5 308.496 75.7 308.616 ;
      RECT 74.78 308.496 74.98 308.616 ;
      RECT 75.86 323.3835 76.06 323.5035 ;
      RECT 77.3 323.3835 77.5 323.5035 ;
      RECT 81.62 323.3835 81.82 323.5035 ;
      RECT 78.38 325.9425 78.58 326.0625 ;
      RECT 80.54 325.9425 80.74 326.0625 ;
      RECT 81.26 325.9425 81.46 326.0625 ;
      RECT 74.78 325.9425 74.98 326.0625 ;
      RECT 75.5 325.9425 75.7 326.0625 ;
      RECT 76.22 325.9425 76.42 326.0625 ;
      RECT 75.5 244.5 75.7 244.62 ;
      RECT 77.66 244.5 77.86 244.62 ;
      RECT 81.26 244.5 81.46 244.62 ;
      RECT 80.54 244.26 80.74 244.38 ;
      RECT 78.38 244.26 78.58 244.38 ;
      RECT 76.94 244.26 77.14 244.38 ;
      RECT 76.22 244.26 76.42 244.38 ;
      RECT 74.78 244.26 74.98 244.38 ;
      RECT 78.38 247.02 78.58 247.14 ;
      RECT 77.66 247.02 77.86 247.14 ;
      RECT 76.94 247.02 77.14 247.14 ;
      RECT 74.78 247.02 74.98 247.14 ;
      RECT 81.26 246.78 81.46 246.9 ;
      RECT 80.54 246.78 80.74 246.9 ;
      RECT 76.22 246.78 76.42 246.9 ;
      RECT 75.5 246.78 75.7 246.9 ;
      RECT 80.9 250.8 81.1 250.92 ;
      RECT 78.02 250.56 78.22 250.68 ;
      RECT 76.58 250.56 76.78 250.68 ;
      RECT 75.14 250.56 75.34 250.68 ;
      RECT 81.26 249.54 81.46 249.66 ;
      RECT 77.66 249.54 77.86 249.66 ;
      RECT 76.22 249.54 76.42 249.66 ;
      RECT 74.78 249.54 74.98 249.66 ;
      RECT 80.54 249.3 80.74 249.42 ;
      RECT 78.38 249.3 78.58 249.42 ;
      RECT 76.94 249.3 77.14 249.42 ;
      RECT 75.5 249.3 75.7 249.42 ;
      RECT 76.58 253.32 76.78 253.44 ;
      RECT 75.14 253.32 75.34 253.44 ;
      RECT 80.9 253.08 81.1 253.2 ;
      RECT 78.02 253.08 78.22 253.2 ;
      RECT 80.54 252.06 80.74 252.18 ;
      RECT 77.66 252.06 77.86 252.18 ;
      RECT 76.94 252.06 77.14 252.18 ;
      RECT 75.5 252.06 75.7 252.18 ;
      RECT 74.78 252.06 74.98 252.18 ;
      RECT 81.26 251.82 81.46 251.94 ;
      RECT 78.38 251.82 78.58 251.94 ;
      RECT 76.22 251.82 76.42 251.94 ;
      RECT 80.9 255.84 81.1 255.96 ;
      RECT 76.58 255.84 76.78 255.96 ;
      RECT 78.02 255.6 78.22 255.72 ;
      RECT 75.14 255.6 75.34 255.72 ;
      RECT 81.26 254.58 81.46 254.7 ;
      RECT 77.66 254.58 77.86 254.7 ;
      RECT 76.22 254.58 76.42 254.7 ;
      RECT 74.78 254.58 74.98 254.7 ;
      RECT 80.54 254.34 80.74 254.46 ;
      RECT 78.38 254.34 78.58 254.46 ;
      RECT 76.94 254.34 77.14 254.46 ;
      RECT 75.5 254.34 75.7 254.46 ;
      RECT 81.26 259.38 81.46 259.5 ;
      RECT 78.38 259.38 78.58 259.5 ;
      RECT 76.94 259.38 77.14 259.5 ;
      RECT 75.5 259.38 75.7 259.5 ;
      RECT 81.62 258.99 81.82 259.11 ;
      RECT 77.3 258.99 77.5 259.11 ;
      RECT 75.86 258.75 76.06 258.87 ;
      RECT 78.02 258.36 78.22 258.48 ;
      RECT 75.14 258.36 75.34 258.48 ;
      RECT 80.9 258.12 81.1 258.24 ;
      RECT 76.58 258.12 76.78 258.24 ;
      RECT 77.66 257.1 77.86 257.22 ;
      RECT 76.22 257.1 76.42 257.22 ;
      RECT 74.78 257.1 74.98 257.22 ;
      RECT 78.38 256.86 78.58 256.98 ;
      RECT 80.54 256.86 80.74 256.98 ;
      RECT 81.26 256.86 81.46 256.98 ;
      RECT 76.94 256.86 77.14 256.98 ;
      RECT 75.5 256.86 75.7 256.98 ;
      RECT 78.38 261.9 78.58 262.02 ;
      RECT 77.66 261.9 77.86 262.02 ;
      RECT 75.5 261.9 75.7 262.02 ;
      RECT 81.62 261.51 81.82 261.63 ;
      RECT 75.86 261.51 76.06 261.63 ;
      RECT 77.3 261.27 77.5 261.39 ;
      RECT 78.02 260.88 78.22 261 ;
      RECT 80.9 260.64 81.1 260.76 ;
      RECT 76.58 260.64 76.78 260.76 ;
      RECT 75.14 260.64 75.34 260.76 ;
      RECT 77.3 260.25 77.5 260.37 ;
      RECT 75.86 260.25 76.06 260.37 ;
      RECT 81.62 260.01 81.82 260.13 ;
      RECT 80.54 259.62 80.74 259.74 ;
      RECT 77.66 259.62 77.86 259.74 ;
      RECT 76.22 259.62 76.42 259.74 ;
      RECT 74.78 259.62 74.98 259.74 ;
      RECT 76.94 264.66 77.14 264.78 ;
      RECT 80.54 264.66 80.74 264.78 ;
      RECT 75.5 264.66 75.7 264.78 ;
      RECT 81.26 264.42 81.46 264.54 ;
      RECT 78.38 264.42 78.58 264.54 ;
      RECT 77.66 264.42 77.86 264.54 ;
      RECT 76.22 264.42 76.42 264.54 ;
      RECT 74.78 264.42 74.98 264.54 ;
      RECT 77.3 264.03 77.5 264.15 ;
      RECT 81.62 263.79 81.82 263.91 ;
      RECT 75.86 263.79 76.06 263.91 ;
      RECT 78.02 263.4 78.22 263.52 ;
      RECT 76.58 263.4 76.78 263.52 ;
      RECT 75.14 263.4 75.34 263.52 ;
      RECT 77.66 211.74 77.86 211.86 ;
      RECT 76.22 211.74 76.42 211.86 ;
      RECT 80.54 211.5 80.74 211.62 ;
      RECT 78.38 211.5 78.58 211.62 ;
      RECT 76.94 211.5 77.14 211.62 ;
      RECT 75.5 211.5 75.7 211.62 ;
      RECT 74.78 211.5 74.98 211.62 ;
      RECT 75.14 211.198 75.34 211.318 ;
      RECT 78.02 211.198 78.22 211.318 ;
      RECT 76.58 210.958 76.78 211.078 ;
      RECT 80.9 210.958 81.1 211.078 ;
      RECT 77.3 215.52 77.5 215.64 ;
      RECT 75.86 215.52 76.06 215.64 ;
      RECT 81.62 215.28 81.82 215.4 ;
      RECT 81.26 214.26 81.46 214.38 ;
      RECT 80.54 214.26 80.74 214.38 ;
      RECT 78.38 214.26 78.58 214.38 ;
      RECT 76.22 214.26 76.42 214.38 ;
      RECT 75.5 214.26 75.7 214.38 ;
      RECT 77.66 214.02 77.86 214.14 ;
      RECT 76.94 214.02 77.14 214.14 ;
      RECT 74.78 214.02 74.98 214.14 ;
      RECT 81.62 213 81.82 213.12 ;
      RECT 81.26 216.78 81.46 216.9 ;
      RECT 78.38 216.78 78.58 216.9 ;
      RECT 76.22 216.78 76.42 216.9 ;
      RECT 75.5 216.78 75.7 216.9 ;
      RECT 80.54 216.54 80.74 216.66 ;
      RECT 77.66 216.54 77.86 216.66 ;
      RECT 76.94 216.54 77.14 216.66 ;
      RECT 74.78 216.54 74.98 216.66 ;
      RECT 81.26 219.3 81.46 219.42 ;
      RECT 80.54 219.3 80.74 219.42 ;
      RECT 77.66 219.3 77.86 219.42 ;
      RECT 76.22 219.3 76.42 219.42 ;
      RECT 75.5 219.3 75.7 219.42 ;
      RECT 74.78 219.06 74.98 219.18 ;
      RECT 76.94 219.06 77.14 219.18 ;
      RECT 78.38 219.06 78.58 219.18 ;
      RECT 74.78 223.798 74.98 223.918 ;
      RECT 76.22 223.798 76.42 223.918 ;
      RECT 76.94 223.798 77.14 223.918 ;
      RECT 77.66 223.798 77.86 223.918 ;
      RECT 78.38 223.798 78.58 223.918 ;
      RECT 75.5 223.558 75.7 223.678 ;
      RECT 80.54 223.558 80.74 223.678 ;
      RECT 81.26 223.558 81.46 223.678 ;
      RECT 75.86 223.08 76.06 223.2 ;
      RECT 77.3 223.08 77.5 223.2 ;
      RECT 81.62 222.84 81.82 222.96 ;
      RECT 75.14 222.362 75.34 222.482 ;
      RECT 78.02 222.362 78.22 222.482 ;
      RECT 76.58 222.122 76.78 222.242 ;
      RECT 80.9 222.122 81.1 222.242 ;
      RECT 76.22 229.14 76.42 229.26 ;
      RECT 76.94 229.14 77.14 229.26 ;
      RECT 78.38 229.14 78.58 229.26 ;
      RECT 80.54 229.14 80.74 229.26 ;
      RECT 81.26 229.14 81.46 229.26 ;
      RECT 81.26 231.9 81.46 232.02 ;
      RECT 80.54 231.9 80.74 232.02 ;
      RECT 76.94 231.9 77.14 232.02 ;
      RECT 76.22 231.9 76.42 232.02 ;
      RECT 74.78 231.9 74.98 232.02 ;
      RECT 78.38 231.66 78.58 231.78 ;
      RECT 77.66 231.66 77.86 231.78 ;
      RECT 75.5 231.66 75.7 231.78 ;
      RECT 74.78 229.38 74.98 229.5 ;
      RECT 75.5 229.38 75.7 229.5 ;
      RECT 77.66 229.38 77.86 229.5 ;
      RECT 77.66 234.42 77.86 234.54 ;
      RECT 76.22 234.42 76.42 234.54 ;
      RECT 80.54 234.42 80.74 234.54 ;
      RECT 78.38 234.42 78.58 234.54 ;
      RECT 74.78 234.18 74.98 234.3 ;
      RECT 75.5 234.18 75.7 234.3 ;
      RECT 76.94 234.18 77.14 234.3 ;
      RECT 81.26 234.18 81.46 234.3 ;
      RECT 81.26 236.94 81.46 237.06 ;
      RECT 80.54 236.94 80.74 237.06 ;
      RECT 77.66 236.94 77.86 237.06 ;
      RECT 76.94 236.94 77.14 237.06 ;
      RECT 76.22 236.94 76.42 237.06 ;
      RECT 74.78 236.7 74.98 236.82 ;
      RECT 75.5 236.7 75.7 236.82 ;
      RECT 78.38 236.7 78.58 236.82 ;
      RECT 81.26 239.46 81.46 239.58 ;
      RECT 80.54 239.46 80.74 239.58 ;
      RECT 77.66 239.46 77.86 239.58 ;
      RECT 75.5 239.46 75.7 239.58 ;
      RECT 78.38 239.22 78.58 239.34 ;
      RECT 76.94 239.22 77.14 239.34 ;
      RECT 76.22 239.22 76.42 239.34 ;
      RECT 74.78 239.22 74.98 239.34 ;
      RECT 74.78 241.98 74.98 242.1 ;
      RECT 75.5 241.98 75.7 242.1 ;
      RECT 76.22 241.98 76.42 242.1 ;
      RECT 76.94 241.98 77.14 242.1 ;
      RECT 80.54 241.98 80.74 242.1 ;
      RECT 77.66 241.74 77.86 241.86 ;
      RECT 78.38 241.74 78.58 241.86 ;
      RECT 81.26 241.74 81.46 241.86 ;
      RECT 81.26 194.1 81.46 194.22 ;
      RECT 78.38 194.1 78.58 194.22 ;
      RECT 77.66 194.1 77.86 194.22 ;
      RECT 76.94 194.1 77.14 194.22 ;
      RECT 75.5 194.1 75.7 194.22 ;
      RECT 74.78 194.1 74.98 194.22 ;
      RECT 77.3 195.12 77.5 195.24 ;
      RECT 75.86 195.12 76.06 195.24 ;
      RECT 81.62 195.36 81.82 195.48 ;
      RECT 76.58 195.662 76.78 195.782 ;
      RECT 78.02 195.662 78.22 195.782 ;
      RECT 80.9 195.662 81.1 195.782 ;
      RECT 75.14 195.902 75.34 196.022 ;
      RECT 81.26 196.38 81.46 196.5 ;
      RECT 77.66 196.38 77.86 196.5 ;
      RECT 76.22 196.38 76.42 196.5 ;
      RECT 75.5 196.38 75.7 196.5 ;
      RECT 74.78 196.62 74.98 196.74 ;
      RECT 76.94 196.62 77.14 196.74 ;
      RECT 78.38 196.62 78.58 196.74 ;
      RECT 80.54 196.62 80.74 196.74 ;
      RECT 75.86 197.64 76.06 197.76 ;
      RECT 81.62 197.64 81.82 197.76 ;
      RECT 77.3 197.88 77.5 198 ;
      RECT 80.9 198.182 81.1 198.302 ;
      RECT 78.02 198.182 78.22 198.302 ;
      RECT 75.14 198.182 75.34 198.302 ;
      RECT 76.58 198.422 76.78 198.542 ;
      RECT 74.78 198.9 74.98 199.02 ;
      RECT 76.22 198.9 76.42 199.02 ;
      RECT 76.94 198.9 77.14 199.02 ;
      RECT 81.26 199.14 81.46 199.26 ;
      RECT 80.54 199.14 80.74 199.26 ;
      RECT 78.38 199.14 78.58 199.26 ;
      RECT 77.66 199.14 77.86 199.26 ;
      RECT 75.5 199.14 75.7 199.26 ;
      RECT 74.78 201.66 74.98 201.78 ;
      RECT 75.5 201.66 75.7 201.78 ;
      RECT 77.66 201.66 77.86 201.78 ;
      RECT 81.26 201.66 81.46 201.78 ;
      RECT 76.22 201.42 76.42 201.54 ;
      RECT 76.94 201.42 77.14 201.54 ;
      RECT 78.38 201.42 78.58 201.54 ;
      RECT 80.54 201.42 80.74 201.54 ;
      RECT 76.58 200.942 76.78 201.062 ;
      RECT 80.9 200.702 81.1 200.822 ;
      RECT 78.02 200.702 78.22 200.822 ;
      RECT 75.14 200.702 75.34 200.822 ;
      RECT 81.62 200.4 81.82 200.52 ;
      RECT 77.3 200.4 77.5 200.52 ;
      RECT 75.86 200.16 76.06 200.28 ;
      RECT 77.66 204.18 77.86 204.3 ;
      RECT 80.54 204.18 80.74 204.3 ;
      RECT 81.26 204.18 81.46 204.3 ;
      RECT 76.22 204.18 76.42 204.3 ;
      RECT 76.94 204.18 77.14 204.3 ;
      RECT 78.38 203.94 78.58 204.06 ;
      RECT 75.5 203.94 75.7 204.06 ;
      RECT 74.78 203.94 74.98 204.06 ;
      RECT 78.02 203.462 78.22 203.582 ;
      RECT 75.14 203.462 75.34 203.582 ;
      RECT 80.9 203.222 81.1 203.342 ;
      RECT 76.58 203.222 76.78 203.342 ;
      RECT 77.3 202.92 77.5 203.04 ;
      RECT 75.86 202.68 76.06 202.8 ;
      RECT 81.62 202.68 81.82 202.8 ;
      RECT 77.66 206.7 77.86 206.82 ;
      RECT 76.22 206.7 76.42 206.82 ;
      RECT 75.5 206.7 75.7 206.82 ;
      RECT 81.26 206.46 81.46 206.58 ;
      RECT 80.54 206.46 80.74 206.58 ;
      RECT 78.38 206.46 78.58 206.58 ;
      RECT 76.94 206.46 77.14 206.58 ;
      RECT 74.78 206.46 74.98 206.58 ;
      RECT 78.02 205.982 78.22 206.102 ;
      RECT 76.58 205.982 76.78 206.102 ;
      RECT 75.14 205.742 75.34 205.862 ;
      RECT 80.9 205.742 81.1 205.862 ;
      RECT 75.86 205.44 76.06 205.56 ;
      RECT 77.3 205.44 77.5 205.56 ;
      RECT 81.62 205.2 81.82 205.32 ;
      RECT 75.86 210.24 76.06 210.36 ;
      RECT 77.3 210.24 77.5 210.36 ;
      RECT 81.62 210.24 81.82 210.36 ;
      RECT 80.54 209.22 80.74 209.34 ;
      RECT 76.22 209.22 76.42 209.34 ;
      RECT 75.5 209.22 75.7 209.34 ;
      RECT 74.78 209.22 74.98 209.34 ;
      RECT 76.94 208.98 77.14 209.1 ;
      RECT 77.66 208.98 77.86 209.1 ;
      RECT 78.38 208.98 78.58 209.1 ;
      RECT 81.26 208.98 81.46 209.1 ;
      RECT 75.14 208.502 75.34 208.622 ;
      RECT 78.02 208.502 78.22 208.622 ;
      RECT 76.58 208.262 76.78 208.382 ;
      RECT 80.9 208.262 81.1 208.382 ;
      RECT 77.3 207.96 77.5 208.08 ;
      RECT 75.86 207.96 76.06 208.08 ;
      RECT 81.62 207.72 81.82 207.84 ;
      RECT 75.86 212.76 76.06 212.88 ;
      RECT 77.3 212.76 77.5 212.88 ;
      RECT 81.26 211.74 81.46 211.86 ;
      RECT 76.94 173.7 77.14 173.82 ;
      RECT 81.62 172.68 81.82 172.8 ;
      RECT 75.86 172.44 76.06 172.56 ;
      RECT 77.3 172.44 77.5 172.56 ;
      RECT 75.86 177.48 76.06 177.6 ;
      RECT 80.54 176.46 80.74 176.58 ;
      RECT 77.66 176.46 77.86 176.58 ;
      RECT 76.22 176.46 76.42 176.58 ;
      RECT 74.78 176.46 74.98 176.58 ;
      RECT 81.26 176.22 81.46 176.34 ;
      RECT 78.38 176.22 78.58 176.34 ;
      RECT 76.94 176.22 77.14 176.34 ;
      RECT 75.5 176.22 75.7 176.34 ;
      RECT 77.3 175.2 77.5 175.32 ;
      RECT 75.86 174.96 76.06 175.08 ;
      RECT 81.62 174.96 81.82 175.08 ;
      RECT 75.86 180 76.06 180.12 ;
      RECT 81.26 178.98 81.46 179.1 ;
      RECT 76.22 178.98 76.42 179.1 ;
      RECT 74.78 178.98 74.98 179.1 ;
      RECT 80.54 178.74 80.74 178.86 ;
      RECT 78.38 178.74 78.58 178.86 ;
      RECT 77.66 178.74 77.86 178.86 ;
      RECT 76.94 178.74 77.14 178.86 ;
      RECT 75.5 178.74 75.7 178.86 ;
      RECT 81.62 177.72 81.82 177.84 ;
      RECT 77.3 177.72 77.5 177.84 ;
      RECT 77.3 182.76 77.5 182.88 ;
      RECT 81.62 182.52 81.82 182.64 ;
      RECT 75.86 182.52 76.06 182.64 ;
      RECT 74.78 181.5 74.98 181.62 ;
      RECT 81.26 181.5 81.46 181.62 ;
      RECT 80.54 181.5 80.74 181.62 ;
      RECT 78.38 181.5 78.58 181.62 ;
      RECT 76.94 181.5 77.14 181.62 ;
      RECT 75.5 181.26 75.7 181.38 ;
      RECT 77.66 181.26 77.86 181.38 ;
      RECT 76.22 181.26 76.42 181.38 ;
      RECT 81.62 180.24 81.82 180.36 ;
      RECT 77.3 180.24 77.5 180.36 ;
      RECT 75.86 185.28 76.06 185.4 ;
      RECT 81.62 185.04 81.82 185.16 ;
      RECT 77.3 185.04 77.5 185.16 ;
      RECT 76.94 184.02 77.14 184.14 ;
      RECT 74.78 184.02 74.98 184.14 ;
      RECT 75.5 183.78 75.7 183.9 ;
      RECT 76.22 183.78 76.42 183.9 ;
      RECT 77.66 183.78 77.86 183.9 ;
      RECT 78.38 183.78 78.58 183.9 ;
      RECT 80.54 183.78 80.74 183.9 ;
      RECT 81.26 183.78 81.46 183.9 ;
      RECT 75.86 187.8 76.06 187.92 ;
      RECT 77.3 187.56 77.5 187.68 ;
      RECT 81.62 187.56 81.82 187.68 ;
      RECT 74.78 186.54 74.98 186.66 ;
      RECT 76.22 186.54 76.42 186.66 ;
      RECT 77.66 186.54 77.86 186.66 ;
      RECT 80.54 186.54 80.74 186.66 ;
      RECT 81.26 186.54 81.46 186.66 ;
      RECT 75.5 186.3 75.7 186.42 ;
      RECT 76.94 186.3 77.14 186.42 ;
      RECT 78.38 186.3 78.58 186.42 ;
      RECT 75.14 190.862 75.34 190.982 ;
      RECT 78.02 190.862 78.22 190.982 ;
      RECT 76.58 190.622 76.78 190.742 ;
      RECT 80.9 190.622 81.1 190.742 ;
      RECT 75.86 190.32 76.06 190.44 ;
      RECT 81.62 190.32 81.82 190.44 ;
      RECT 77.3 190.08 77.5 190.2 ;
      RECT 74.78 189.06 74.98 189.18 ;
      RECT 76.94 189.06 77.14 189.18 ;
      RECT 77.66 189.06 77.86 189.18 ;
      RECT 81.26 189.06 81.46 189.18 ;
      RECT 80.54 188.82 80.74 188.94 ;
      RECT 78.38 188.82 78.58 188.94 ;
      RECT 76.22 188.82 76.42 188.94 ;
      RECT 75.5 188.82 75.7 188.94 ;
      RECT 76.22 193.86 76.42 193.98 ;
      RECT 80.54 193.86 80.74 193.98 ;
      RECT 75.14 193.382 75.34 193.502 ;
      RECT 76.58 193.142 76.78 193.262 ;
      RECT 78.02 193.142 78.22 193.262 ;
      RECT 80.9 193.142 81.1 193.262 ;
      RECT 81.62 192.84 81.82 192.96 ;
      RECT 75.86 192.84 76.06 192.96 ;
      RECT 77.3 192.6 77.5 192.72 ;
      RECT 75.14 192.122 75.34 192.242 ;
      RECT 80.9 192.122 81.1 192.242 ;
      RECT 76.58 191.882 76.78 192.002 ;
      RECT 78.02 191.882 78.22 192.002 ;
      RECT 80.54 191.58 80.74 191.7 ;
      RECT 78.38 191.58 78.58 191.7 ;
      RECT 76.94 191.58 77.14 191.7 ;
      RECT 75.5 191.58 75.7 191.7 ;
      RECT 74.78 191.58 74.98 191.7 ;
      RECT 76.22 191.34 76.42 191.46 ;
      RECT 77.66 191.34 77.86 191.46 ;
      RECT 81.26 191.34 81.46 191.46 ;
      RECT 76.58 194.642 76.78 194.762 ;
      RECT 80.9 194.402 81.1 194.522 ;
      RECT 78.02 194.402 78.22 194.522 ;
      RECT 75.14 194.402 75.34 194.522 ;
      RECT 76.94 151.02 77.14 151.14 ;
      RECT 75.5 151.02 75.7 151.14 ;
      RECT 81.62 155.04 81.82 155.16 ;
      RECT 75.86 155.04 76.06 155.16 ;
      RECT 77.3 154.8 77.5 154.92 ;
      RECT 80.54 153.78 80.74 153.9 ;
      RECT 77.66 153.78 77.86 153.9 ;
      RECT 75.5 153.78 75.7 153.9 ;
      RECT 74.78 153.54 74.98 153.66 ;
      RECT 76.22 153.54 76.42 153.66 ;
      RECT 76.94 153.54 77.14 153.66 ;
      RECT 78.38 153.54 78.58 153.66 ;
      RECT 81.26 153.54 81.46 153.66 ;
      RECT 76.58 158.278 76.78 158.398 ;
      RECT 75.14 158.278 75.34 158.398 ;
      RECT 80.9 158.038 81.1 158.158 ;
      RECT 78.02 158.038 78.22 158.158 ;
      RECT 81.62 157.56 81.82 157.68 ;
      RECT 75.86 157.56 76.06 157.68 ;
      RECT 77.3 157.32 77.5 157.44 ;
      RECT 80.9 156.602 81.1 156.722 ;
      RECT 78.02 156.602 78.22 156.722 ;
      RECT 76.58 156.602 76.78 156.722 ;
      RECT 75.14 156.602 75.34 156.722 ;
      RECT 75.5 156.3 75.7 156.42 ;
      RECT 77.66 156.3 77.86 156.42 ;
      RECT 76.22 156.3 76.42 156.42 ;
      RECT 81.26 156.3 81.46 156.42 ;
      RECT 80.54 156.06 80.74 156.18 ;
      RECT 78.38 156.06 78.58 156.18 ;
      RECT 76.94 156.06 77.14 156.18 ;
      RECT 74.78 156.06 74.98 156.18 ;
      RECT 75.86 160.08 76.06 160.2 ;
      RECT 81.62 160.08 81.82 160.2 ;
      RECT 77.3 159.84 77.5 159.96 ;
      RECT 81.26 158.82 81.46 158.94 ;
      RECT 77.66 158.82 77.86 158.94 ;
      RECT 74.78 158.82 74.98 158.94 ;
      RECT 80.54 158.58 80.74 158.7 ;
      RECT 78.38 158.58 78.58 158.7 ;
      RECT 76.94 158.58 77.14 158.7 ;
      RECT 76.22 158.58 76.42 158.7 ;
      RECT 75.5 158.58 75.7 158.7 ;
      RECT 74.78 163.62 74.98 163.74 ;
      RECT 76.94 163.62 77.14 163.74 ;
      RECT 77.66 163.62 77.86 163.74 ;
      RECT 81.26 163.62 81.46 163.74 ;
      RECT 81.62 162.6 81.82 162.72 ;
      RECT 77.3 162.6 77.5 162.72 ;
      RECT 75.86 162.6 76.06 162.72 ;
      RECT 74.78 161.1 74.98 161.22 ;
      RECT 75.5 161.1 75.7 161.22 ;
      RECT 76.22 161.1 76.42 161.22 ;
      RECT 76.94 161.1 77.14 161.22 ;
      RECT 77.66 161.1 77.86 161.22 ;
      RECT 78.38 161.1 78.58 161.22 ;
      RECT 80.54 161.1 80.74 161.22 ;
      RECT 81.26 161.1 81.46 161.22 ;
      RECT 76.22 166.38 76.42 166.5 ;
      RECT 75.5 166.38 75.7 166.5 ;
      RECT 76.94 166.38 77.14 166.5 ;
      RECT 78.38 166.38 78.58 166.5 ;
      RECT 80.54 166.38 80.74 166.5 ;
      RECT 81.26 166.38 81.46 166.5 ;
      RECT 77.66 166.14 77.86 166.26 ;
      RECT 74.78 166.14 74.98 166.26 ;
      RECT 81.62 165.12 81.82 165.24 ;
      RECT 75.86 165.12 76.06 165.24 ;
      RECT 77.3 164.88 77.5 165 ;
      RECT 80.54 163.86 80.74 163.98 ;
      RECT 78.38 163.86 78.58 163.98 ;
      RECT 76.22 163.86 76.42 163.98 ;
      RECT 75.5 163.86 75.7 163.98 ;
      RECT 80.54 168.9 80.74 169.02 ;
      RECT 78.38 168.9 78.58 169.02 ;
      RECT 76.94 168.9 77.14 169.02 ;
      RECT 76.22 168.9 76.42 169.02 ;
      RECT 74.78 168.66 74.98 168.78 ;
      RECT 75.5 168.66 75.7 168.78 ;
      RECT 77.66 168.66 77.86 168.78 ;
      RECT 81.26 168.66 81.46 168.78 ;
      RECT 81.62 167.64 81.82 167.76 ;
      RECT 77.3 167.64 77.5 167.76 ;
      RECT 75.86 167.4 76.06 167.52 ;
      RECT 80.54 171.42 80.74 171.54 ;
      RECT 77.66 171.42 77.86 171.54 ;
      RECT 76.22 171.42 76.42 171.54 ;
      RECT 75.5 171.42 75.7 171.54 ;
      RECT 81.26 171.18 81.46 171.3 ;
      RECT 78.38 171.18 78.58 171.3 ;
      RECT 76.94 171.18 77.14 171.3 ;
      RECT 74.78 171.18 74.98 171.3 ;
      RECT 81.62 170.16 81.82 170.28 ;
      RECT 77.3 170.16 77.5 170.28 ;
      RECT 75.86 169.92 76.06 170.04 ;
      RECT 80.54 173.94 80.74 174.06 ;
      RECT 78.38 173.94 78.58 174.06 ;
      RECT 74.78 173.94 74.98 174.06 ;
      RECT 75.5 173.7 75.7 173.82 ;
      RECT 76.22 173.7 76.42 173.82 ;
      RECT 81.26 173.7 81.46 173.82 ;
      RECT 77.66 173.7 77.86 173.82 ;
      RECT 78.38 131.578 78.58 131.698 ;
      RECT 74.78 131.1 74.98 131.22 ;
      RECT 77.66 131.1 77.86 131.22 ;
      RECT 76.22 136.14 76.42 136.26 ;
      RECT 77.66 136.14 77.86 136.26 ;
      RECT 81.26 136.14 81.46 136.26 ;
      RECT 80.54 135.9 80.74 136.02 ;
      RECT 78.38 135.9 78.58 136.02 ;
      RECT 76.94 135.9 77.14 136.02 ;
      RECT 75.5 135.9 75.7 136.02 ;
      RECT 74.78 135.9 74.98 136.02 ;
      RECT 81.62 134.64 81.82 134.76 ;
      RECT 77.3 134.64 77.5 134.76 ;
      RECT 75.86 134.64 76.06 134.76 ;
      RECT 74.78 134.098 74.98 134.218 ;
      RECT 75.5 134.098 75.7 134.218 ;
      RECT 76.22 134.098 76.42 134.218 ;
      RECT 76.94 134.098 77.14 134.218 ;
      RECT 77.66 134.098 77.86 134.218 ;
      RECT 78.38 134.098 78.58 134.218 ;
      RECT 80.54 134.098 80.74 134.218 ;
      RECT 81.26 134.098 81.46 134.218 ;
      RECT 74.78 139.138 74.98 139.258 ;
      RECT 75.5 139.138 75.7 139.258 ;
      RECT 76.22 139.138 76.42 139.258 ;
      RECT 76.94 139.138 77.14 139.258 ;
      RECT 77.66 139.138 77.86 139.258 ;
      RECT 78.38 139.138 78.58 139.258 ;
      RECT 80.54 139.138 80.74 139.258 ;
      RECT 81.26 139.138 81.46 139.258 ;
      RECT 81.26 138.66 81.46 138.78 ;
      RECT 77.66 138.66 77.86 138.78 ;
      RECT 76.22 138.66 76.42 138.78 ;
      RECT 74.78 138.66 74.98 138.78 ;
      RECT 80.54 138.42 80.74 138.54 ;
      RECT 78.38 138.42 78.58 138.54 ;
      RECT 76.94 138.42 77.14 138.54 ;
      RECT 75.5 138.42 75.7 138.54 ;
      RECT 75.86 137.4 76.06 137.52 ;
      RECT 77.3 137.16 77.5 137.28 ;
      RECT 81.62 137.16 81.82 137.28 ;
      RECT 74.78 136.618 74.98 136.738 ;
      RECT 75.5 136.618 75.7 136.738 ;
      RECT 76.22 136.618 76.42 136.738 ;
      RECT 76.94 136.618 77.14 136.738 ;
      RECT 77.66 136.618 77.86 136.738 ;
      RECT 78.38 136.618 78.58 136.738 ;
      RECT 80.54 136.618 80.74 136.738 ;
      RECT 81.26 136.618 81.46 136.738 ;
      RECT 81.26 141.18 81.46 141.3 ;
      RECT 77.66 141.18 77.86 141.3 ;
      RECT 76.22 141.18 76.42 141.3 ;
      RECT 74.78 140.94 74.98 141.06 ;
      RECT 75.5 140.94 75.7 141.06 ;
      RECT 76.94 140.94 77.14 141.06 ;
      RECT 78.38 140.94 78.58 141.06 ;
      RECT 80.54 140.94 80.74 141.06 ;
      RECT 75.86 139.92 76.06 140.04 ;
      RECT 81.62 139.68 81.82 139.8 ;
      RECT 77.3 139.68 77.5 139.8 ;
      RECT 81.26 143.7 81.46 143.82 ;
      RECT 77.66 143.7 77.86 143.82 ;
      RECT 76.22 143.7 76.42 143.82 ;
      RECT 80.54 143.46 80.74 143.58 ;
      RECT 78.38 143.46 78.58 143.58 ;
      RECT 76.94 143.46 77.14 143.58 ;
      RECT 75.5 143.46 75.7 143.58 ;
      RECT 74.78 143.46 74.98 143.58 ;
      RECT 81.62 142.44 81.82 142.56 ;
      RECT 75.86 142.44 76.06 142.56 ;
      RECT 77.3 142.2 77.5 142.32 ;
      RECT 74.78 145.98 74.98 146.1 ;
      RECT 75.5 145.98 75.7 146.1 ;
      RECT 76.22 145.98 76.42 146.1 ;
      RECT 76.94 145.98 77.14 146.1 ;
      RECT 77.66 145.98 77.86 146.1 ;
      RECT 78.38 145.98 78.58 146.1 ;
      RECT 80.54 145.98 80.74 146.1 ;
      RECT 81.26 145.98 81.46 146.1 ;
      RECT 75.86 144.96 76.06 145.08 ;
      RECT 77.3 144.72 77.5 144.84 ;
      RECT 81.62 144.72 81.82 144.84 ;
      RECT 81.62 150 81.82 150.12 ;
      RECT 75.86 150 76.06 150.12 ;
      RECT 77.3 149.76 77.5 149.88 ;
      RECT 81.26 148.74 81.46 148.86 ;
      RECT 80.54 148.74 80.74 148.86 ;
      RECT 78.38 148.74 78.58 148.86 ;
      RECT 77.66 148.74 77.86 148.86 ;
      RECT 76.94 148.74 77.14 148.86 ;
      RECT 74.78 148.5 74.98 148.62 ;
      RECT 75.5 148.5 75.7 148.62 ;
      RECT 76.22 148.5 76.42 148.62 ;
      RECT 81.62 152.28 81.82 152.4 ;
      RECT 77.3 152.28 77.5 152.4 ;
      RECT 75.86 152.28 76.06 152.4 ;
      RECT 74.78 151.26 74.98 151.38 ;
      RECT 76.22 151.26 76.42 151.38 ;
      RECT 78.38 151.26 78.58 151.38 ;
      RECT 80.54 151.26 80.74 151.38 ;
      RECT 81.26 151.26 81.46 151.38 ;
      RECT 77.66 151.02 77.86 151.14 ;
      RECT 66.5 265.68 66.7 265.8 ;
      RECT 71.9 269.7 72.1 269.82 ;
      RECT 71.18 269.7 71.38 269.82 ;
      RECT 70.46 269.7 70.66 269.82 ;
      RECT 69.74 269.7 69.94 269.82 ;
      RECT 69.02 269.7 69.22 269.82 ;
      RECT 72.62 269.46 72.82 269.58 ;
      RECT 72.26 268.44 72.46 268.56 ;
      RECT 69.38 268.44 69.58 268.56 ;
      RECT 70.82 268.2 71.02 268.32 ;
      RECT 66.86 269.46 67.06 269.58 ;
      RECT 66.14 269.46 66.34 269.58 ;
      RECT 66.5 268.2 66.7 268.32 ;
      RECT 71.9 272.22 72.1 272.34 ;
      RECT 69.02 272.22 69.22 272.34 ;
      RECT 72.62 271.98 72.82 272.1 ;
      RECT 71.18 271.98 71.38 272.1 ;
      RECT 70.46 271.98 70.66 272.1 ;
      RECT 69.74 271.98 69.94 272.1 ;
      RECT 70.82 270.96 71.02 271.08 ;
      RECT 72.26 270.72 72.46 270.84 ;
      RECT 69.38 270.72 69.58 270.84 ;
      RECT 66.5 270.96 66.7 271.08 ;
      RECT 66.86 271.98 67.06 272.1 ;
      RECT 66.14 271.98 66.34 272.1 ;
      RECT 70.82 275.76 71.02 275.88 ;
      RECT 72.62 274.74 72.82 274.86 ;
      RECT 70.46 274.74 70.66 274.86 ;
      RECT 69.02 274.74 69.22 274.86 ;
      RECT 71.9 274.5 72.1 274.62 ;
      RECT 71.18 274.5 71.38 274.62 ;
      RECT 69.74 274.5 69.94 274.62 ;
      RECT 72.26 273.48 72.46 273.6 ;
      RECT 70.82 273.48 71.02 273.6 ;
      RECT 69.38 273.24 69.58 273.36 ;
      RECT 66.5 275.76 66.7 275.88 ;
      RECT 66.86 274.74 67.06 274.86 ;
      RECT 66.14 274.5 66.34 274.62 ;
      RECT 66.5 273.48 66.7 273.6 ;
      RECT 70.82 278.28 71.02 278.4 ;
      RECT 71.9 277.26 72.1 277.38 ;
      RECT 70.46 277.26 70.66 277.38 ;
      RECT 69.74 277.26 69.94 277.38 ;
      RECT 69.02 277.26 69.22 277.38 ;
      RECT 72.62 277.02 72.82 277.14 ;
      RECT 71.18 277.02 71.38 277.14 ;
      RECT 72.26 276 72.46 276.12 ;
      RECT 69.38 276 69.58 276.12 ;
      RECT 66.14 277.26 66.34 277.38 ;
      RECT 66.86 277.02 67.06 277.14 ;
      RECT 72.26 278.52 72.46 278.64 ;
      RECT 69.38 278.52 69.58 278.64 ;
      RECT 66.5 278.52 66.7 278.64 ;
      RECT 66.86 308.496 67.06 308.616 ;
      RECT 66.14 308.496 66.34 308.616 ;
      RECT 71.9 308.496 72.1 308.616 ;
      RECT 71.18 308.496 71.38 308.616 ;
      RECT 70.46 308.496 70.66 308.616 ;
      RECT 69.74 308.496 69.94 308.616 ;
      RECT 69.02 308.496 69.22 308.616 ;
      RECT 72.62 308.496 72.82 308.616 ;
      RECT 65.78 323.3835 65.98 323.5035 ;
      RECT 70.1 323.3835 70.3 323.5035 ;
      RECT 71.54 323.3835 71.74 323.5035 ;
      RECT 66.14 325.9425 66.34 326.0625 ;
      RECT 66.86 325.9425 67.06 326.0625 ;
      RECT 69.02 325.9425 69.22 326.0625 ;
      RECT 69.74 325.9425 69.94 326.0625 ;
      RECT 70.46 325.9425 70.66 326.0625 ;
      RECT 71.18 325.9425 71.38 326.0625 ;
      RECT 71.9 325.9425 72.1 326.0625 ;
      RECT 72.62 325.9425 72.82 326.0625 ;
      RECT 65.78 348.339 65.98 348.459 ;
      RECT 70.1 348.339 70.3 348.459 ;
      RECT 71.54 348.339 71.74 348.459 ;
      RECT 81.26 118.5 81.46 118.62 ;
      RECT 77.66 118.5 77.86 118.62 ;
      RECT 76.22 118.5 76.42 118.62 ;
      RECT 80.54 118.26 80.74 118.38 ;
      RECT 78.38 118.26 78.58 118.38 ;
      RECT 76.94 118.26 77.14 118.38 ;
      RECT 75.5 118.26 75.7 118.38 ;
      RECT 74.78 118.26 74.98 118.38 ;
      RECT 75.5 130.86 75.7 130.98 ;
      RECT 76.22 130.86 76.42 130.98 ;
      RECT 78.38 130.86 78.58 130.98 ;
      RECT 76.94 130.86 77.14 130.98 ;
      RECT 74.78 133.62 74.98 133.74 ;
      RECT 78.38 133.38 78.58 133.5 ;
      RECT 80.54 133.38 80.74 133.5 ;
      RECT 81.26 133.38 81.46 133.5 ;
      RECT 77.66 133.38 77.86 133.5 ;
      RECT 76.94 133.38 77.14 133.5 ;
      RECT 76.22 133.38 76.42 133.5 ;
      RECT 75.5 133.38 75.7 133.5 ;
      RECT 77.3 132.12 77.5 132.24 ;
      RECT 75.86 132.12 76.06 132.24 ;
      RECT 74.78 131.578 74.98 131.698 ;
      RECT 75.5 131.578 75.7 131.698 ;
      RECT 76.22 131.578 76.42 131.698 ;
      RECT 76.94 131.578 77.14 131.698 ;
      RECT 77.66 131.578 77.86 131.698 ;
      RECT 71.9 247.02 72.1 247.14 ;
      RECT 71.18 247.02 71.38 247.14 ;
      RECT 69.02 247.02 69.22 247.14 ;
      RECT 72.62 246.78 72.82 246.9 ;
      RECT 70.46 246.78 70.66 246.9 ;
      RECT 69.74 246.78 69.94 246.9 ;
      RECT 66.5 248.28 66.7 248.4 ;
      RECT 66.14 247.02 66.34 247.14 ;
      RECT 66.86 246.78 67.06 246.9 ;
      RECT 70.82 245.76 71.02 245.88 ;
      RECT 66.5 245.76 66.7 245.88 ;
      RECT 72.26 250.8 72.46 250.92 ;
      RECT 70.82 250.8 71.02 250.92 ;
      RECT 69.38 250.56 69.58 250.68 ;
      RECT 71.9 249.54 72.1 249.66 ;
      RECT 69.74 249.54 69.94 249.66 ;
      RECT 72.62 249.3 72.82 249.42 ;
      RECT 71.18 249.3 71.38 249.42 ;
      RECT 70.46 249.3 70.66 249.42 ;
      RECT 69.02 249.3 69.22 249.42 ;
      RECT 66.5 250.8 66.7 250.92 ;
      RECT 66.86 249.54 67.06 249.66 ;
      RECT 66.14 249.3 66.34 249.42 ;
      RECT 70.82 253.32 71.02 253.44 ;
      RECT 72.26 253.08 72.46 253.2 ;
      RECT 69.38 253.08 69.58 253.2 ;
      RECT 71.9 252.06 72.1 252.18 ;
      RECT 70.46 252.06 70.66 252.18 ;
      RECT 69.02 252.06 69.22 252.18 ;
      RECT 72.62 251.82 72.82 251.94 ;
      RECT 71.18 251.82 71.38 251.94 ;
      RECT 69.74 251.82 69.94 251.94 ;
      RECT 66.5 253.32 66.7 253.44 ;
      RECT 66.14 252.06 66.34 252.18 ;
      RECT 66.86 251.82 67.06 251.94 ;
      RECT 69.38 255.84 69.58 255.96 ;
      RECT 72.26 255.84 72.46 255.96 ;
      RECT 70.82 255.84 71.02 255.96 ;
      RECT 70.46 254.58 70.66 254.7 ;
      RECT 69.02 254.58 69.22 254.7 ;
      RECT 72.62 254.58 72.82 254.7 ;
      RECT 71.9 254.58 72.1 254.7 ;
      RECT 71.18 254.58 71.38 254.7 ;
      RECT 69.74 254.34 69.94 254.46 ;
      RECT 66.5 255.6 66.7 255.72 ;
      RECT 66.86 254.34 67.06 254.46 ;
      RECT 66.14 254.34 66.34 254.46 ;
      RECT 72.62 259.38 72.82 259.5 ;
      RECT 70.46 259.38 70.66 259.5 ;
      RECT 69.02 259.38 69.22 259.5 ;
      RECT 69.38 258.36 69.58 258.48 ;
      RECT 72.26 258.12 72.46 258.24 ;
      RECT 70.82 258.12 71.02 258.24 ;
      RECT 72.62 257.1 72.82 257.22 ;
      RECT 70.46 257.1 70.66 257.22 ;
      RECT 69.02 257.1 69.22 257.22 ;
      RECT 71.9 256.86 72.1 256.98 ;
      RECT 71.18 256.86 71.38 256.98 ;
      RECT 69.74 256.86 69.94 256.98 ;
      RECT 66.14 259.38 66.34 259.5 ;
      RECT 66.5 258.36 66.7 258.48 ;
      RECT 66.86 257.1 67.06 257.22 ;
      RECT 66.14 256.86 66.34 256.98 ;
      RECT 71.9 261.9 72.1 262.02 ;
      RECT 71.18 261.9 71.38 262.02 ;
      RECT 69.02 261.9 69.22 262.02 ;
      RECT 72.26 260.88 72.46 261 ;
      RECT 70.82 260.88 71.02 261 ;
      RECT 69.38 260.64 69.58 260.76 ;
      RECT 71.9 259.62 72.1 259.74 ;
      RECT 71.18 259.62 71.38 259.74 ;
      RECT 69.74 259.62 69.94 259.74 ;
      RECT 66.14 261.9 66.34 262.02 ;
      RECT 66.5 260.88 66.7 261 ;
      RECT 66.86 259.62 67.06 259.74 ;
      RECT 72.62 264.66 72.82 264.78 ;
      RECT 71.9 264.66 72.1 264.78 ;
      RECT 69.74 264.66 69.94 264.78 ;
      RECT 71.18 264.42 71.38 264.54 ;
      RECT 70.46 264.42 70.66 264.54 ;
      RECT 69.02 264.42 69.22 264.54 ;
      RECT 72.26 263.16 72.46 263.28 ;
      RECT 70.82 263.16 71.02 263.28 ;
      RECT 69.38 263.16 69.58 263.28 ;
      RECT 72.62 262.14 72.82 262.26 ;
      RECT 70.46 262.14 70.66 262.26 ;
      RECT 69.74 262.14 69.94 262.26 ;
      RECT 66.86 264.66 67.06 264.78 ;
      RECT 66.14 264.66 66.34 264.78 ;
      RECT 66.5 263.16 66.7 263.28 ;
      RECT 66.86 262.14 67.06 262.26 ;
      RECT 72.62 267.18 72.82 267.3 ;
      RECT 71.9 267.18 72.1 267.3 ;
      RECT 71.18 267.18 71.38 267.3 ;
      RECT 69.74 267.18 69.94 267.3 ;
      RECT 69.02 267.18 69.22 267.3 ;
      RECT 70.46 266.94 70.66 267.06 ;
      RECT 72.26 265.92 72.46 266.04 ;
      RECT 69.38 265.92 69.58 266.04 ;
      RECT 70.82 265.68 71.02 265.8 ;
      RECT 66.86 267.18 67.06 267.3 ;
      RECT 66.14 267.18 66.34 267.3 ;
      RECT 69.74 223.558 69.94 223.678 ;
      RECT 72.62 223.558 72.82 223.678 ;
      RECT 71.54 223.08 71.74 223.2 ;
      RECT 70.1 222.84 70.3 222.96 ;
      RECT 72.26 222.362 72.46 222.482 ;
      RECT 69.38 222.122 69.58 222.242 ;
      RECT 70.82 222.122 71.02 222.242 ;
      RECT 69.38 221.278 69.58 221.398 ;
      RECT 66.14 223.798 66.34 223.918 ;
      RECT 66.86 223.558 67.06 223.678 ;
      RECT 65.78 223.08 65.98 223.2 ;
      RECT 66.5 222.122 66.7 222.242 ;
      RECT 66.5 221.278 66.7 221.398 ;
      RECT 69.02 229.14 69.22 229.26 ;
      RECT 71.18 229.14 71.38 229.26 ;
      RECT 71.9 229.14 72.1 229.26 ;
      RECT 70.82 228.12 71.02 228.24 ;
      RECT 72.26 227.88 72.46 228 ;
      RECT 69.38 227.88 69.58 228 ;
      RECT 66.86 229.14 67.06 229.26 ;
      RECT 66.5 228.12 66.7 228.24 ;
      RECT 72.62 231.9 72.82 232.02 ;
      RECT 71.9 231.9 72.1 232.02 ;
      RECT 69.74 231.9 69.94 232.02 ;
      RECT 69.02 231.9 69.22 232.02 ;
      RECT 71.18 231.66 71.38 231.78 ;
      RECT 70.46 231.66 70.66 231.78 ;
      RECT 70.82 230.64 71.02 230.76 ;
      RECT 72.26 230.4 72.46 230.52 ;
      RECT 69.38 230.4 69.58 230.52 ;
      RECT 69.74 229.38 69.94 229.5 ;
      RECT 70.46 229.38 70.66 229.5 ;
      RECT 72.62 229.38 72.82 229.5 ;
      RECT 66.86 231.66 67.06 231.78 ;
      RECT 66.14 231.66 66.34 231.78 ;
      RECT 66.5 230.64 66.7 230.76 ;
      RECT 66.14 229.38 66.34 229.5 ;
      RECT 69.02 234.42 69.22 234.54 ;
      RECT 69.74 234.42 69.94 234.54 ;
      RECT 71.18 234.42 71.38 234.54 ;
      RECT 71.9 234.42 72.1 234.54 ;
      RECT 72.62 234.42 72.82 234.54 ;
      RECT 70.46 234.18 70.66 234.3 ;
      RECT 69.38 233.16 69.58 233.28 ;
      RECT 72.26 232.92 72.46 233.04 ;
      RECT 70.82 232.92 71.02 233.04 ;
      RECT 66.14 234.42 66.34 234.54 ;
      RECT 66.86 234.18 67.06 234.3 ;
      RECT 66.5 233.16 66.7 233.28 ;
      RECT 72.62 236.94 72.82 237.06 ;
      RECT 71.9 236.94 72.1 237.06 ;
      RECT 70.46 236.94 70.66 237.06 ;
      RECT 69.74 236.94 69.94 237.06 ;
      RECT 71.18 236.7 71.38 236.82 ;
      RECT 69.02 236.7 69.22 236.82 ;
      RECT 72.26 235.68 72.46 235.8 ;
      RECT 69.38 235.68 69.58 235.8 ;
      RECT 70.82 235.44 71.02 235.56 ;
      RECT 66.86 236.7 67.06 236.82 ;
      RECT 66.14 236.7 66.34 236.82 ;
      RECT 66.5 235.44 66.7 235.56 ;
      RECT 71.9 239.46 72.1 239.58 ;
      RECT 72.62 239.22 72.82 239.34 ;
      RECT 71.18 239.22 71.38 239.34 ;
      RECT 70.46 239.22 70.66 239.34 ;
      RECT 69.74 239.22 69.94 239.34 ;
      RECT 69.02 239.22 69.22 239.34 ;
      RECT 69.38 238.2 69.58 238.32 ;
      RECT 70.82 237.96 71.02 238.08 ;
      RECT 72.26 237.96 72.46 238.08 ;
      RECT 66.14 239.46 66.34 239.58 ;
      RECT 66.86 239.22 67.06 239.34 ;
      RECT 66.5 238.2 66.7 238.32 ;
      RECT 72.26 243 72.46 243.12 ;
      RECT 69.38 243 69.58 243.12 ;
      RECT 69.02 241.98 69.22 242.1 ;
      RECT 69.74 241.74 69.94 241.86 ;
      RECT 70.46 241.74 70.66 241.86 ;
      RECT 71.18 241.74 71.38 241.86 ;
      RECT 71.9 241.74 72.1 241.86 ;
      RECT 72.62 241.74 72.82 241.86 ;
      RECT 70.82 240.72 71.02 240.84 ;
      RECT 69.38 240.48 69.58 240.6 ;
      RECT 72.26 240.48 72.46 240.6 ;
      RECT 66.14 241.98 66.34 242.1 ;
      RECT 66.86 241.74 67.06 241.86 ;
      RECT 66.5 240.72 66.7 240.84 ;
      RECT 69.38 245.52 69.58 245.64 ;
      RECT 72.26 245.52 72.46 245.64 ;
      RECT 69.02 244.5 69.22 244.62 ;
      RECT 69.74 244.5 69.94 244.62 ;
      RECT 70.46 244.5 70.66 244.62 ;
      RECT 72.62 244.5 72.82 244.62 ;
      RECT 71.9 244.26 72.1 244.38 ;
      RECT 71.18 244.26 71.38 244.38 ;
      RECT 70.82 243.24 71.02 243.36 ;
      RECT 66.14 244.5 66.34 244.62 ;
      RECT 66.86 244.26 67.06 244.38 ;
      RECT 66.5 243.24 66.7 243.36 ;
      RECT 70.82 248.28 71.02 248.4 ;
      RECT 72.26 248.04 72.46 248.16 ;
      RECT 69.38 248.04 69.58 248.16 ;
      RECT 72.26 203.462 72.46 203.582 ;
      RECT 69.38 203.462 69.58 203.582 ;
      RECT 70.82 203.222 71.02 203.342 ;
      RECT 71.54 202.92 71.74 203.04 ;
      RECT 70.1 202.92 70.3 203.04 ;
      RECT 65.78 202.92 65.98 203.04 ;
      RECT 66.5 203.222 66.7 203.342 ;
      RECT 66.14 203.94 66.34 204.06 ;
      RECT 66.86 204.18 67.06 204.3 ;
      RECT 70.46 206.7 70.66 206.82 ;
      RECT 69.02 206.7 69.22 206.82 ;
      RECT 72.62 206.46 72.82 206.58 ;
      RECT 71.9 206.46 72.1 206.58 ;
      RECT 71.18 206.46 71.38 206.58 ;
      RECT 69.74 206.46 69.94 206.58 ;
      RECT 70.82 205.982 71.02 206.102 ;
      RECT 69.38 205.982 69.58 206.102 ;
      RECT 72.26 205.742 72.46 205.862 ;
      RECT 71.54 205.2 71.74 205.32 ;
      RECT 70.1 205.2 70.3 205.32 ;
      RECT 65.78 205.44 65.98 205.56 ;
      RECT 66.5 205.742 66.7 205.862 ;
      RECT 66.14 206.7 66.34 206.82 ;
      RECT 66.86 206.7 67.06 206.82 ;
      RECT 70.1 210.24 70.3 210.36 ;
      RECT 71.9 209.22 72.1 209.34 ;
      RECT 70.46 209.22 70.66 209.34 ;
      RECT 69.74 209.22 69.94 209.34 ;
      RECT 69.02 209.22 69.22 209.34 ;
      RECT 71.18 208.98 71.38 209.1 ;
      RECT 72.62 208.98 72.82 209.1 ;
      RECT 70.82 208.502 71.02 208.622 ;
      RECT 69.38 208.262 69.58 208.382 ;
      RECT 72.26 208.262 72.46 208.382 ;
      RECT 71.54 207.96 71.74 208.08 ;
      RECT 70.1 207.72 70.3 207.84 ;
      RECT 65.78 207.72 65.98 207.84 ;
      RECT 66.5 208.502 66.7 208.622 ;
      RECT 66.14 208.98 66.34 209.1 ;
      RECT 66.86 209.22 67.06 209.34 ;
      RECT 65.78 210.24 65.98 210.36 ;
      RECT 71.54 212.76 71.74 212.88 ;
      RECT 71.9 211.74 72.1 211.86 ;
      RECT 71.18 211.74 71.38 211.86 ;
      RECT 70.46 211.74 70.66 211.86 ;
      RECT 69.02 211.5 69.22 211.62 ;
      RECT 69.74 211.5 69.94 211.62 ;
      RECT 72.62 211.5 72.82 211.62 ;
      RECT 70.82 211.198 71.02 211.318 ;
      RECT 69.38 210.958 69.58 211.078 ;
      RECT 72.26 210.958 72.46 211.078 ;
      RECT 71.54 210.48 71.74 210.6 ;
      RECT 66.5 211.198 66.7 211.318 ;
      RECT 66.86 211.5 67.06 211.62 ;
      RECT 66.14 211.74 66.34 211.86 ;
      RECT 71.54 215.52 71.74 215.64 ;
      RECT 70.1 215.52 70.3 215.64 ;
      RECT 71.9 214.26 72.1 214.38 ;
      RECT 69.02 214.26 69.22 214.38 ;
      RECT 72.62 214.02 72.82 214.14 ;
      RECT 71.18 214.02 71.38 214.14 ;
      RECT 70.46 214.02 70.66 214.14 ;
      RECT 69.74 214.02 69.94 214.14 ;
      RECT 72.26 213.718 72.46 213.838 ;
      RECT 69.38 213.478 69.58 213.598 ;
      RECT 70.82 213.478 71.02 213.598 ;
      RECT 70.1 213 70.3 213.12 ;
      RECT 65.78 213 65.98 213.12 ;
      RECT 66.5 213.478 66.7 213.598 ;
      RECT 66.86 214.02 67.06 214.14 ;
      RECT 66.14 214.26 66.34 214.38 ;
      RECT 65.78 215.28 65.98 215.4 ;
      RECT 72.62 216.78 72.82 216.9 ;
      RECT 71.9 216.78 72.1 216.9 ;
      RECT 70.46 216.78 70.66 216.9 ;
      RECT 69.02 216.78 69.22 216.9 ;
      RECT 71.18 216.54 71.38 216.66 ;
      RECT 69.74 216.54 69.94 216.66 ;
      RECT 72.26 216.238 72.46 216.358 ;
      RECT 69.38 216.238 69.58 216.358 ;
      RECT 70.82 215.998 71.02 216.118 ;
      RECT 66.5 215.998 66.7 216.118 ;
      RECT 66.14 216.54 66.34 216.66 ;
      RECT 66.86 216.54 67.06 216.66 ;
      RECT 70.82 221.038 71.02 221.158 ;
      RECT 72.26 221.038 72.46 221.158 ;
      RECT 71.9 219.3 72.1 219.42 ;
      RECT 70.46 219.3 70.66 219.42 ;
      RECT 69.02 219.3 69.22 219.42 ;
      RECT 71.18 219.06 71.38 219.18 ;
      RECT 72.62 219.06 72.82 219.18 ;
      RECT 69.74 219.06 69.94 219.18 ;
      RECT 70.82 218.758 71.02 218.878 ;
      RECT 69.38 218.518 69.58 218.638 ;
      RECT 72.26 218.518 72.46 218.638 ;
      RECT 66.5 218.518 66.7 218.638 ;
      RECT 66.14 219.06 66.34 219.18 ;
      RECT 66.86 219.3 67.06 219.42 ;
      RECT 69.02 223.798 69.22 223.918 ;
      RECT 70.46 223.798 70.66 223.918 ;
      RECT 71.18 223.798 71.38 223.918 ;
      RECT 71.9 223.798 72.1 223.918 ;
      RECT 69.74 186.3 69.94 186.42 ;
      RECT 71.9 186.3 72.1 186.42 ;
      RECT 65.78 187.56 65.98 187.68 ;
      RECT 66.14 186.3 66.34 186.42 ;
      RECT 66.86 186.3 67.06 186.42 ;
      RECT 69.38 190.862 69.58 190.982 ;
      RECT 70.82 190.622 71.02 190.742 ;
      RECT 72.26 190.622 72.46 190.742 ;
      RECT 70.1 190.08 70.3 190.2 ;
      RECT 71.54 190.08 71.74 190.2 ;
      RECT 69.02 189.06 69.22 189.18 ;
      RECT 70.46 189.06 70.66 189.18 ;
      RECT 72.62 189.06 72.82 189.18 ;
      RECT 71.9 188.82 72.1 188.94 ;
      RECT 71.18 188.82 71.38 188.94 ;
      RECT 69.74 188.82 69.94 188.94 ;
      RECT 66.5 190.622 66.7 190.742 ;
      RECT 65.78 190.32 65.98 190.44 ;
      RECT 66.86 188.82 67.06 188.94 ;
      RECT 66.14 188.82 66.34 188.94 ;
      RECT 70.46 193.86 70.66 193.98 ;
      RECT 71.18 193.86 71.38 193.98 ;
      RECT 71.9 193.86 72.1 193.98 ;
      RECT 69.38 193.382 69.58 193.502 ;
      RECT 72.26 193.382 72.46 193.502 ;
      RECT 70.82 193.142 71.02 193.262 ;
      RECT 71.54 192.84 71.74 192.96 ;
      RECT 70.1 192.6 70.3 192.72 ;
      RECT 70.82 192.122 71.02 192.242 ;
      RECT 72.26 192.122 72.46 192.242 ;
      RECT 69.38 191.882 69.58 192.002 ;
      RECT 71.9 191.58 72.1 191.7 ;
      RECT 71.18 191.58 71.38 191.7 ;
      RECT 69.02 191.34 69.22 191.46 ;
      RECT 69.74 191.34 69.94 191.46 ;
      RECT 70.46 191.34 70.66 191.46 ;
      RECT 72.62 191.34 72.82 191.46 ;
      RECT 66.86 193.86 67.06 193.98 ;
      RECT 66.5 193.142 66.7 193.262 ;
      RECT 65.78 192.6 65.98 192.72 ;
      RECT 66.5 191.882 66.7 192.002 ;
      RECT 66.86 191.58 67.06 191.7 ;
      RECT 66.14 191.34 66.34 191.46 ;
      RECT 70.82 194.642 71.02 194.762 ;
      RECT 72.26 194.402 72.46 194.522 ;
      RECT 69.38 194.402 69.58 194.522 ;
      RECT 72.62 194.1 72.82 194.22 ;
      RECT 69.74 194.1 69.94 194.22 ;
      RECT 69.02 194.1 69.22 194.22 ;
      RECT 66.5 194.642 66.7 194.762 ;
      RECT 66.14 194.1 66.34 194.22 ;
      RECT 65.78 195.36 65.98 195.48 ;
      RECT 66.5 195.902 66.7 196.022 ;
      RECT 66.14 196.38 66.34 196.5 ;
      RECT 71.54 195.12 71.74 195.24 ;
      RECT 70.1 195.36 70.3 195.48 ;
      RECT 69.38 195.662 69.58 195.782 ;
      RECT 70.82 195.662 71.02 195.782 ;
      RECT 72.26 195.902 72.46 196.022 ;
      RECT 71.9 196.38 72.1 196.5 ;
      RECT 70.46 196.38 70.66 196.5 ;
      RECT 69.02 196.38 69.22 196.5 ;
      RECT 69.74 199.14 69.94 199.26 ;
      RECT 71.18 199.14 71.38 199.26 ;
      RECT 71.9 199.14 72.1 199.26 ;
      RECT 66.86 196.62 67.06 196.74 ;
      RECT 65.78 197.88 65.98 198 ;
      RECT 66.5 198.182 66.7 198.302 ;
      RECT 66.86 199.14 67.06 199.26 ;
      RECT 66.14 199.14 66.34 199.26 ;
      RECT 69.74 196.62 69.94 196.74 ;
      RECT 71.18 196.62 71.38 196.74 ;
      RECT 72.62 196.62 72.82 196.74 ;
      RECT 71.54 197.64 71.74 197.76 ;
      RECT 70.1 197.88 70.3 198 ;
      RECT 72.26 198.182 72.46 198.302 ;
      RECT 69.38 198.182 69.58 198.302 ;
      RECT 70.82 198.422 71.02 198.542 ;
      RECT 69.02 198.9 69.22 199.02 ;
      RECT 70.46 198.9 70.66 199.02 ;
      RECT 72.62 199.14 72.82 199.26 ;
      RECT 69.74 201.66 69.94 201.78 ;
      RECT 71.18 201.66 71.38 201.78 ;
      RECT 72.62 201.66 72.82 201.78 ;
      RECT 69.02 201.66 69.22 201.78 ;
      RECT 70.46 201.42 70.66 201.54 ;
      RECT 71.9 201.42 72.1 201.54 ;
      RECT 69.38 200.942 69.58 201.062 ;
      RECT 70.82 200.942 71.02 201.062 ;
      RECT 72.26 200.702 72.46 200.822 ;
      RECT 71.54 200.4 71.74 200.52 ;
      RECT 70.1 200.16 70.3 200.28 ;
      RECT 65.78 200.16 65.98 200.28 ;
      RECT 66.5 200.702 66.7 200.822 ;
      RECT 66.14 201.66 66.34 201.78 ;
      RECT 66.86 201.66 67.06 201.78 ;
      RECT 69.02 204.18 69.22 204.3 ;
      RECT 69.74 204.18 69.94 204.3 ;
      RECT 70.46 204.18 70.66 204.3 ;
      RECT 71.18 204.18 71.38 204.3 ;
      RECT 72.62 203.94 72.82 204.06 ;
      RECT 71.9 203.94 72.1 204.06 ;
      RECT 71.9 161.1 72.1 161.22 ;
      RECT 72.62 161.1 72.82 161.22 ;
      RECT 66.14 166.38 66.34 166.5 ;
      RECT 66.86 166.14 67.06 166.26 ;
      RECT 65.78 164.88 65.98 165 ;
      RECT 71.9 166.38 72.1 166.5 ;
      RECT 70.46 166.38 70.66 166.5 ;
      RECT 69.74 166.38 69.94 166.5 ;
      RECT 69.02 166.38 69.22 166.5 ;
      RECT 72.62 166.14 72.82 166.26 ;
      RECT 71.18 166.14 71.38 166.26 ;
      RECT 71.54 165.12 71.74 165.24 ;
      RECT 70.1 164.88 70.3 165 ;
      RECT 72.62 163.86 72.82 163.98 ;
      RECT 69.74 163.86 69.94 163.98 ;
      RECT 69.02 163.86 69.22 163.98 ;
      RECT 66.14 168.9 66.34 169.02 ;
      RECT 66.86 168.66 67.06 168.78 ;
      RECT 65.78 167.4 65.98 167.52 ;
      RECT 72.62 168.9 72.82 169.02 ;
      RECT 71.18 168.9 71.38 169.02 ;
      RECT 69.74 168.9 69.94 169.02 ;
      RECT 69.02 168.66 69.22 168.78 ;
      RECT 70.46 168.66 70.66 168.78 ;
      RECT 71.9 168.66 72.1 168.78 ;
      RECT 71.54 167.64 71.74 167.76 ;
      RECT 70.1 167.4 70.3 167.52 ;
      RECT 72.62 171.42 72.82 171.54 ;
      RECT 71.9 171.42 72.1 171.54 ;
      RECT 69.02 171.42 69.22 171.54 ;
      RECT 71.18 171.18 71.38 171.3 ;
      RECT 70.46 171.18 70.66 171.3 ;
      RECT 69.74 171.18 69.94 171.3 ;
      RECT 71.54 170.16 71.74 170.28 ;
      RECT 70.1 169.92 70.3 170.04 ;
      RECT 66.14 171.42 66.34 171.54 ;
      RECT 66.86 171.18 67.06 171.3 ;
      RECT 65.78 170.16 65.98 170.28 ;
      RECT 72.62 173.94 72.82 174.06 ;
      RECT 71.18 173.94 71.38 174.06 ;
      RECT 69.74 173.94 69.94 174.06 ;
      RECT 69.02 173.7 69.22 173.82 ;
      RECT 70.46 173.7 70.66 173.82 ;
      RECT 71.9 173.7 72.1 173.82 ;
      RECT 71.54 172.68 71.74 172.8 ;
      RECT 70.1 172.44 70.3 172.56 ;
      RECT 66.86 173.94 67.06 174.06 ;
      RECT 66.14 173.7 66.34 173.82 ;
      RECT 65.78 172.68 65.98 172.8 ;
      RECT 71.54 177.48 71.74 177.6 ;
      RECT 71.18 176.46 71.38 176.58 ;
      RECT 70.46 176.46 70.66 176.58 ;
      RECT 72.62 176.22 72.82 176.34 ;
      RECT 71.9 176.22 72.1 176.34 ;
      RECT 69.74 176.22 69.94 176.34 ;
      RECT 69.02 176.22 69.22 176.34 ;
      RECT 71.54 175.2 71.74 175.32 ;
      RECT 70.1 174.96 70.3 175.08 ;
      RECT 66.86 176.46 67.06 176.58 ;
      RECT 66.14 176.46 66.34 176.58 ;
      RECT 65.78 175.2 65.98 175.32 ;
      RECT 71.54 180 71.74 180.12 ;
      RECT 72.62 178.98 72.82 179.1 ;
      RECT 69.74 178.98 69.94 179.1 ;
      RECT 71.9 178.74 72.1 178.86 ;
      RECT 71.18 178.74 71.38 178.86 ;
      RECT 70.46 178.74 70.66 178.86 ;
      RECT 69.02 178.74 69.22 178.86 ;
      RECT 70.1 177.72 70.3 177.84 ;
      RECT 65.78 180 65.98 180.12 ;
      RECT 66.86 178.98 67.06 179.1 ;
      RECT 66.14 178.98 66.34 179.1 ;
      RECT 65.78 177.72 65.98 177.84 ;
      RECT 71.54 182.76 71.74 182.88 ;
      RECT 70.1 182.52 70.3 182.64 ;
      RECT 69.02 181.5 69.22 181.62 ;
      RECT 70.46 181.5 70.66 181.62 ;
      RECT 72.62 181.5 72.82 181.62 ;
      RECT 71.9 181.26 72.1 181.38 ;
      RECT 71.18 181.26 71.38 181.38 ;
      RECT 69.74 181.26 69.94 181.38 ;
      RECT 70.1 180.24 70.3 180.36 ;
      RECT 65.78 182.52 65.98 182.64 ;
      RECT 66.14 181.5 66.34 181.62 ;
      RECT 66.86 181.5 67.06 181.62 ;
      RECT 71.54 185.28 71.74 185.4 ;
      RECT 70.1 185.04 70.3 185.16 ;
      RECT 69.74 184.02 69.94 184.14 ;
      RECT 70.46 184.02 70.66 184.14 ;
      RECT 69.02 184.02 69.22 184.14 ;
      RECT 71.9 183.78 72.1 183.9 ;
      RECT 72.62 183.78 72.82 183.9 ;
      RECT 71.18 183.78 71.38 183.9 ;
      RECT 65.78 185.28 65.98 185.4 ;
      RECT 66.14 184.02 66.34 184.14 ;
      RECT 66.86 183.78 67.06 183.9 ;
      RECT 71.54 187.8 71.74 187.92 ;
      RECT 70.1 187.8 70.3 187.92 ;
      RECT 69.02 186.54 69.22 186.66 ;
      RECT 70.46 186.54 70.66 186.66 ;
      RECT 71.18 186.54 71.38 186.66 ;
      RECT 72.62 186.54 72.82 186.66 ;
      RECT 71.9 140.94 72.1 141.06 ;
      RECT 70.1 139.92 70.3 140.04 ;
      RECT 71.54 139.68 71.74 139.8 ;
      RECT 66.86 143.7 67.06 143.82 ;
      RECT 72.62 143.7 72.82 143.82 ;
      RECT 71.18 143.7 71.38 143.82 ;
      RECT 66.14 143.46 66.34 143.58 ;
      RECT 65.78 142.2 65.98 142.32 ;
      RECT 71.9 143.46 72.1 143.58 ;
      RECT 70.46 143.46 70.66 143.58 ;
      RECT 69.74 143.46 69.94 143.58 ;
      RECT 69.02 143.46 69.22 143.58 ;
      RECT 71.54 142.44 71.74 142.56 ;
      RECT 70.1 142.2 70.3 142.32 ;
      RECT 66.14 145.98 66.34 146.1 ;
      RECT 66.86 145.98 67.06 146.1 ;
      RECT 65.78 144.96 65.98 145.08 ;
      RECT 69.02 145.98 69.22 146.1 ;
      RECT 69.74 145.98 69.94 146.1 ;
      RECT 70.46 145.98 70.66 146.1 ;
      RECT 71.18 145.98 71.38 146.1 ;
      RECT 71.9 145.98 72.1 146.1 ;
      RECT 72.62 145.98 72.82 146.1 ;
      RECT 70.1 144.72 70.3 144.84 ;
      RECT 71.54 144.72 71.74 144.84 ;
      RECT 65.78 149.76 65.98 149.88 ;
      RECT 66.14 148.74 66.34 148.86 ;
      RECT 66.86 148.5 67.06 148.62 ;
      RECT 70.1 150 70.3 150.12 ;
      RECT 71.54 149.76 71.74 149.88 ;
      RECT 71.9 148.74 72.1 148.86 ;
      RECT 70.46 148.74 70.66 148.86 ;
      RECT 69.74 148.74 69.94 148.86 ;
      RECT 69.02 148.74 69.22 148.86 ;
      RECT 71.18 148.5 71.38 148.62 ;
      RECT 72.62 148.5 72.82 148.62 ;
      RECT 65.78 152.28 65.98 152.4 ;
      RECT 66.86 151.26 67.06 151.38 ;
      RECT 66.14 151.02 66.34 151.14 ;
      RECT 70.1 152.52 70.3 152.64 ;
      RECT 71.54 152.28 71.74 152.4 ;
      RECT 70.46 151.26 70.66 151.38 ;
      RECT 71.18 151.26 71.38 151.38 ;
      RECT 72.62 151.02 72.82 151.14 ;
      RECT 71.9 151.02 72.1 151.14 ;
      RECT 69.74 151.02 69.94 151.14 ;
      RECT 69.02 151.02 69.22 151.14 ;
      RECT 65.78 154.8 65.98 154.92 ;
      RECT 66.14 153.54 66.34 153.66 ;
      RECT 66.86 153.54 67.06 153.66 ;
      RECT 70.1 155.04 70.3 155.16 ;
      RECT 71.54 154.8 71.74 154.92 ;
      RECT 72.62 153.78 72.82 153.9 ;
      RECT 71.18 153.78 71.38 153.9 ;
      RECT 69.74 153.78 69.94 153.9 ;
      RECT 69.02 153.54 69.22 153.66 ;
      RECT 70.46 153.54 70.66 153.66 ;
      RECT 71.9 153.54 72.1 153.66 ;
      RECT 66.5 158.278 66.7 158.398 ;
      RECT 65.78 157.56 65.98 157.68 ;
      RECT 66.5 156.842 66.7 156.962 ;
      RECT 66.14 156.3 66.34 156.42 ;
      RECT 66.86 156.3 67.06 156.42 ;
      RECT 70.82 158.278 71.02 158.398 ;
      RECT 72.26 158.038 72.46 158.158 ;
      RECT 69.38 158.038 69.58 158.158 ;
      RECT 70.1 157.56 70.3 157.68 ;
      RECT 71.54 157.32 71.74 157.44 ;
      RECT 70.82 156.842 71.02 156.962 ;
      RECT 72.26 156.602 72.46 156.722 ;
      RECT 69.38 156.602 69.58 156.722 ;
      RECT 69.74 156.3 69.94 156.42 ;
      RECT 71.9 156.3 72.1 156.42 ;
      RECT 72.62 156.06 72.82 156.18 ;
      RECT 71.18 156.06 71.38 156.18 ;
      RECT 70.46 156.06 70.66 156.18 ;
      RECT 69.02 156.06 69.22 156.18 ;
      RECT 65.78 159.84 65.98 159.96 ;
      RECT 66.14 158.82 66.34 158.94 ;
      RECT 66.86 158.82 67.06 158.94 ;
      RECT 70.1 160.08 70.3 160.2 ;
      RECT 71.54 160.08 71.74 160.2 ;
      RECT 70.46 158.82 70.66 158.94 ;
      RECT 71.9 158.82 72.1 158.94 ;
      RECT 69.02 158.58 69.22 158.7 ;
      RECT 69.74 158.58 69.94 158.7 ;
      RECT 71.18 158.58 71.38 158.7 ;
      RECT 72.62 158.58 72.82 158.7 ;
      RECT 66.14 163.62 66.34 163.74 ;
      RECT 66.86 163.62 67.06 163.74 ;
      RECT 65.78 162.36 65.98 162.48 ;
      RECT 66.14 161.1 66.34 161.22 ;
      RECT 66.86 161.1 67.06 161.22 ;
      RECT 70.46 163.62 70.66 163.74 ;
      RECT 71.18 163.62 71.38 163.74 ;
      RECT 71.9 163.62 72.1 163.74 ;
      RECT 70.1 162.6 70.3 162.72 ;
      RECT 71.54 162.36 71.74 162.48 ;
      RECT 69.02 161.1 69.22 161.22 ;
      RECT 69.74 161.1 69.94 161.22 ;
      RECT 70.46 161.1 70.66 161.22 ;
      RECT 71.18 161.1 71.38 161.22 ;
      RECT 71.18 125.82 71.38 125.94 ;
      RECT 72.62 125.82 72.82 125.94 ;
      RECT 66.86 130.86 67.06 130.98 ;
      RECT 65.78 129.6 65.98 129.72 ;
      RECT 66.14 129.058 66.34 129.178 ;
      RECT 66.86 129.058 67.06 129.178 ;
      RECT 66.14 128.58 66.34 128.7 ;
      RECT 66.86 128.58 67.06 128.7 ;
      RECT 69.74 130.86 69.94 130.98 ;
      RECT 71.18 130.86 71.38 130.98 ;
      RECT 72.62 130.86 72.82 130.98 ;
      RECT 70.1 129.84 70.3 129.96 ;
      RECT 71.54 129.6 71.74 129.72 ;
      RECT 69.02 129.058 69.22 129.178 ;
      RECT 69.74 129.058 69.94 129.178 ;
      RECT 70.46 129.058 70.66 129.178 ;
      RECT 71.18 129.058 71.38 129.178 ;
      RECT 71.9 129.058 72.1 129.178 ;
      RECT 72.62 129.058 72.82 129.178 ;
      RECT 71.9 128.58 72.1 128.7 ;
      RECT 70.46 128.58 70.66 128.7 ;
      RECT 72.62 128.34 72.82 128.46 ;
      RECT 71.18 128.34 71.38 128.46 ;
      RECT 69.74 128.34 69.94 128.46 ;
      RECT 69.02 128.34 69.22 128.46 ;
      RECT 66.14 133.62 66.34 133.74 ;
      RECT 66.86 133.38 67.06 133.5 ;
      RECT 65.78 132.36 65.98 132.48 ;
      RECT 66.14 131.578 66.34 131.698 ;
      RECT 66.86 131.578 67.06 131.698 ;
      RECT 66.14 131.1 66.34 131.22 ;
      RECT 71.18 133.62 71.38 133.74 ;
      RECT 69.74 133.62 69.94 133.74 ;
      RECT 69.02 133.62 69.22 133.74 ;
      RECT 72.62 133.38 72.82 133.5 ;
      RECT 71.9 133.38 72.1 133.5 ;
      RECT 70.46 133.38 70.66 133.5 ;
      RECT 70.1 132.36 70.3 132.48 ;
      RECT 71.54 132.12 71.74 132.24 ;
      RECT 69.02 131.578 69.22 131.698 ;
      RECT 69.74 131.578 69.94 131.698 ;
      RECT 70.46 131.578 70.66 131.698 ;
      RECT 71.18 131.578 71.38 131.698 ;
      RECT 71.9 131.578 72.1 131.698 ;
      RECT 72.62 131.578 72.82 131.698 ;
      RECT 71.9 131.1 72.1 131.22 ;
      RECT 70.46 131.1 70.66 131.22 ;
      RECT 69.02 131.1 69.22 131.22 ;
      RECT 66.86 135.9 67.06 136.02 ;
      RECT 66.14 135.9 66.34 136.02 ;
      RECT 65.78 134.64 65.98 134.76 ;
      RECT 66.14 134.098 66.34 134.218 ;
      RECT 66.86 134.098 67.06 134.218 ;
      RECT 69.74 136.14 69.94 136.26 ;
      RECT 71.9 136.14 72.1 136.26 ;
      RECT 72.62 135.9 72.82 136.02 ;
      RECT 71.18 135.9 71.38 136.02 ;
      RECT 70.46 135.9 70.66 136.02 ;
      RECT 69.02 135.9 69.22 136.02 ;
      RECT 70.1 134.88 70.3 135 ;
      RECT 71.54 134.64 71.74 134.76 ;
      RECT 69.02 134.098 69.22 134.218 ;
      RECT 69.74 134.098 69.94 134.218 ;
      RECT 70.46 134.098 70.66 134.218 ;
      RECT 71.18 134.098 71.38 134.218 ;
      RECT 71.9 134.098 72.1 134.218 ;
      RECT 72.62 134.098 72.82 134.218 ;
      RECT 66.14 139.138 66.34 139.258 ;
      RECT 66.86 139.138 67.06 139.258 ;
      RECT 66.86 138.66 67.06 138.78 ;
      RECT 66.14 138.42 66.34 138.54 ;
      RECT 65.78 137.16 65.98 137.28 ;
      RECT 66.14 136.618 66.34 136.738 ;
      RECT 66.86 136.618 67.06 136.738 ;
      RECT 69.02 139.138 69.22 139.258 ;
      RECT 69.74 139.138 69.94 139.258 ;
      RECT 70.46 139.138 70.66 139.258 ;
      RECT 71.18 139.138 71.38 139.258 ;
      RECT 71.9 139.138 72.1 139.258 ;
      RECT 72.62 139.138 72.82 139.258 ;
      RECT 69.74 138.66 69.94 138.78 ;
      RECT 69.02 138.66 69.22 138.78 ;
      RECT 72.62 138.42 72.82 138.54 ;
      RECT 71.9 138.42 72.1 138.54 ;
      RECT 71.18 138.42 71.38 138.54 ;
      RECT 70.46 138.42 70.66 138.54 ;
      RECT 70.1 137.4 70.3 137.52 ;
      RECT 71.54 137.16 71.74 137.28 ;
      RECT 69.02 136.618 69.22 136.738 ;
      RECT 69.74 136.618 69.94 136.738 ;
      RECT 70.46 136.618 70.66 136.738 ;
      RECT 71.18 136.618 71.38 136.738 ;
      RECT 71.9 136.618 72.1 136.738 ;
      RECT 72.62 136.618 72.82 136.738 ;
      RECT 66.14 140.94 66.34 141.06 ;
      RECT 66.86 140.94 67.06 141.06 ;
      RECT 65.78 139.68 65.98 139.8 ;
      RECT 72.62 141.18 72.82 141.3 ;
      RECT 71.18 141.18 71.38 141.3 ;
      RECT 69.74 141.18 69.94 141.3 ;
      RECT 69.02 140.94 69.22 141.06 ;
      RECT 70.46 140.94 70.66 141.06 ;
      RECT 57.5 283.087 57.7 283.207 ;
      RECT 58.58 305.498 58.78 305.618 ;
      RECT 63.98 308.496 64.18 308.616 ;
      RECT 63.26 308.496 63.46 308.616 ;
      RECT 61.1 308.496 61.3 308.616 ;
      RECT 60.38 308.496 60.58 308.616 ;
      RECT 65.42 308.496 65.62 308.616 ;
      RECT 64.7 308.496 64.9 308.616 ;
      RECT 59.66 305.967 59.86 306.087 ;
      RECT 58.94 305.967 59.14 306.087 ;
      RECT 58.22 305.967 58.42 306.087 ;
      RECT 57.5 305.967 57.7 306.087 ;
      RECT 64.34 323.3835 64.54 323.5035 ;
      RECT 60.02 323.3835 60.22 323.5035 ;
      RECT 58.58 323.3835 58.78 323.5035 ;
      RECT 65.42 325.9425 65.62 326.0625 ;
      RECT 64.7 325.9425 64.9 326.0625 ;
      RECT 63.98 325.9425 64.18 326.0625 ;
      RECT 63.26 325.9425 63.46 326.0625 ;
      RECT 61.1 325.9425 61.3 326.0625 ;
      RECT 60.38 325.9425 60.58 326.0625 ;
      RECT 57.5 325.9425 57.7 326.0625 ;
      RECT 58.22 325.9425 58.42 326.0625 ;
      RECT 58.94 325.9425 59.14 326.0625 ;
      RECT 59.66 325.9425 59.86 326.0625 ;
      RECT 58.58 348.339 58.78 348.459 ;
      RECT 64.34 348.339 64.54 348.459 ;
      RECT 60.02 348.339 60.22 348.459 ;
      RECT 65.78 119.52 65.98 119.64 ;
      RECT 66.14 118.978 66.34 119.098 ;
      RECT 66.86 118.978 67.06 119.098 ;
      RECT 66.86 118.26 67.06 118.38 ;
      RECT 66.14 118.26 66.34 118.38 ;
      RECT 70.1 119.76 70.3 119.88 ;
      RECT 71.54 119.52 71.74 119.64 ;
      RECT 69.02 118.978 69.22 119.098 ;
      RECT 69.74 118.978 69.94 119.098 ;
      RECT 70.46 118.978 70.66 119.098 ;
      RECT 71.18 118.978 71.38 119.098 ;
      RECT 71.9 118.978 72.1 119.098 ;
      RECT 72.62 118.978 72.82 119.098 ;
      RECT 71.9 118.5 72.1 118.62 ;
      RECT 70.46 118.5 70.66 118.62 ;
      RECT 72.62 118.26 72.82 118.38 ;
      RECT 71.18 118.26 71.38 118.38 ;
      RECT 69.74 118.26 69.94 118.38 ;
      RECT 69.02 118.26 69.22 118.38 ;
      RECT 65.78 122.04 65.98 122.16 ;
      RECT 66.14 121.498 66.34 121.618 ;
      RECT 66.86 121.498 67.06 121.618 ;
      RECT 66.14 121.02 66.34 121.14 ;
      RECT 66.86 120.78 67.06 120.9 ;
      RECT 70.1 122.28 70.3 122.4 ;
      RECT 71.54 122.04 71.74 122.16 ;
      RECT 69.02 121.498 69.22 121.618 ;
      RECT 69.74 121.498 69.94 121.618 ;
      RECT 70.46 121.498 70.66 121.618 ;
      RECT 71.18 121.498 71.38 121.618 ;
      RECT 71.9 121.498 72.1 121.618 ;
      RECT 72.62 121.498 72.82 121.618 ;
      RECT 69.02 121.02 69.22 121.14 ;
      RECT 71.18 121.02 71.38 121.14 ;
      RECT 70.46 120.78 70.66 120.9 ;
      RECT 71.9 120.78 72.1 120.9 ;
      RECT 72.62 120.78 72.82 120.9 ;
      RECT 69.74 120.78 69.94 120.9 ;
      RECT 65.78 124.56 65.98 124.68 ;
      RECT 66.14 124.018 66.34 124.138 ;
      RECT 66.86 124.018 67.06 124.138 ;
      RECT 66.14 123.54 66.34 123.66 ;
      RECT 66.86 123.3 67.06 123.42 ;
      RECT 70.1 124.8 70.3 124.92 ;
      RECT 71.54 124.56 71.74 124.68 ;
      RECT 69.02 124.018 69.22 124.138 ;
      RECT 69.74 124.018 69.94 124.138 ;
      RECT 70.46 124.018 70.66 124.138 ;
      RECT 71.18 124.018 71.38 124.138 ;
      RECT 71.9 124.018 72.1 124.138 ;
      RECT 72.62 124.018 72.82 124.138 ;
      RECT 69.02 123.54 69.22 123.66 ;
      RECT 71.18 123.54 71.38 123.66 ;
      RECT 69.74 123.3 69.94 123.42 ;
      RECT 70.46 123.3 70.66 123.42 ;
      RECT 71.9 123.3 72.1 123.42 ;
      RECT 72.62 123.3 72.82 123.42 ;
      RECT 65.78 127.08 65.98 127.2 ;
      RECT 66.14 126.538 66.34 126.658 ;
      RECT 66.86 126.538 67.06 126.658 ;
      RECT 66.14 125.82 66.34 125.94 ;
      RECT 66.86 125.82 67.06 125.94 ;
      RECT 70.1 127.32 70.3 127.44 ;
      RECT 71.54 127.08 71.74 127.2 ;
      RECT 69.02 126.538 69.22 126.658 ;
      RECT 69.74 126.538 69.94 126.658 ;
      RECT 70.46 126.538 70.66 126.658 ;
      RECT 71.18 126.538 71.38 126.658 ;
      RECT 71.9 126.538 72.1 126.658 ;
      RECT 72.62 126.538 72.82 126.658 ;
      RECT 69.02 126.06 69.22 126.18 ;
      RECT 70.46 126.06 70.66 126.18 ;
      RECT 71.9 126.06 72.1 126.18 ;
      RECT 69.74 125.82 69.94 125.94 ;
      RECT 65.06 235.44 65.26 235.56 ;
      RECT 64.7 239.46 64.9 239.58 ;
      RECT 63.98 239.46 64.18 239.58 ;
      RECT 63.26 239.46 63.46 239.58 ;
      RECT 65.42 239.22 65.62 239.34 ;
      RECT 63.62 238.2 63.82 238.32 ;
      RECT 65.06 237.96 65.26 238.08 ;
      RECT 65.06 243 65.26 243.12 ;
      RECT 63.98 241.98 64.18 242.1 ;
      RECT 64.7 241.98 64.9 242.1 ;
      RECT 63.26 241.74 63.46 241.86 ;
      RECT 65.42 241.74 65.62 241.86 ;
      RECT 63.62 240.72 63.82 240.84 ;
      RECT 65.06 240.48 65.26 240.6 ;
      RECT 65.06 245.52 65.26 245.64 ;
      RECT 65.42 244.5 65.62 244.62 ;
      RECT 63.98 244.5 64.18 244.62 ;
      RECT 64.7 244.26 64.9 244.38 ;
      RECT 63.26 244.26 63.46 244.38 ;
      RECT 63.62 243.24 63.82 243.36 ;
      RECT 63.62 248.28 63.82 248.4 ;
      RECT 65.06 248.04 65.26 248.16 ;
      RECT 65.42 247.02 65.62 247.14 ;
      RECT 64.7 247.02 64.9 247.14 ;
      RECT 63.98 247.02 64.18 247.14 ;
      RECT 63.26 246.78 63.46 246.9 ;
      RECT 63.62 245.76 63.82 245.88 ;
      RECT 65.06 250.8 65.26 250.92 ;
      RECT 63.62 250.8 63.82 250.92 ;
      RECT 65.42 249.54 65.62 249.66 ;
      RECT 64.7 249.54 64.9 249.66 ;
      RECT 63.98 249.54 64.18 249.66 ;
      RECT 63.26 249.3 63.46 249.42 ;
      RECT 63.62 253.32 63.82 253.44 ;
      RECT 65.06 253.08 65.26 253.2 ;
      RECT 64.7 252.06 64.9 252.18 ;
      RECT 63.98 252.06 64.18 252.18 ;
      RECT 65.42 251.82 65.62 251.94 ;
      RECT 63.26 251.82 63.46 251.94 ;
      RECT 65.06 255.84 65.26 255.96 ;
      RECT 63.62 255.6 63.82 255.72 ;
      RECT 65.42 254.58 65.62 254.7 ;
      RECT 64.7 254.34 64.9 254.46 ;
      RECT 63.98 254.34 64.18 254.46 ;
      RECT 63.26 254.34 63.46 254.46 ;
      RECT 64.7 259.38 64.9 259.5 ;
      RECT 63.26 259.38 63.46 259.5 ;
      RECT 63.62 258.36 63.82 258.48 ;
      RECT 65.06 258.12 65.26 258.24 ;
      RECT 65.42 257.1 65.62 257.22 ;
      RECT 64.7 257.1 64.9 257.22 ;
      RECT 63.98 257.1 64.18 257.22 ;
      RECT 63.26 256.86 63.46 256.98 ;
      RECT 63.62 260.88 63.82 261 ;
      RECT 65.06 260.64 65.26 260.76 ;
      RECT 65.42 259.62 65.62 259.74 ;
      RECT 63.98 259.62 64.18 259.74 ;
      RECT 64.7 264.66 64.9 264.78 ;
      RECT 65.42 264.42 65.62 264.54 ;
      RECT 63.98 264.42 64.18 264.54 ;
      RECT 63.26 264.42 63.46 264.54 ;
      RECT 65.06 263.4 65.26 263.52 ;
      RECT 63.62 263.4 63.82 263.52 ;
      RECT 65.42 262.14 65.62 262.26 ;
      RECT 64.7 262.14 64.9 262.26 ;
      RECT 63.98 262.14 64.18 262.26 ;
      RECT 63.26 262.14 63.46 262.26 ;
      RECT 63.98 267.18 64.18 267.3 ;
      RECT 65.42 266.94 65.62 267.06 ;
      RECT 64.7 266.94 64.9 267.06 ;
      RECT 63.26 266.94 63.46 267.06 ;
      RECT 65.06 265.92 65.26 266.04 ;
      RECT 63.62 265.68 63.82 265.8 ;
      RECT 65.42 269.7 65.62 269.82 ;
      RECT 63.98 269.7 64.18 269.82 ;
      RECT 64.7 269.46 64.9 269.58 ;
      RECT 63.26 269.46 63.46 269.58 ;
      RECT 65.06 268.44 65.26 268.56 ;
      RECT 63.62 268.2 63.82 268.32 ;
      RECT 65.06 270.96 65.26 271.08 ;
      RECT 63.62 270.72 63.82 270.84 ;
      RECT 64.7 272.22 64.9 272.34 ;
      RECT 63.26 272.22 63.46 272.34 ;
      RECT 65.42 271.98 65.62 272.1 ;
      RECT 63.98 271.98 64.18 272.1 ;
      RECT 63.62 275.76 63.82 275.88 ;
      RECT 65.42 274.74 65.62 274.86 ;
      RECT 63.26 274.74 63.46 274.86 ;
      RECT 64.7 274.5 64.9 274.62 ;
      RECT 63.98 274.5 64.18 274.62 ;
      RECT 65.06 273.24 65.26 273.36 ;
      RECT 63.62 273.24 63.82 273.36 ;
      RECT 63.62 278.28 63.82 278.4 ;
      RECT 65.42 277.26 65.62 277.38 ;
      RECT 64.7 277.26 64.9 277.38 ;
      RECT 63.26 277.26 63.46 277.38 ;
      RECT 63.98 277.02 64.18 277.14 ;
      RECT 65.06 276 65.26 276.12 ;
      RECT 65.06 278.52 65.26 278.64 ;
      RECT 59.66 283.087 59.86 283.207 ;
      RECT 58.94 283.087 59.14 283.207 ;
      RECT 58.22 283.087 58.42 283.207 ;
      RECT 60.74 210.958 60.94 211.078 ;
      RECT 65.06 210.958 65.26 211.078 ;
      RECT 58.58 210.48 58.78 210.6 ;
      RECT 60.02 210.48 60.22 210.6 ;
      RECT 64.34 210.48 64.54 210.6 ;
      RECT 58.58 215.52 58.78 215.64 ;
      RECT 64.34 215.52 64.54 215.64 ;
      RECT 60.02 215.28 60.22 215.4 ;
      RECT 65.42 214.26 65.62 214.38 ;
      RECT 63.98 214.26 64.18 214.38 ;
      RECT 63.26 214.26 63.46 214.38 ;
      RECT 58.94 214.26 59.14 214.38 ;
      RECT 58.22 214.26 58.42 214.38 ;
      RECT 64.7 214.02 64.9 214.14 ;
      RECT 61.1 214.02 61.3 214.14 ;
      RECT 60.38 214.02 60.58 214.14 ;
      RECT 59.66 214.02 59.86 214.14 ;
      RECT 59.3 213.718 59.5 213.838 ;
      RECT 63.62 213.718 63.82 213.838 ;
      RECT 65.06 213.718 65.26 213.838 ;
      RECT 57.86 213.478 58.06 213.598 ;
      RECT 60.74 213.478 60.94 213.598 ;
      RECT 58.58 213 58.78 213.12 ;
      RECT 64.34 213 64.54 213.12 ;
      RECT 65.42 216.78 65.62 216.9 ;
      RECT 64.7 216.78 64.9 216.9 ;
      RECT 63.26 216.78 63.46 216.9 ;
      RECT 60.38 216.78 60.58 216.9 ;
      RECT 59.66 216.78 59.86 216.9 ;
      RECT 63.98 216.54 64.18 216.66 ;
      RECT 61.1 216.54 61.3 216.66 ;
      RECT 58.94 216.54 59.14 216.66 ;
      RECT 58.22 216.54 58.42 216.66 ;
      RECT 63.62 216.238 63.82 216.358 ;
      RECT 59.3 216.238 59.5 216.358 ;
      RECT 57.86 215.998 58.06 216.118 ;
      RECT 60.74 215.998 60.94 216.118 ;
      RECT 65.06 215.998 65.26 216.118 ;
      RECT 57.86 221.038 58.06 221.158 ;
      RECT 63.62 221.038 63.82 221.158 ;
      RECT 65.06 221.038 65.26 221.158 ;
      RECT 65.42 219.3 65.62 219.42 ;
      RECT 64.7 219.3 64.9 219.42 ;
      RECT 63.26 219.3 63.46 219.42 ;
      RECT 60.38 219.3 60.58 219.42 ;
      RECT 58.22 219.3 58.42 219.42 ;
      RECT 58.94 219.06 59.14 219.18 ;
      RECT 59.66 219.06 59.86 219.18 ;
      RECT 61.1 219.06 61.3 219.18 ;
      RECT 63.98 219.06 64.18 219.18 ;
      RECT 57.86 218.758 58.06 218.878 ;
      RECT 60.74 218.758 60.94 218.878 ;
      RECT 65.06 218.758 65.26 218.878 ;
      RECT 59.3 218.518 59.5 218.638 ;
      RECT 63.62 218.518 63.82 218.638 ;
      RECT 58.22 223.798 58.42 223.918 ;
      RECT 58.94 223.798 59.14 223.918 ;
      RECT 61.1 223.798 61.3 223.918 ;
      RECT 63.98 223.798 64.18 223.918 ;
      RECT 65.42 223.798 65.62 223.918 ;
      RECT 59.66 223.558 59.86 223.678 ;
      RECT 60.38 223.558 60.58 223.678 ;
      RECT 63.26 223.558 63.46 223.678 ;
      RECT 64.7 223.558 64.9 223.678 ;
      RECT 60.02 223.08 60.22 223.2 ;
      RECT 58.58 222.84 58.78 222.96 ;
      RECT 64.34 222.84 64.54 222.96 ;
      RECT 65.06 222.362 65.26 222.482 ;
      RECT 63.62 222.122 63.82 222.242 ;
      RECT 59.3 221.278 59.5 221.398 ;
      RECT 60.74 221.278 60.94 221.398 ;
      RECT 63.26 229.14 63.46 229.26 ;
      RECT 64.7 229.14 64.9 229.26 ;
      RECT 65.42 229.14 65.62 229.26 ;
      RECT 57.5 228.36 57.7 228.48 ;
      RECT 58.22 228.36 58.42 228.48 ;
      RECT 58.94 228.36 59.14 228.48 ;
      RECT 59.66 228.36 59.86 228.48 ;
      RECT 60.38 228.36 60.58 228.48 ;
      RECT 63.62 228.12 63.82 228.24 ;
      RECT 65.06 227.88 65.26 228 ;
      RECT 60.74 227.73 60.94 227.85 ;
      RECT 59.3 227.73 59.5 227.85 ;
      RECT 57.86 227.73 58.06 227.85 ;
      RECT 65.42 231.9 65.62 232.02 ;
      RECT 63.98 231.9 64.18 232.02 ;
      RECT 64.7 231.66 64.9 231.78 ;
      RECT 63.26 231.66 63.46 231.78 ;
      RECT 63.62 230.64 63.82 230.76 ;
      RECT 65.06 230.4 65.26 230.52 ;
      RECT 63.98 229.38 64.18 229.5 ;
      RECT 63.26 234.42 63.46 234.54 ;
      RECT 64.7 234.42 64.9 234.54 ;
      RECT 63.98 234.18 64.18 234.3 ;
      RECT 65.42 234.18 65.62 234.3 ;
      RECT 63.62 233.16 63.82 233.28 ;
      RECT 65.06 232.92 65.26 233.04 ;
      RECT 63.26 236.94 63.46 237.06 ;
      RECT 64.7 236.94 64.9 237.06 ;
      RECT 65.42 236.7 65.62 236.82 ;
      RECT 63.98 236.7 64.18 236.82 ;
      RECT 63.62 235.68 63.82 235.8 ;
      RECT 63.98 198.9 64.18 199.02 ;
      RECT 63.26 198.9 63.46 199.02 ;
      RECT 61.1 198.9 61.3 199.02 ;
      RECT 60.38 198.9 60.58 199.02 ;
      RECT 58.94 198.9 59.14 199.02 ;
      RECT 60.74 198.422 60.94 198.542 ;
      RECT 63.62 198.422 63.82 198.542 ;
      RECT 65.06 198.422 65.26 198.542 ;
      RECT 57.86 198.182 58.06 198.302 ;
      RECT 59.3 198.182 59.5 198.302 ;
      RECT 60.02 197.88 60.22 198 ;
      RECT 64.34 197.88 64.54 198 ;
      RECT 58.58 197.64 58.78 197.76 ;
      RECT 65.42 196.62 65.62 196.74 ;
      RECT 63.98 196.62 64.18 196.74 ;
      RECT 59.66 196.62 59.86 196.74 ;
      RECT 58.22 196.62 58.42 196.74 ;
      RECT 57.5 196.62 57.7 196.74 ;
      RECT 63.98 201.66 64.18 201.78 ;
      RECT 61.1 201.66 61.3 201.78 ;
      RECT 59.66 201.66 59.86 201.78 ;
      RECT 57.5 201.42 57.7 201.54 ;
      RECT 58.22 201.42 58.42 201.54 ;
      RECT 58.94 201.42 59.14 201.54 ;
      RECT 60.38 201.42 60.58 201.54 ;
      RECT 63.26 201.42 63.46 201.54 ;
      RECT 64.7 201.42 64.9 201.54 ;
      RECT 65.42 201.42 65.62 201.54 ;
      RECT 57.86 200.942 58.06 201.062 ;
      RECT 59.3 200.942 59.5 201.062 ;
      RECT 65.06 200.702 65.26 200.822 ;
      RECT 63.62 200.702 63.82 200.822 ;
      RECT 60.74 200.702 60.94 200.822 ;
      RECT 64.34 200.4 64.54 200.52 ;
      RECT 58.58 200.4 58.78 200.52 ;
      RECT 60.02 200.16 60.22 200.28 ;
      RECT 57.5 204.18 57.7 204.3 ;
      RECT 58.94 204.18 59.14 204.3 ;
      RECT 61.1 204.18 61.3 204.3 ;
      RECT 65.42 203.94 65.62 204.06 ;
      RECT 64.7 203.94 64.9 204.06 ;
      RECT 63.98 203.94 64.18 204.06 ;
      RECT 63.26 203.94 63.46 204.06 ;
      RECT 60.38 203.94 60.58 204.06 ;
      RECT 59.66 203.94 59.86 204.06 ;
      RECT 58.22 203.94 58.42 204.06 ;
      RECT 65.06 203.462 65.26 203.582 ;
      RECT 59.3 203.462 59.5 203.582 ;
      RECT 63.62 203.222 63.82 203.342 ;
      RECT 60.74 203.222 60.94 203.342 ;
      RECT 57.86 203.222 58.06 203.342 ;
      RECT 60.02 202.92 60.22 203.04 ;
      RECT 58.58 202.92 58.78 203.04 ;
      RECT 64.34 202.68 64.54 202.8 ;
      RECT 64.7 206.7 64.9 206.82 ;
      RECT 61.1 206.7 61.3 206.82 ;
      RECT 60.38 206.7 60.58 206.82 ;
      RECT 58.94 206.7 59.14 206.82 ;
      RECT 58.22 206.7 58.42 206.82 ;
      RECT 65.42 206.46 65.62 206.58 ;
      RECT 63.98 206.46 64.18 206.58 ;
      RECT 63.26 206.46 63.46 206.58 ;
      RECT 59.66 206.46 59.86 206.58 ;
      RECT 57.5 206.46 57.7 206.58 ;
      RECT 63.62 205.982 63.82 206.102 ;
      RECT 59.3 205.982 59.5 206.102 ;
      RECT 57.86 205.982 58.06 206.102 ;
      RECT 60.74 205.742 60.94 205.862 ;
      RECT 65.06 205.742 65.26 205.862 ;
      RECT 64.34 205.44 64.54 205.56 ;
      RECT 60.02 205.2 60.22 205.32 ;
      RECT 58.58 205.2 58.78 205.32 ;
      RECT 63.26 209.22 63.46 209.34 ;
      RECT 61.1 209.22 61.3 209.34 ;
      RECT 60.38 209.22 60.58 209.34 ;
      RECT 58.94 209.22 59.14 209.34 ;
      RECT 58.22 209.22 58.42 209.34 ;
      RECT 59.66 208.98 59.86 209.1 ;
      RECT 63.98 208.98 64.18 209.1 ;
      RECT 64.7 208.98 64.9 209.1 ;
      RECT 65.42 208.98 65.62 209.1 ;
      RECT 59.3 208.502 59.5 208.622 ;
      RECT 63.62 208.502 63.82 208.622 ;
      RECT 57.86 208.262 58.06 208.382 ;
      RECT 60.74 208.262 60.94 208.382 ;
      RECT 65.06 208.262 65.26 208.382 ;
      RECT 58.58 207.96 58.78 208.08 ;
      RECT 60.02 207.96 60.22 208.08 ;
      RECT 64.34 207.72 64.54 207.84 ;
      RECT 60.02 212.76 60.22 212.88 ;
      RECT 64.7 211.74 64.9 211.86 ;
      RECT 63.26 211.74 63.46 211.86 ;
      RECT 59.66 211.74 59.86 211.86 ;
      RECT 58.94 211.74 59.14 211.86 ;
      RECT 58.22 211.74 58.42 211.86 ;
      RECT 60.38 211.5 60.58 211.62 ;
      RECT 61.1 211.5 61.3 211.62 ;
      RECT 65.42 211.5 65.62 211.62 ;
      RECT 63.98 211.5 64.18 211.62 ;
      RECT 59.3 211.198 59.5 211.318 ;
      RECT 63.62 211.198 63.82 211.318 ;
      RECT 57.86 210.958 58.06 211.078 ;
      RECT 58.22 181.26 58.42 181.38 ;
      RECT 64.34 180.24 64.54 180.36 ;
      RECT 60.02 185.28 60.22 185.4 ;
      RECT 64.34 185.04 64.54 185.16 ;
      RECT 58.58 185.04 58.78 185.16 ;
      RECT 64.7 184.02 64.9 184.14 ;
      RECT 59.66 184.02 59.86 184.14 ;
      RECT 58.94 184.02 59.14 184.14 ;
      RECT 57.5 184.02 57.7 184.14 ;
      RECT 65.42 183.78 65.62 183.9 ;
      RECT 63.98 183.78 64.18 183.9 ;
      RECT 63.26 183.78 63.46 183.9 ;
      RECT 61.1 183.78 61.3 183.9 ;
      RECT 60.38 183.78 60.58 183.9 ;
      RECT 58.22 183.78 58.42 183.9 ;
      RECT 60.02 187.8 60.22 187.92 ;
      RECT 64.34 187.56 64.54 187.68 ;
      RECT 58.58 187.56 58.78 187.68 ;
      RECT 58.94 186.54 59.14 186.66 ;
      RECT 63.26 186.54 63.46 186.66 ;
      RECT 63.98 186.54 64.18 186.66 ;
      RECT 65.42 186.54 65.62 186.66 ;
      RECT 57.5 186.3 57.7 186.42 ;
      RECT 58.22 186.3 58.42 186.42 ;
      RECT 59.66 186.3 59.86 186.42 ;
      RECT 60.38 186.3 60.58 186.42 ;
      RECT 61.1 186.3 61.3 186.42 ;
      RECT 64.7 186.3 64.9 186.42 ;
      RECT 57.86 190.862 58.06 190.982 ;
      RECT 59.3 190.862 59.5 190.982 ;
      RECT 60.74 190.862 60.94 190.982 ;
      RECT 63.62 190.622 63.82 190.742 ;
      RECT 65.06 190.622 65.26 190.742 ;
      RECT 64.34 190.32 64.54 190.44 ;
      RECT 58.58 190.32 58.78 190.44 ;
      RECT 60.02 190.08 60.22 190.2 ;
      RECT 58.94 189.06 59.14 189.18 ;
      RECT 61.1 189.06 61.3 189.18 ;
      RECT 63.26 189.06 63.46 189.18 ;
      RECT 63.98 189.06 64.18 189.18 ;
      RECT 65.42 189.06 65.62 189.18 ;
      RECT 64.7 188.82 64.9 188.94 ;
      RECT 60.38 188.82 60.58 188.94 ;
      RECT 59.66 188.82 59.86 188.94 ;
      RECT 58.22 188.82 58.42 188.94 ;
      RECT 57.5 188.82 57.7 188.94 ;
      RECT 59.66 193.86 59.86 193.98 ;
      RECT 60.38 193.86 60.58 193.98 ;
      RECT 63.26 193.86 63.46 193.98 ;
      RECT 64.7 193.86 64.9 193.98 ;
      RECT 65.42 193.86 65.62 193.98 ;
      RECT 57.86 193.382 58.06 193.502 ;
      RECT 60.74 193.382 60.94 193.502 ;
      RECT 63.62 193.382 63.82 193.502 ;
      RECT 59.3 193.142 59.5 193.262 ;
      RECT 65.06 193.142 65.26 193.262 ;
      RECT 58.58 192.84 58.78 192.96 ;
      RECT 60.02 192.6 60.22 192.72 ;
      RECT 64.34 192.6 64.54 192.72 ;
      RECT 59.3 192.122 59.5 192.242 ;
      RECT 60.74 192.122 60.94 192.242 ;
      RECT 63.62 192.122 63.82 192.242 ;
      RECT 57.86 191.882 58.06 192.002 ;
      RECT 65.06 191.882 65.26 192.002 ;
      RECT 64.7 191.58 64.9 191.7 ;
      RECT 63.98 191.58 64.18 191.7 ;
      RECT 61.1 191.58 61.3 191.7 ;
      RECT 59.66 191.58 59.86 191.7 ;
      RECT 58.94 191.58 59.14 191.7 ;
      RECT 57.5 191.58 57.7 191.7 ;
      RECT 58.22 191.34 58.42 191.46 ;
      RECT 60.38 191.34 60.58 191.46 ;
      RECT 63.26 191.34 63.46 191.46 ;
      RECT 65.42 191.34 65.62 191.46 ;
      RECT 57.86 194.642 58.06 194.762 ;
      RECT 60.74 194.642 60.94 194.762 ;
      RECT 63.62 194.642 63.82 194.762 ;
      RECT 65.06 194.402 65.26 194.522 ;
      RECT 59.3 194.402 59.5 194.522 ;
      RECT 63.98 194.1 64.18 194.22 ;
      RECT 61.1 194.1 61.3 194.22 ;
      RECT 58.94 194.1 59.14 194.22 ;
      RECT 58.22 194.1 58.42 194.22 ;
      RECT 57.5 194.1 57.7 194.22 ;
      RECT 58.94 196.38 59.14 196.5 ;
      RECT 60.38 196.38 60.58 196.5 ;
      RECT 61.1 196.38 61.3 196.5 ;
      RECT 63.26 196.38 63.46 196.5 ;
      RECT 64.7 196.38 64.9 196.5 ;
      RECT 59.3 195.902 59.5 196.022 ;
      RECT 63.62 195.902 63.82 196.022 ;
      RECT 65.06 195.662 65.26 195.782 ;
      RECT 60.74 195.662 60.94 195.782 ;
      RECT 57.86 195.662 58.06 195.782 ;
      RECT 64.34 195.36 64.54 195.48 ;
      RECT 58.58 195.12 58.78 195.24 ;
      RECT 60.02 195.12 60.22 195.24 ;
      RECT 57.5 199.14 57.7 199.26 ;
      RECT 58.22 199.14 58.42 199.26 ;
      RECT 59.66 199.14 59.86 199.26 ;
      RECT 65.42 199.14 65.62 199.26 ;
      RECT 64.7 198.9 64.9 199.02 ;
      RECT 61.1 161.1 61.3 161.22 ;
      RECT 63.26 161.1 63.46 161.22 ;
      RECT 63.98 161.1 64.18 161.22 ;
      RECT 64.7 161.1 64.9 161.22 ;
      RECT 65.42 161.1 65.62 161.22 ;
      RECT 64.7 166.38 64.9 166.5 ;
      RECT 63.98 166.38 64.18 166.5 ;
      RECT 59.66 166.38 59.86 166.5 ;
      RECT 58.94 166.38 59.14 166.5 ;
      RECT 65.42 166.14 65.62 166.26 ;
      RECT 63.26 166.14 63.46 166.26 ;
      RECT 61.1 166.14 61.3 166.26 ;
      RECT 60.38 166.14 60.58 166.26 ;
      RECT 58.22 166.14 58.42 166.26 ;
      RECT 57.5 166.14 57.7 166.26 ;
      RECT 60.02 165.12 60.22 165.24 ;
      RECT 58.58 165.12 58.78 165.24 ;
      RECT 64.34 164.88 64.54 165 ;
      RECT 65.42 163.86 65.62 163.98 ;
      RECT 63.98 163.86 64.18 163.98 ;
      RECT 61.1 163.86 61.3 163.98 ;
      RECT 58.94 163.86 59.14 163.98 ;
      RECT 57.5 163.86 57.7 163.98 ;
      RECT 65.42 168.9 65.62 169.02 ;
      RECT 63.98 168.9 64.18 169.02 ;
      RECT 61.1 168.9 61.3 169.02 ;
      RECT 60.38 168.9 60.58 169.02 ;
      RECT 58.22 168.9 58.42 169.02 ;
      RECT 57.5 168.66 57.7 168.78 ;
      RECT 58.94 168.66 59.14 168.78 ;
      RECT 59.66 168.66 59.86 168.78 ;
      RECT 63.26 168.66 63.46 168.78 ;
      RECT 64.7 168.66 64.9 168.78 ;
      RECT 64.34 167.64 64.54 167.76 ;
      RECT 58.58 167.4 58.78 167.52 ;
      RECT 60.02 167.4 60.22 167.52 ;
      RECT 63.98 171.42 64.18 171.54 ;
      RECT 63.26 171.42 63.46 171.54 ;
      RECT 59.66 171.42 59.86 171.54 ;
      RECT 58.22 171.42 58.42 171.54 ;
      RECT 57.5 171.42 57.7 171.54 ;
      RECT 58.94 171.18 59.14 171.3 ;
      RECT 65.42 171.18 65.62 171.3 ;
      RECT 64.7 171.18 64.9 171.3 ;
      RECT 61.1 171.18 61.3 171.3 ;
      RECT 60.38 171.18 60.58 171.3 ;
      RECT 64.34 170.16 64.54 170.28 ;
      RECT 60.02 170.16 60.22 170.28 ;
      RECT 58.58 170.16 58.78 170.28 ;
      RECT 65.42 173.94 65.62 174.06 ;
      RECT 63.98 173.94 64.18 174.06 ;
      RECT 59.66 173.94 59.86 174.06 ;
      RECT 58.94 173.94 59.14 174.06 ;
      RECT 58.22 173.94 58.42 174.06 ;
      RECT 57.5 173.7 57.7 173.82 ;
      RECT 60.38 173.7 60.58 173.82 ;
      RECT 61.1 173.7 61.3 173.82 ;
      RECT 63.26 173.7 63.46 173.82 ;
      RECT 64.7 173.7 64.9 173.82 ;
      RECT 64.34 172.68 64.54 172.8 ;
      RECT 60.02 172.68 60.22 172.8 ;
      RECT 58.58 172.44 58.78 172.56 ;
      RECT 64.34 177.48 64.54 177.6 ;
      RECT 58.58 177.48 58.78 177.6 ;
      RECT 64.7 176.46 64.9 176.58 ;
      RECT 63.98 176.46 64.18 176.58 ;
      RECT 63.26 176.46 63.46 176.58 ;
      RECT 60.38 176.46 60.58 176.58 ;
      RECT 59.66 176.46 59.86 176.58 ;
      RECT 58.94 176.46 59.14 176.58 ;
      RECT 58.22 176.46 58.42 176.58 ;
      RECT 65.42 176.22 65.62 176.34 ;
      RECT 61.1 176.22 61.3 176.34 ;
      RECT 57.5 176.22 57.7 176.34 ;
      RECT 58.58 174.96 58.78 175.08 ;
      RECT 60.02 174.96 60.22 175.08 ;
      RECT 64.34 174.96 64.54 175.08 ;
      RECT 60.02 180 60.22 180.12 ;
      RECT 58.58 180 58.78 180.12 ;
      RECT 65.42 178.98 65.62 179.1 ;
      RECT 64.7 178.98 64.9 179.1 ;
      RECT 58.94 178.98 59.14 179.1 ;
      RECT 58.22 178.98 58.42 179.1 ;
      RECT 57.5 178.98 57.7 179.1 ;
      RECT 63.98 178.74 64.18 178.86 ;
      RECT 63.26 178.74 63.46 178.86 ;
      RECT 61.1 178.74 61.3 178.86 ;
      RECT 60.38 178.74 60.58 178.86 ;
      RECT 59.66 178.74 59.86 178.86 ;
      RECT 60.02 177.72 60.22 177.84 ;
      RECT 60.02 182.76 60.22 182.88 ;
      RECT 58.58 182.76 58.78 182.88 ;
      RECT 64.34 182.52 64.54 182.64 ;
      RECT 57.5 181.5 57.7 181.62 ;
      RECT 58.94 181.5 59.14 181.62 ;
      RECT 59.66 181.5 59.86 181.62 ;
      RECT 60.38 181.5 60.58 181.62 ;
      RECT 64.7 181.5 64.9 181.62 ;
      RECT 65.42 181.26 65.62 181.38 ;
      RECT 63.98 181.26 64.18 181.38 ;
      RECT 63.26 181.26 63.46 181.38 ;
      RECT 61.1 181.26 61.3 181.38 ;
      RECT 58.58 142.2 58.78 142.32 ;
      RECT 57.5 145.98 57.7 146.1 ;
      RECT 58.22 145.98 58.42 146.1 ;
      RECT 58.94 145.98 59.14 146.1 ;
      RECT 59.66 145.98 59.86 146.1 ;
      RECT 60.38 145.98 60.58 146.1 ;
      RECT 61.1 145.98 61.3 146.1 ;
      RECT 63.26 145.98 63.46 146.1 ;
      RECT 63.98 145.98 64.18 146.1 ;
      RECT 64.7 145.98 64.9 146.1 ;
      RECT 65.42 145.98 65.62 146.1 ;
      RECT 58.58 144.96 58.78 145.08 ;
      RECT 64.34 144.96 64.54 145.08 ;
      RECT 60.02 144.72 60.22 144.84 ;
      RECT 64.34 150 64.54 150.12 ;
      RECT 58.58 150 58.78 150.12 ;
      RECT 60.02 149.76 60.22 149.88 ;
      RECT 59.66 148.74 59.86 148.86 ;
      RECT 63.98 148.74 64.18 148.86 ;
      RECT 61.1 148.5 61.3 148.62 ;
      RECT 63.26 148.5 63.46 148.62 ;
      RECT 64.7 148.5 64.9 148.62 ;
      RECT 65.42 148.5 65.62 148.62 ;
      RECT 60.38 148.5 60.58 148.62 ;
      RECT 58.94 148.5 59.14 148.62 ;
      RECT 58.22 148.5 58.42 148.62 ;
      RECT 57.5 148.5 57.7 148.62 ;
      RECT 64.34 152.52 64.54 152.64 ;
      RECT 60.02 152.52 60.22 152.64 ;
      RECT 58.58 152.28 58.78 152.4 ;
      RECT 61.1 151.26 61.3 151.38 ;
      RECT 63.98 151.26 64.18 151.38 ;
      RECT 65.42 151.26 65.62 151.38 ;
      RECT 64.7 151.02 64.9 151.14 ;
      RECT 63.26 151.02 63.46 151.14 ;
      RECT 60.38 151.02 60.58 151.14 ;
      RECT 59.66 151.02 59.86 151.14 ;
      RECT 58.94 151.02 59.14 151.14 ;
      RECT 58.22 151.02 58.42 151.14 ;
      RECT 57.5 151.02 57.7 151.14 ;
      RECT 64.34 155.04 64.54 155.16 ;
      RECT 60.02 154.8 60.22 154.92 ;
      RECT 58.58 154.8 58.78 154.92 ;
      RECT 65.42 153.78 65.62 153.9 ;
      RECT 63.98 153.78 64.18 153.9 ;
      RECT 61.1 153.78 61.3 153.9 ;
      RECT 64.7 153.54 64.9 153.66 ;
      RECT 63.26 153.54 63.46 153.66 ;
      RECT 60.38 153.54 60.58 153.66 ;
      RECT 59.66 153.54 59.86 153.66 ;
      RECT 58.94 153.54 59.14 153.66 ;
      RECT 58.22 153.54 58.42 153.66 ;
      RECT 57.5 153.54 57.7 153.66 ;
      RECT 63.62 158.278 63.82 158.398 ;
      RECT 59.3 158.278 59.5 158.398 ;
      RECT 65.06 158.038 65.26 158.158 ;
      RECT 60.74 158.038 60.94 158.158 ;
      RECT 57.86 158.038 58.06 158.158 ;
      RECT 60.02 157.56 60.22 157.68 ;
      RECT 58.58 157.56 58.78 157.68 ;
      RECT 64.34 157.32 64.54 157.44 ;
      RECT 63.62 156.842 63.82 156.962 ;
      RECT 59.3 156.842 59.5 156.962 ;
      RECT 65.06 156.602 65.26 156.722 ;
      RECT 60.74 156.602 60.94 156.722 ;
      RECT 57.86 156.602 58.06 156.722 ;
      RECT 58.22 156.3 58.42 156.42 ;
      RECT 58.94 156.3 59.14 156.42 ;
      RECT 63.26 156.3 63.46 156.42 ;
      RECT 65.42 156.3 65.62 156.42 ;
      RECT 64.7 156.06 64.9 156.18 ;
      RECT 63.98 156.06 64.18 156.18 ;
      RECT 61.1 156.06 61.3 156.18 ;
      RECT 60.38 156.06 60.58 156.18 ;
      RECT 59.66 156.06 59.86 156.18 ;
      RECT 57.5 156.06 57.7 156.18 ;
      RECT 60.02 160.08 60.22 160.2 ;
      RECT 64.34 159.84 64.54 159.96 ;
      RECT 58.58 159.84 58.78 159.96 ;
      RECT 58.22 158.82 58.42 158.94 ;
      RECT 60.38 158.82 60.58 158.94 ;
      RECT 64.7 158.82 64.9 158.94 ;
      RECT 57.5 158.58 57.7 158.7 ;
      RECT 58.94 158.58 59.14 158.7 ;
      RECT 59.66 158.58 59.86 158.7 ;
      RECT 61.1 158.58 61.3 158.7 ;
      RECT 63.26 158.58 63.46 158.7 ;
      RECT 63.98 158.58 64.18 158.7 ;
      RECT 65.42 158.58 65.62 158.7 ;
      RECT 58.22 163.62 58.42 163.74 ;
      RECT 59.66 163.62 59.86 163.74 ;
      RECT 60.38 163.62 60.58 163.74 ;
      RECT 63.26 163.62 63.46 163.74 ;
      RECT 64.7 163.62 64.9 163.74 ;
      RECT 64.34 162.36 64.54 162.48 ;
      RECT 60.02 162.36 60.22 162.48 ;
      RECT 58.58 162.36 58.78 162.48 ;
      RECT 57.5 161.1 57.7 161.22 ;
      RECT 58.22 161.1 58.42 161.22 ;
      RECT 58.94 161.1 59.14 161.22 ;
      RECT 59.66 161.1 59.86 161.22 ;
      RECT 60.38 161.1 60.58 161.22 ;
      RECT 60.38 133.38 60.58 133.5 ;
      RECT 59.66 133.38 59.86 133.5 ;
      RECT 58.94 133.38 59.14 133.5 ;
      RECT 58.22 133.38 58.42 133.5 ;
      RECT 58.58 132.36 58.78 132.48 ;
      RECT 64.34 132.12 64.54 132.24 ;
      RECT 60.02 132.12 60.22 132.24 ;
      RECT 57.5 131.578 57.7 131.698 ;
      RECT 58.22 131.578 58.42 131.698 ;
      RECT 58.94 131.578 59.14 131.698 ;
      RECT 59.66 131.578 59.86 131.698 ;
      RECT 60.38 131.578 60.58 131.698 ;
      RECT 61.1 131.578 61.3 131.698 ;
      RECT 63.26 131.578 63.46 131.698 ;
      RECT 63.98 131.578 64.18 131.698 ;
      RECT 64.7 131.578 64.9 131.698 ;
      RECT 65.42 131.578 65.62 131.698 ;
      RECT 64.7 131.1 64.9 131.22 ;
      RECT 63.26 131.1 63.46 131.22 ;
      RECT 59.66 131.1 59.86 131.22 ;
      RECT 58.22 131.1 58.42 131.22 ;
      RECT 58.22 136.14 58.42 136.26 ;
      RECT 59.66 136.14 59.86 136.26 ;
      RECT 63.26 136.14 63.46 136.26 ;
      RECT 63.98 136.14 64.18 136.26 ;
      RECT 64.7 136.14 64.9 136.26 ;
      RECT 65.42 136.14 65.62 136.26 ;
      RECT 61.1 135.9 61.3 136.02 ;
      RECT 60.38 135.9 60.58 136.02 ;
      RECT 58.94 135.9 59.14 136.02 ;
      RECT 57.5 135.9 57.7 136.02 ;
      RECT 64.34 134.88 64.54 135 ;
      RECT 58.58 134.88 58.78 135 ;
      RECT 60.02 134.64 60.22 134.76 ;
      RECT 57.5 134.098 57.7 134.218 ;
      RECT 58.22 134.098 58.42 134.218 ;
      RECT 58.94 134.098 59.14 134.218 ;
      RECT 59.66 134.098 59.86 134.218 ;
      RECT 60.38 134.098 60.58 134.218 ;
      RECT 61.1 134.098 61.3 134.218 ;
      RECT 63.26 134.098 63.46 134.218 ;
      RECT 63.98 134.098 64.18 134.218 ;
      RECT 64.7 134.098 64.9 134.218 ;
      RECT 65.42 134.098 65.62 134.218 ;
      RECT 57.5 139.138 57.7 139.258 ;
      RECT 58.22 139.138 58.42 139.258 ;
      RECT 58.94 139.138 59.14 139.258 ;
      RECT 59.66 139.138 59.86 139.258 ;
      RECT 60.38 139.138 60.58 139.258 ;
      RECT 61.1 139.138 61.3 139.258 ;
      RECT 63.26 139.138 63.46 139.258 ;
      RECT 63.98 139.138 64.18 139.258 ;
      RECT 64.7 139.138 64.9 139.258 ;
      RECT 65.42 139.138 65.62 139.258 ;
      RECT 64.7 138.66 64.9 138.78 ;
      RECT 63.98 138.66 64.18 138.78 ;
      RECT 61.1 138.66 61.3 138.78 ;
      RECT 58.22 138.66 58.42 138.78 ;
      RECT 65.42 138.42 65.62 138.54 ;
      RECT 63.26 138.42 63.46 138.54 ;
      RECT 60.38 138.42 60.58 138.54 ;
      RECT 59.66 138.42 59.86 138.54 ;
      RECT 58.94 138.42 59.14 138.54 ;
      RECT 57.5 138.42 57.7 138.54 ;
      RECT 58.58 137.4 58.78 137.52 ;
      RECT 64.34 137.4 64.54 137.52 ;
      RECT 60.02 137.16 60.22 137.28 ;
      RECT 57.5 136.618 57.7 136.738 ;
      RECT 58.22 136.618 58.42 136.738 ;
      RECT 58.94 136.618 59.14 136.738 ;
      RECT 59.66 136.618 59.86 136.738 ;
      RECT 60.38 136.618 60.58 136.738 ;
      RECT 61.1 136.618 61.3 136.738 ;
      RECT 63.26 136.618 63.46 136.738 ;
      RECT 63.98 136.618 64.18 136.738 ;
      RECT 64.7 136.618 64.9 136.738 ;
      RECT 65.42 136.618 65.62 136.738 ;
      RECT 65.42 141.18 65.62 141.3 ;
      RECT 64.7 141.18 64.9 141.3 ;
      RECT 63.26 141.18 63.46 141.3 ;
      RECT 58.94 141.18 59.14 141.3 ;
      RECT 57.5 140.94 57.7 141.06 ;
      RECT 58.22 140.94 58.42 141.06 ;
      RECT 59.66 140.94 59.86 141.06 ;
      RECT 60.38 140.94 60.58 141.06 ;
      RECT 61.1 140.94 61.3 141.06 ;
      RECT 63.98 140.94 64.18 141.06 ;
      RECT 64.34 139.92 64.54 140.04 ;
      RECT 60.02 139.92 60.22 140.04 ;
      RECT 58.58 139.68 58.78 139.8 ;
      RECT 64.7 143.7 64.9 143.82 ;
      RECT 63.98 143.7 64.18 143.82 ;
      RECT 63.26 143.7 63.46 143.82 ;
      RECT 60.38 143.7 60.58 143.82 ;
      RECT 59.66 143.7 59.86 143.82 ;
      RECT 58.22 143.7 58.42 143.82 ;
      RECT 65.42 143.46 65.62 143.58 ;
      RECT 61.1 143.46 61.3 143.58 ;
      RECT 58.94 143.46 59.14 143.58 ;
      RECT 57.5 143.46 57.7 143.58 ;
      RECT 64.34 142.44 64.54 142.56 ;
      RECT 60.02 142.44 60.22 142.56 ;
      RECT 60.02 122.04 60.22 122.16 ;
      RECT 57.5 121.498 57.7 121.618 ;
      RECT 58.22 121.498 58.42 121.618 ;
      RECT 58.94 121.498 59.14 121.618 ;
      RECT 59.66 121.498 59.86 121.618 ;
      RECT 60.38 121.498 60.58 121.618 ;
      RECT 61.1 121.498 61.3 121.618 ;
      RECT 63.26 121.498 63.46 121.618 ;
      RECT 63.98 121.498 64.18 121.618 ;
      RECT 64.7 121.498 64.9 121.618 ;
      RECT 65.42 121.498 65.62 121.618 ;
      RECT 61.1 121.02 61.3 121.14 ;
      RECT 63.26 121.02 63.46 121.14 ;
      RECT 63.98 121.02 64.18 121.14 ;
      RECT 60.38 120.78 60.58 120.9 ;
      RECT 64.7 120.78 64.9 120.9 ;
      RECT 57.5 120.78 57.7 120.9 ;
      RECT 65.42 120.78 65.62 120.9 ;
      RECT 58.22 120.78 58.42 120.9 ;
      RECT 58.94 120.78 59.14 120.9 ;
      RECT 59.66 120.78 59.86 120.9 ;
      RECT 64.34 124.8 64.54 124.92 ;
      RECT 58.58 124.56 58.78 124.68 ;
      RECT 60.02 124.56 60.22 124.68 ;
      RECT 57.5 124.018 57.7 124.138 ;
      RECT 58.22 124.018 58.42 124.138 ;
      RECT 58.94 124.018 59.14 124.138 ;
      RECT 59.66 124.018 59.86 124.138 ;
      RECT 60.38 124.018 60.58 124.138 ;
      RECT 61.1 124.018 61.3 124.138 ;
      RECT 63.26 124.018 63.46 124.138 ;
      RECT 63.98 124.018 64.18 124.138 ;
      RECT 64.7 124.018 64.9 124.138 ;
      RECT 65.42 124.018 65.62 124.138 ;
      RECT 63.26 123.54 63.46 123.66 ;
      RECT 65.42 123.54 65.62 123.66 ;
      RECT 57.5 123.3 57.7 123.42 ;
      RECT 58.22 123.3 58.42 123.42 ;
      RECT 58.94 123.3 59.14 123.42 ;
      RECT 59.66 123.3 59.86 123.42 ;
      RECT 60.38 123.3 60.58 123.42 ;
      RECT 61.1 123.3 61.3 123.42 ;
      RECT 63.98 123.3 64.18 123.42 ;
      RECT 64.7 123.3 64.9 123.42 ;
      RECT 64.34 127.32 64.54 127.44 ;
      RECT 58.58 127.08 58.78 127.2 ;
      RECT 60.02 127.08 60.22 127.2 ;
      RECT 57.5 126.538 57.7 126.658 ;
      RECT 58.22 126.538 58.42 126.658 ;
      RECT 58.94 126.538 59.14 126.658 ;
      RECT 59.66 126.538 59.86 126.658 ;
      RECT 60.38 126.538 60.58 126.658 ;
      RECT 61.1 126.538 61.3 126.658 ;
      RECT 63.26 126.538 63.46 126.658 ;
      RECT 63.98 126.538 64.18 126.658 ;
      RECT 64.7 126.538 64.9 126.658 ;
      RECT 65.42 126.538 65.62 126.658 ;
      RECT 63.26 126.06 63.46 126.18 ;
      RECT 63.98 126.06 64.18 126.18 ;
      RECT 64.7 126.06 64.9 126.18 ;
      RECT 57.5 125.82 57.7 125.94 ;
      RECT 58.22 125.82 58.42 125.94 ;
      RECT 58.94 125.82 59.14 125.94 ;
      RECT 59.66 125.82 59.86 125.94 ;
      RECT 60.38 125.82 60.58 125.94 ;
      RECT 61.1 125.82 61.3 125.94 ;
      RECT 65.42 125.82 65.62 125.94 ;
      RECT 57.5 130.86 57.7 130.98 ;
      RECT 58.94 130.86 59.14 130.98 ;
      RECT 60.38 130.86 60.58 130.98 ;
      RECT 61.1 130.86 61.3 130.98 ;
      RECT 63.98 130.86 64.18 130.98 ;
      RECT 65.42 130.86 65.62 130.98 ;
      RECT 58.58 129.84 58.78 129.96 ;
      RECT 64.34 129.84 64.54 129.96 ;
      RECT 60.02 129.6 60.22 129.72 ;
      RECT 57.5 129.058 57.7 129.178 ;
      RECT 58.22 129.058 58.42 129.178 ;
      RECT 58.94 129.058 59.14 129.178 ;
      RECT 59.66 129.058 59.86 129.178 ;
      RECT 60.38 129.058 60.58 129.178 ;
      RECT 61.1 129.058 61.3 129.178 ;
      RECT 63.26 129.058 63.46 129.178 ;
      RECT 63.98 129.058 64.18 129.178 ;
      RECT 64.7 129.058 64.9 129.178 ;
      RECT 65.42 129.058 65.62 129.178 ;
      RECT 64.7 128.58 64.9 128.7 ;
      RECT 63.26 128.58 63.46 128.7 ;
      RECT 58.22 128.58 58.42 128.7 ;
      RECT 65.42 128.34 65.62 128.46 ;
      RECT 63.98 128.34 64.18 128.46 ;
      RECT 61.1 128.34 61.3 128.46 ;
      RECT 60.38 128.34 60.58 128.46 ;
      RECT 59.66 128.34 59.86 128.46 ;
      RECT 58.94 128.34 59.14 128.46 ;
      RECT 57.5 128.34 57.7 128.46 ;
      RECT 65.42 133.62 65.62 133.74 ;
      RECT 63.98 133.62 64.18 133.74 ;
      RECT 57.5 133.62 57.7 133.74 ;
      RECT 64.7 133.38 64.9 133.5 ;
      RECT 63.26 133.38 63.46 133.5 ;
      RECT 61.1 133.38 61.3 133.5 ;
      RECT 54.62 262.38 54.82 262.5 ;
      RECT 53.9 262.38 54.1 262.5 ;
      RECT 54.98 264.27 55.18 264.39 ;
      RECT 53.54 264.27 53.74 264.39 ;
      RECT 55.34 263.64 55.54 263.76 ;
      RECT 54.62 263.64 54.82 263.76 ;
      RECT 53.9 263.64 54.1 263.76 ;
      RECT 55.34 266.16 55.54 266.28 ;
      RECT 54.62 266.16 54.82 266.28 ;
      RECT 53.9 266.16 54.1 266.28 ;
      RECT 54.98 265.53 55.18 265.65 ;
      RECT 53.54 265.53 53.74 265.65 ;
      RECT 55.34 264.9 55.54 265.02 ;
      RECT 54.62 264.9 54.82 265.02 ;
      RECT 53.9 264.9 54.1 265.02 ;
      RECT 55.34 267.42 55.54 267.54 ;
      RECT 54.62 267.42 54.82 267.54 ;
      RECT 53.9 267.42 54.1 267.54 ;
      RECT 54.98 266.79 55.18 266.91 ;
      RECT 53.54 266.79 53.74 266.91 ;
      RECT 55.34 268.68 55.54 268.8 ;
      RECT 54.62 268.68 54.82 268.8 ;
      RECT 53.9 268.68 54.1 268.8 ;
      RECT 54.98 268.05 55.18 268.17 ;
      RECT 53.54 268.05 53.74 268.17 ;
      RECT 55.34 269.94 55.54 270.06 ;
      RECT 54.62 269.94 54.82 270.06 ;
      RECT 53.9 269.94 54.1 270.06 ;
      RECT 54.98 269.31 55.18 269.43 ;
      RECT 53.54 269.31 53.74 269.43 ;
      RECT 55.34 271.2 55.54 271.32 ;
      RECT 54.62 271.2 54.82 271.32 ;
      RECT 53.9 271.2 54.1 271.32 ;
      RECT 54.98 270.57 55.18 270.69 ;
      RECT 53.54 270.57 53.74 270.69 ;
      RECT 55.34 272.46 55.54 272.58 ;
      RECT 54.62 272.46 54.82 272.58 ;
      RECT 53.9 272.46 54.1 272.58 ;
      RECT 54.98 271.83 55.18 271.95 ;
      RECT 53.54 271.83 53.74 271.95 ;
      RECT 54.98 274.35 55.18 274.47 ;
      RECT 53.54 274.35 53.74 274.47 ;
      RECT 55.34 273.72 55.54 273.84 ;
      RECT 54.62 273.72 54.82 273.84 ;
      RECT 53.9 273.72 54.1 273.84 ;
      RECT 54.98 273.09 55.18 273.21 ;
      RECT 53.54 273.09 53.74 273.21 ;
      RECT 54.98 275.61 55.18 275.73 ;
      RECT 53.54 275.61 53.74 275.73 ;
      RECT 55.34 274.98 55.54 275.1 ;
      RECT 54.62 274.98 54.82 275.1 ;
      RECT 53.9 274.98 54.1 275.1 ;
      RECT 54.98 276.87 55.18 276.99 ;
      RECT 53.54 276.87 53.74 276.99 ;
      RECT 55.34 276.24 55.54 276.36 ;
      RECT 54.62 276.24 54.82 276.36 ;
      RECT 53.9 276.24 54.1 276.36 ;
      RECT 54.98 278.13 55.18 278.25 ;
      RECT 53.54 278.13 53.74 278.25 ;
      RECT 55.34 277.5 55.54 277.62 ;
      RECT 54.62 277.5 54.82 277.62 ;
      RECT 53.9 277.5 54.1 277.62 ;
      RECT 55.34 278.76 55.54 278.88 ;
      RECT 54.62 278.76 54.82 278.88 ;
      RECT 53.9 278.76 54.1 278.88 ;
      RECT 55.34 283.087 55.54 283.207 ;
      RECT 54.62 283.087 54.82 283.207 ;
      RECT 53.9 283.087 54.1 283.207 ;
      RECT 54.26 305.498 54.46 305.618 ;
      RECT 53.9 305.967 54.1 306.087 ;
      RECT 54.62 305.967 54.82 306.087 ;
      RECT 55.34 305.967 55.54 306.087 ;
      RECT 54.26 323.3835 54.46 323.5035 ;
      RECT 55.34 325.9425 55.54 326.0625 ;
      RECT 54.62 325.9425 54.82 326.0625 ;
      RECT 53.9 325.9425 54.1 326.0625 ;
      RECT 54.26 348.339 54.46 348.459 ;
      RECT 64.34 119.76 64.54 119.88 ;
      RECT 60.02 119.52 60.22 119.64 ;
      RECT 58.58 119.52 58.78 119.64 ;
      RECT 57.5 118.978 57.7 119.098 ;
      RECT 58.22 118.978 58.42 119.098 ;
      RECT 58.94 118.978 59.14 119.098 ;
      RECT 59.66 118.978 59.86 119.098 ;
      RECT 60.38 118.978 60.58 119.098 ;
      RECT 61.1 118.978 61.3 119.098 ;
      RECT 63.26 118.978 63.46 119.098 ;
      RECT 63.98 118.978 64.18 119.098 ;
      RECT 64.7 118.978 64.9 119.098 ;
      RECT 65.42 118.978 65.62 119.098 ;
      RECT 65.42 118.5 65.62 118.62 ;
      RECT 64.7 118.5 64.9 118.62 ;
      RECT 60.38 118.5 60.58 118.62 ;
      RECT 59.66 118.5 59.86 118.62 ;
      RECT 58.94 118.5 59.14 118.62 ;
      RECT 58.22 118.5 58.42 118.62 ;
      RECT 63.98 118.26 64.18 118.38 ;
      RECT 63.26 118.26 63.46 118.38 ;
      RECT 61.1 118.26 61.3 118.38 ;
      RECT 57.5 118.26 57.7 118.38 ;
      RECT 64.34 122.28 64.54 122.4 ;
      RECT 58.58 122.04 58.78 122.16 ;
      RECT 54.62 237.18 54.82 237.3 ;
      RECT 53.9 237.18 54.1 237.3 ;
      RECT 55.34 238.44 55.54 238.56 ;
      RECT 54.62 238.44 54.82 238.56 ;
      RECT 53.9 238.44 54.1 238.56 ;
      RECT 53.54 237.81 53.74 237.93 ;
      RECT 54.98 237.81 55.18 237.93 ;
      RECT 55.34 239.7 55.54 239.82 ;
      RECT 54.62 239.7 54.82 239.82 ;
      RECT 53.9 239.7 54.1 239.82 ;
      RECT 54.98 239.07 55.18 239.19 ;
      RECT 53.54 239.07 53.74 239.19 ;
      RECT 53.54 241.59 53.74 241.71 ;
      RECT 54.98 241.59 55.18 241.71 ;
      RECT 53.9 240.96 54.1 241.08 ;
      RECT 54.62 240.96 54.82 241.08 ;
      RECT 55.34 240.96 55.54 241.08 ;
      RECT 53.54 240.33 53.74 240.45 ;
      RECT 54.98 240.33 55.18 240.45 ;
      RECT 54.98 242.85 55.18 242.97 ;
      RECT 53.54 242.85 53.74 242.97 ;
      RECT 55.34 242.22 55.54 242.34 ;
      RECT 54.62 242.22 54.82 242.34 ;
      RECT 53.9 242.22 54.1 242.34 ;
      RECT 54.98 244.11 55.18 244.23 ;
      RECT 53.54 244.11 53.74 244.23 ;
      RECT 55.34 243.48 55.54 243.6 ;
      RECT 54.62 243.48 54.82 243.6 ;
      RECT 53.9 243.48 54.1 243.6 ;
      RECT 53.54 245.37 53.74 245.49 ;
      RECT 54.98 245.37 55.18 245.49 ;
      RECT 53.9 244.74 54.1 244.86 ;
      RECT 54.62 244.74 54.82 244.86 ;
      RECT 55.34 244.74 55.54 244.86 ;
      RECT 54.98 246.63 55.18 246.75 ;
      RECT 53.54 246.63 53.74 246.75 ;
      RECT 53.9 246 54.1 246.12 ;
      RECT 54.62 246 54.82 246.12 ;
      RECT 55.34 246 55.54 246.12 ;
      RECT 54.98 247.89 55.18 248.01 ;
      RECT 53.54 247.89 53.74 248.01 ;
      RECT 55.34 247.26 55.54 247.38 ;
      RECT 54.62 247.26 54.82 247.38 ;
      RECT 53.9 247.26 54.1 247.38 ;
      RECT 54.62 249.78 54.82 249.9 ;
      RECT 53.9 249.78 54.1 249.9 ;
      RECT 55.34 249.78 55.54 249.9 ;
      RECT 54.98 249.15 55.18 249.27 ;
      RECT 53.54 249.15 53.74 249.27 ;
      RECT 55.34 248.52 55.54 248.64 ;
      RECT 54.62 248.52 54.82 248.64 ;
      RECT 53.9 248.52 54.1 248.64 ;
      RECT 55.34 251.04 55.54 251.16 ;
      RECT 54.62 251.04 54.82 251.16 ;
      RECT 53.9 251.04 54.1 251.16 ;
      RECT 54.98 250.41 55.18 250.53 ;
      RECT 53.54 250.41 53.74 250.53 ;
      RECT 55.34 252.3 55.54 252.42 ;
      RECT 54.62 252.3 54.82 252.42 ;
      RECT 53.9 252.3 54.1 252.42 ;
      RECT 54.98 251.67 55.18 251.79 ;
      RECT 53.54 251.67 53.74 251.79 ;
      RECT 55.34 253.56 55.54 253.68 ;
      RECT 54.62 253.56 54.82 253.68 ;
      RECT 53.9 253.56 54.1 253.68 ;
      RECT 54.98 252.93 55.18 253.05 ;
      RECT 53.54 252.93 53.74 253.05 ;
      RECT 55.34 254.82 55.54 254.94 ;
      RECT 54.62 254.82 54.82 254.94 ;
      RECT 53.9 254.82 54.1 254.94 ;
      RECT 54.98 254.19 55.18 254.31 ;
      RECT 53.54 254.19 53.74 254.31 ;
      RECT 55.34 256.08 55.54 256.2 ;
      RECT 53.9 256.08 54.1 256.2 ;
      RECT 54.62 256.08 54.82 256.2 ;
      RECT 54.98 255.45 55.18 255.57 ;
      RECT 53.54 255.45 53.74 255.57 ;
      RECT 54.98 257.97 55.18 258.09 ;
      RECT 53.54 257.97 53.74 258.09 ;
      RECT 55.34 257.34 55.54 257.46 ;
      RECT 54.62 257.34 54.82 257.46 ;
      RECT 53.9 257.34 54.1 257.46 ;
      RECT 54.98 256.71 55.18 256.83 ;
      RECT 53.54 256.71 53.74 256.83 ;
      RECT 54.98 259.23 55.18 259.35 ;
      RECT 53.54 259.23 53.74 259.35 ;
      RECT 55.34 258.6 55.54 258.72 ;
      RECT 54.62 258.6 54.82 258.72 ;
      RECT 53.9 258.6 54.1 258.72 ;
      RECT 54.98 260.49 55.18 260.61 ;
      RECT 53.54 260.49 53.74 260.61 ;
      RECT 55.34 259.86 55.54 259.98 ;
      RECT 54.62 259.86 54.82 259.98 ;
      RECT 53.9 259.86 54.1 259.98 ;
      RECT 54.98 261.75 55.18 261.87 ;
      RECT 53.54 261.75 53.74 261.87 ;
      RECT 53.9 261.12 54.1 261.24 ;
      RECT 55.34 261.12 55.54 261.24 ;
      RECT 54.62 261.12 54.82 261.24 ;
      RECT 54.98 263.01 55.18 263.13 ;
      RECT 53.54 263.01 53.74 263.13 ;
      RECT 55.34 262.38 55.54 262.5 ;
      RECT 53.54 211.35 53.74 211.47 ;
      RECT 55.34 211.98 55.54 212.1 ;
      RECT 54.62 211.98 54.82 212.1 ;
      RECT 53.9 211.98 54.1 212.1 ;
      RECT 54.98 212.61 55.18 212.73 ;
      RECT 53.54 212.61 53.74 212.73 ;
      RECT 55.34 213.24 55.54 213.36 ;
      RECT 54.62 213.24 54.82 213.36 ;
      RECT 53.9 213.24 54.1 213.36 ;
      RECT 53.54 213.87 53.74 213.99 ;
      RECT 54.98 213.87 55.18 213.99 ;
      RECT 55.34 214.5 55.54 214.62 ;
      RECT 54.62 214.5 54.82 214.62 ;
      RECT 53.9 214.5 54.1 214.62 ;
      RECT 54.98 215.13 55.18 215.25 ;
      RECT 53.54 215.13 53.74 215.25 ;
      RECT 55.34 215.76 55.54 215.88 ;
      RECT 54.62 215.76 54.82 215.88 ;
      RECT 53.9 215.76 54.1 215.88 ;
      RECT 53.54 216.39 53.74 216.51 ;
      RECT 54.98 216.39 55.18 216.51 ;
      RECT 55.34 217.02 55.54 217.14 ;
      RECT 54.62 217.02 54.82 217.14 ;
      RECT 53.9 217.02 54.1 217.14 ;
      RECT 53.54 217.65 53.74 217.77 ;
      RECT 54.98 217.65 55.18 217.77 ;
      RECT 55.34 218.28 55.54 218.4 ;
      RECT 54.62 218.28 54.82 218.4 ;
      RECT 53.9 218.28 54.1 218.4 ;
      RECT 54.98 218.91 55.18 219.03 ;
      RECT 53.54 218.91 53.74 219.03 ;
      RECT 53.9 219.54 54.1 219.66 ;
      RECT 54.62 219.54 54.82 219.66 ;
      RECT 55.34 219.54 55.54 219.66 ;
      RECT 54.98 220.17 55.18 220.29 ;
      RECT 53.54 220.17 53.74 220.29 ;
      RECT 55.34 220.8 55.54 220.92 ;
      RECT 54.62 220.8 54.82 220.92 ;
      RECT 53.9 220.8 54.1 220.92 ;
      RECT 53.54 221.43 53.74 221.55 ;
      RECT 54.98 221.43 55.18 221.55 ;
      RECT 53.9 222.06 54.1 222.18 ;
      RECT 55.34 222.06 55.54 222.18 ;
      RECT 54.62 222.06 54.82 222.18 ;
      RECT 54.98 222.69 55.18 222.81 ;
      RECT 53.54 222.69 53.74 222.81 ;
      RECT 55.34 223.32 55.54 223.44 ;
      RECT 54.62 223.32 54.82 223.44 ;
      RECT 53.9 223.32 54.1 223.44 ;
      RECT 54.98 223.95 55.18 224.07 ;
      RECT 53.54 223.95 53.74 224.07 ;
      RECT 55.34 224.58 55.54 224.7 ;
      RECT 54.62 224.58 54.82 224.7 ;
      RECT 53.9 224.58 54.1 224.7 ;
      RECT 54.98 225.21 55.18 225.33 ;
      RECT 53.54 225.21 53.74 225.33 ;
      RECT 55.34 225.84 55.54 225.96 ;
      RECT 54.62 225.84 54.82 225.96 ;
      RECT 53.9 225.84 54.1 225.96 ;
      RECT 54.98 226.47 55.18 226.59 ;
      RECT 53.54 226.47 53.74 226.59 ;
      RECT 55.34 227.1 55.54 227.22 ;
      RECT 54.62 227.1 54.82 227.22 ;
      RECT 53.9 227.1 54.1 227.22 ;
      RECT 53.54 227.73 53.74 227.85 ;
      RECT 54.98 227.73 55.18 227.85 ;
      RECT 55.34 228.36 55.54 228.48 ;
      RECT 54.62 228.36 54.82 228.48 ;
      RECT 53.9 228.36 54.1 228.48 ;
      RECT 54.98 228.99 55.18 229.11 ;
      RECT 53.54 228.99 53.74 229.11 ;
      RECT 53.9 229.62 54.1 229.74 ;
      RECT 54.62 229.62 54.82 229.74 ;
      RECT 55.34 229.62 55.54 229.74 ;
      RECT 53.54 230.25 53.74 230.37 ;
      RECT 54.98 230.25 55.18 230.37 ;
      RECT 53.9 230.88 54.1 231 ;
      RECT 54.62 230.88 54.82 231 ;
      RECT 55.34 230.88 55.54 231 ;
      RECT 53.54 231.51 53.74 231.63 ;
      RECT 54.98 231.51 55.18 231.63 ;
      RECT 53.9 232.14 54.1 232.26 ;
      RECT 54.62 232.14 54.82 232.26 ;
      RECT 55.34 232.14 55.54 232.26 ;
      RECT 53.54 232.77 53.74 232.89 ;
      RECT 54.98 232.77 55.18 232.89 ;
      RECT 55.34 233.4 55.54 233.52 ;
      RECT 54.62 233.4 54.82 233.52 ;
      RECT 53.9 233.4 54.1 233.52 ;
      RECT 54.98 234.03 55.18 234.15 ;
      RECT 53.54 234.03 53.74 234.15 ;
      RECT 53.9 234.66 54.1 234.78 ;
      RECT 54.62 234.66 54.82 234.78 ;
      RECT 55.34 234.66 55.54 234.78 ;
      RECT 53.54 235.29 53.74 235.41 ;
      RECT 54.98 235.29 55.18 235.41 ;
      RECT 53.9 235.92 54.1 236.04 ;
      RECT 54.62 235.92 54.82 236.04 ;
      RECT 55.34 235.92 55.54 236.04 ;
      RECT 53.54 236.55 53.74 236.67 ;
      RECT 54.98 236.55 55.18 236.67 ;
      RECT 55.34 237.18 55.54 237.3 ;
      RECT 55.34 161.1 55.54 161.22 ;
      RECT 53.9 163.62 54.1 163.74 ;
      RECT 55.34 163.62 55.54 163.74 ;
      RECT 54.26 164.88 54.46 165 ;
      RECT 54.62 163.86 54.82 163.98 ;
      RECT 55.34 166.38 55.54 166.5 ;
      RECT 53.9 166.38 54.1 166.5 ;
      RECT 54.62 166.14 54.82 166.26 ;
      RECT 54.26 167.4 54.46 167.52 ;
      RECT 55.34 168.9 55.54 169.02 ;
      RECT 54.62 168.9 54.82 169.02 ;
      RECT 53.9 168.66 54.1 168.78 ;
      RECT 54.26 169.92 54.46 170.04 ;
      RECT 54.62 171.42 54.82 171.54 ;
      RECT 53.9 171.18 54.1 171.3 ;
      RECT 55.34 171.18 55.54 171.3 ;
      RECT 54.26 172.44 54.46 172.56 ;
      RECT 53.9 173.94 54.1 174.06 ;
      RECT 54.62 173.7 54.82 173.82 ;
      RECT 55.34 173.7 55.54 173.82 ;
      RECT 54.26 175.2 54.46 175.32 ;
      RECT 55.34 176.46 55.54 176.58 ;
      RECT 54.62 176.46 54.82 176.58 ;
      RECT 53.9 176.22 54.1 176.34 ;
      RECT 55.34 178.74 55.54 178.86 ;
      RECT 53.9 178.74 54.1 178.86 ;
      RECT 54.26 177.48 54.46 177.6 ;
      RECT 54.26 180 54.46 180.12 ;
      RECT 54.62 178.98 54.82 179.1 ;
      RECT 53.9 181.5 54.1 181.62 ;
      RECT 55.34 181.26 55.54 181.38 ;
      RECT 54.62 181.26 54.82 181.38 ;
      RECT 54.26 182.76 54.46 182.88 ;
      RECT 54.62 184.02 54.82 184.14 ;
      RECT 55.34 183.78 55.54 183.9 ;
      RECT 53.9 183.78 54.1 183.9 ;
      RECT 54.26 185.28 54.46 185.4 ;
      RECT 54.62 186.54 54.82 186.66 ;
      RECT 55.34 186.3 55.54 186.42 ;
      RECT 53.9 186.3 54.1 186.42 ;
      RECT 54.26 187.8 54.46 187.92 ;
      RECT 53.9 189.06 54.1 189.18 ;
      RECT 54.62 189.06 54.82 189.18 ;
      RECT 55.34 188.82 55.54 188.94 ;
      RECT 53.54 190.862 53.74 190.982 ;
      RECT 54.98 190.622 55.18 190.742 ;
      RECT 54.26 190.08 54.46 190.2 ;
      RECT 53.54 191.882 53.74 192.002 ;
      RECT 54.98 191.882 55.18 192.002 ;
      RECT 55.34 191.58 55.54 191.7 ;
      RECT 53.9 191.58 54.1 191.7 ;
      RECT 54.62 191.34 54.82 191.46 ;
      RECT 53.54 193.382 53.74 193.502 ;
      RECT 54.98 193.142 55.18 193.262 ;
      RECT 54.26 192.6 54.46 192.72 ;
      RECT 54.98 194.402 55.18 194.522 ;
      RECT 53.54 194.402 53.74 194.522 ;
      RECT 53.9 193.86 54.1 193.98 ;
      RECT 54.62 193.86 54.82 193.98 ;
      RECT 55.34 193.86 55.54 193.98 ;
      RECT 54.26 195.12 54.46 195.24 ;
      RECT 53.54 195.662 53.74 195.782 ;
      RECT 54.98 195.662 55.18 195.782 ;
      RECT 55.34 196.38 55.54 196.5 ;
      RECT 53.9 196.38 54.1 196.5 ;
      RECT 54.62 196.62 54.82 196.74 ;
      RECT 54.26 197.88 54.46 198 ;
      RECT 54.98 198.182 55.18 198.302 ;
      RECT 53.54 198.422 53.74 198.542 ;
      RECT 53.9 198.9 54.1 199.02 ;
      RECT 55.34 198.9 55.54 199.02 ;
      RECT 54.62 199.14 54.82 199.26 ;
      RECT 54.26 200.4 54.46 200.52 ;
      RECT 53.54 200.942 53.74 201.062 ;
      RECT 54.98 200.942 55.18 201.062 ;
      RECT 55.34 201.42 55.54 201.54 ;
      RECT 53.9 201.66 54.1 201.78 ;
      RECT 54.62 201.66 54.82 201.78 ;
      RECT 54.26 202.68 54.46 202.8 ;
      RECT 53.54 203.222 53.74 203.342 ;
      RECT 54.98 203.462 55.18 203.582 ;
      RECT 54.62 203.94 54.82 204.06 ;
      RECT 55.34 204.18 55.54 204.3 ;
      RECT 53.9 204.18 54.1 204.3 ;
      RECT 54.26 205.44 54.46 205.56 ;
      RECT 54.98 205.742 55.18 205.862 ;
      RECT 53.54 205.982 53.74 206.102 ;
      RECT 53.9 206.46 54.1 206.58 ;
      RECT 54.62 206.46 54.82 206.58 ;
      RECT 55.34 206.7 55.54 206.82 ;
      RECT 54.26 207.72 54.46 207.84 ;
      RECT 54.98 208.262 55.18 208.382 ;
      RECT 53.54 208.502 53.74 208.622 ;
      RECT 53.9 209.46 54.1 209.58 ;
      RECT 54.62 209.46 54.82 209.58 ;
      RECT 55.34 209.46 55.54 209.58 ;
      RECT 54.98 210.09 55.18 210.21 ;
      RECT 53.54 210.09 53.74 210.21 ;
      RECT 55.34 210.72 55.54 210.84 ;
      RECT 54.62 210.72 54.82 210.84 ;
      RECT 53.9 210.72 54.1 210.84 ;
      RECT 54.98 211.35 55.18 211.47 ;
      RECT 52.82 348.339 53.02 348.459 ;
      RECT 55.34 118.5 55.54 118.62 ;
      RECT 53.9 118.5 54.1 118.62 ;
      RECT 54.62 118.26 54.82 118.38 ;
      RECT 54.26 119.76 54.46 119.88 ;
      RECT 53.9 118.978 54.1 119.098 ;
      RECT 54.62 118.978 54.82 119.098 ;
      RECT 55.34 118.978 55.54 119.098 ;
      RECT 53.9 121.02 54.1 121.14 ;
      RECT 55.34 121.02 55.54 121.14 ;
      RECT 54.62 120.78 54.82 120.9 ;
      RECT 54.26 122.28 54.46 122.4 ;
      RECT 53.9 121.498 54.1 121.618 ;
      RECT 54.62 121.498 54.82 121.618 ;
      RECT 55.34 121.498 55.54 121.618 ;
      RECT 53.9 124.018 54.1 124.138 ;
      RECT 54.62 124.018 54.82 124.138 ;
      RECT 55.34 124.018 55.54 124.138 ;
      RECT 54.62 123.54 54.82 123.66 ;
      RECT 53.9 123.3 54.1 123.42 ;
      RECT 55.34 123.3 55.54 123.42 ;
      RECT 54.26 124.8 54.46 124.92 ;
      RECT 53.9 126.538 54.1 126.658 ;
      RECT 54.62 126.538 54.82 126.658 ;
      RECT 55.34 126.538 55.54 126.658 ;
      RECT 54.62 126.06 54.82 126.18 ;
      RECT 53.9 125.82 54.1 125.94 ;
      RECT 55.34 125.82 55.54 125.94 ;
      RECT 54.26 127.32 54.46 127.44 ;
      RECT 54.26 129.6 54.46 129.72 ;
      RECT 53.9 129.058 54.1 129.178 ;
      RECT 54.62 129.058 54.82 129.178 ;
      RECT 55.34 129.058 55.54 129.178 ;
      RECT 54.62 128.58 54.82 128.7 ;
      RECT 53.9 128.58 54.1 128.7 ;
      RECT 55.34 128.34 55.54 128.46 ;
      RECT 53.9 130.86 54.1 130.98 ;
      RECT 55.34 130.86 55.54 130.98 ;
      RECT 54.26 132.12 54.46 132.24 ;
      RECT 53.9 131.578 54.1 131.698 ;
      RECT 54.62 131.578 54.82 131.698 ;
      RECT 55.34 131.578 55.54 131.698 ;
      RECT 54.62 131.1 54.82 131.22 ;
      RECT 55.34 133.62 55.54 133.74 ;
      RECT 54.62 133.38 54.82 133.5 ;
      RECT 53.9 133.38 54.1 133.5 ;
      RECT 54.26 134.64 54.46 134.76 ;
      RECT 53.9 134.098 54.1 134.218 ;
      RECT 54.62 134.098 54.82 134.218 ;
      RECT 55.34 134.098 55.54 134.218 ;
      RECT 54.62 136.14 54.82 136.26 ;
      RECT 55.34 135.9 55.54 136.02 ;
      RECT 53.9 135.9 54.1 136.02 ;
      RECT 54.26 137.16 54.46 137.28 ;
      RECT 53.9 136.618 54.1 136.738 ;
      RECT 54.62 136.618 54.82 136.738 ;
      RECT 55.34 136.618 55.54 136.738 ;
      RECT 53.9 139.138 54.1 139.258 ;
      RECT 54.62 139.138 54.82 139.258 ;
      RECT 55.34 139.138 55.54 139.258 ;
      RECT 54.62 138.66 54.82 138.78 ;
      RECT 55.34 138.42 55.54 138.54 ;
      RECT 53.9 138.42 54.1 138.54 ;
      RECT 54.26 139.68 54.46 139.8 ;
      RECT 53.9 141.18 54.1 141.3 ;
      RECT 54.62 140.94 54.82 141.06 ;
      RECT 55.34 140.94 55.54 141.06 ;
      RECT 54.26 142.44 54.46 142.56 ;
      RECT 55.34 143.7 55.54 143.82 ;
      RECT 53.9 143.7 54.1 143.82 ;
      RECT 54.62 143.46 54.82 143.58 ;
      RECT 53.9 145.98 54.1 146.1 ;
      RECT 54.62 145.98 54.82 146.1 ;
      RECT 55.34 145.98 55.54 146.1 ;
      RECT 54.26 144.72 54.46 144.84 ;
      RECT 53.9 148.74 54.1 148.86 ;
      RECT 55.34 148.5 55.54 148.62 ;
      RECT 54.62 148.5 54.82 148.62 ;
      RECT 54.26 150 54.46 150.12 ;
      RECT 53.9 151.26 54.1 151.38 ;
      RECT 54.62 151.26 54.82 151.38 ;
      RECT 55.34 151.02 55.54 151.14 ;
      RECT 54.26 152.28 54.46 152.4 ;
      RECT 54.62 153.78 54.82 153.9 ;
      RECT 53.9 153.78 54.1 153.9 ;
      RECT 55.34 153.54 55.54 153.66 ;
      RECT 54.26 154.8 54.46 154.92 ;
      RECT 54.98 156.842 55.18 156.962 ;
      RECT 53.54 156.602 53.74 156.722 ;
      RECT 53.9 156.3 54.1 156.42 ;
      RECT 54.62 156.3 54.82 156.42 ;
      RECT 55.34 156.06 55.54 156.18 ;
      RECT 53.54 158.278 53.74 158.398 ;
      RECT 54.98 158.038 55.18 158.158 ;
      RECT 54.26 157.32 54.46 157.44 ;
      RECT 53.9 158.82 54.1 158.94 ;
      RECT 54.62 158.82 54.82 158.94 ;
      RECT 55.34 158.58 55.54 158.7 ;
      RECT 54.26 159.84 54.46 159.96 ;
      RECT 54.26 162.36 54.46 162.48 ;
      RECT 53.9 161.1 54.1 161.22 ;
      RECT 54.62 161.1 54.82 161.22 ;
      RECT 52.1 261.75 52.3 261.87 ;
      RECT 49.22 261.75 49.42 261.87 ;
      RECT 52.46 261.12 52.66 261.24 ;
      RECT 53.18 261.12 53.38 261.24 ;
      RECT 51.74 261.12 51.94 261.24 ;
      RECT 49.58 261.12 49.78 261.24 ;
      RECT 52.1 263.01 52.3 263.13 ;
      RECT 49.22 263.01 49.42 263.13 ;
      RECT 53.18 262.38 53.38 262.5 ;
      RECT 52.46 262.38 52.66 262.5 ;
      RECT 51.74 262.38 51.94 262.5 ;
      RECT 49.58 262.38 49.78 262.5 ;
      RECT 52.1 264.27 52.3 264.39 ;
      RECT 49.22 264.27 49.42 264.39 ;
      RECT 53.18 263.64 53.38 263.76 ;
      RECT 52.46 263.64 52.66 263.76 ;
      RECT 51.74 263.64 51.94 263.76 ;
      RECT 49.58 263.64 49.78 263.76 ;
      RECT 53.18 266.16 53.38 266.28 ;
      RECT 52.46 266.16 52.66 266.28 ;
      RECT 51.74 266.16 51.94 266.28 ;
      RECT 49.58 266.16 49.78 266.28 ;
      RECT 52.1 265.53 52.3 265.65 ;
      RECT 49.22 265.53 49.42 265.65 ;
      RECT 53.18 264.9 53.38 265.02 ;
      RECT 52.46 264.9 52.66 265.02 ;
      RECT 51.74 264.9 51.94 265.02 ;
      RECT 49.58 264.9 49.78 265.02 ;
      RECT 53.18 267.42 53.38 267.54 ;
      RECT 52.46 267.42 52.66 267.54 ;
      RECT 51.74 267.42 51.94 267.54 ;
      RECT 49.58 267.42 49.78 267.54 ;
      RECT 52.1 266.79 52.3 266.91 ;
      RECT 49.22 266.79 49.42 266.91 ;
      RECT 53.18 268.68 53.38 268.8 ;
      RECT 52.46 268.68 52.66 268.8 ;
      RECT 51.74 268.68 51.94 268.8 ;
      RECT 49.58 268.68 49.78 268.8 ;
      RECT 52.1 268.05 52.3 268.17 ;
      RECT 49.22 268.05 49.42 268.17 ;
      RECT 53.18 269.94 53.38 270.06 ;
      RECT 52.46 269.94 52.66 270.06 ;
      RECT 51.74 269.94 51.94 270.06 ;
      RECT 49.58 269.94 49.78 270.06 ;
      RECT 52.1 269.31 52.3 269.43 ;
      RECT 49.22 269.31 49.42 269.43 ;
      RECT 53.18 271.2 53.38 271.32 ;
      RECT 52.46 271.2 52.66 271.32 ;
      RECT 51.74 271.2 51.94 271.32 ;
      RECT 49.58 271.2 49.78 271.32 ;
      RECT 52.1 270.57 52.3 270.69 ;
      RECT 49.22 270.57 49.42 270.69 ;
      RECT 53.18 272.46 53.38 272.58 ;
      RECT 52.46 272.46 52.66 272.58 ;
      RECT 51.74 272.46 51.94 272.58 ;
      RECT 49.58 272.46 49.78 272.58 ;
      RECT 52.1 271.83 52.3 271.95 ;
      RECT 49.22 271.83 49.42 271.95 ;
      RECT 52.1 274.35 52.3 274.47 ;
      RECT 49.22 274.35 49.42 274.47 ;
      RECT 53.18 273.72 53.38 273.84 ;
      RECT 52.46 273.72 52.66 273.84 ;
      RECT 51.74 273.72 51.94 273.84 ;
      RECT 49.58 273.72 49.78 273.84 ;
      RECT 49.22 273.09 49.42 273.21 ;
      RECT 52.1 273.09 52.3 273.21 ;
      RECT 52.1 275.61 52.3 275.73 ;
      RECT 49.22 275.61 49.42 275.73 ;
      RECT 53.18 274.98 53.38 275.1 ;
      RECT 52.46 274.98 52.66 275.1 ;
      RECT 51.74 274.98 51.94 275.1 ;
      RECT 49.58 274.98 49.78 275.1 ;
      RECT 52.1 276.87 52.3 276.99 ;
      RECT 49.22 276.87 49.42 276.99 ;
      RECT 53.18 276.24 53.38 276.36 ;
      RECT 52.46 276.24 52.66 276.36 ;
      RECT 51.74 276.24 51.94 276.36 ;
      RECT 49.58 276.24 49.78 276.36 ;
      RECT 52.1 278.13 52.3 278.25 ;
      RECT 49.22 278.13 49.42 278.25 ;
      RECT 53.18 277.5 53.38 277.62 ;
      RECT 52.46 277.5 52.66 277.62 ;
      RECT 51.74 277.5 51.94 277.62 ;
      RECT 49.58 277.5 49.78 277.62 ;
      RECT 53.18 278.76 53.38 278.88 ;
      RECT 51.74 278.76 51.94 278.88 ;
      RECT 52.46 278.76 52.66 278.88 ;
      RECT 49.58 278.76 49.78 278.88 ;
      RECT 52.46 283.087 52.66 283.207 ;
      RECT 51.74 283.087 51.94 283.207 ;
      RECT 49.58 283.087 49.78 283.207 ;
      RECT 53.18 283.087 53.38 283.207 ;
      RECT 52.82 305.498 53.02 305.618 ;
      RECT 51.74 305.967 51.94 306.087 ;
      RECT 53.18 305.967 53.38 306.087 ;
      RECT 52.46 305.967 52.66 306.087 ;
      RECT 49.58 305.967 49.78 306.087 ;
      RECT 52.82 323.3835 53.02 323.5035 ;
      RECT 53.18 325.9425 53.38 326.0625 ;
      RECT 49.58 325.9425 49.78 326.0625 ;
      RECT 51.74 325.9425 51.94 326.0625 ;
      RECT 52.46 325.9425 52.66 326.0625 ;
      RECT 51.74 239.7 51.94 239.82 ;
      RECT 49.58 239.7 49.78 239.82 ;
      RECT 52.1 239.07 52.3 239.19 ;
      RECT 49.22 239.07 49.42 239.19 ;
      RECT 49.22 241.59 49.42 241.71 ;
      RECT 52.1 241.59 52.3 241.71 ;
      RECT 53.18 240.96 53.38 241.08 ;
      RECT 52.46 240.96 52.66 241.08 ;
      RECT 51.74 240.96 51.94 241.08 ;
      RECT 49.58 240.96 49.78 241.08 ;
      RECT 52.1 240.33 52.3 240.45 ;
      RECT 49.22 240.33 49.42 240.45 ;
      RECT 52.1 242.85 52.3 242.97 ;
      RECT 49.22 242.85 49.42 242.97 ;
      RECT 53.18 242.22 53.38 242.34 ;
      RECT 52.46 242.22 52.66 242.34 ;
      RECT 51.74 242.22 51.94 242.34 ;
      RECT 49.58 242.22 49.78 242.34 ;
      RECT 52.1 244.11 52.3 244.23 ;
      RECT 49.22 244.11 49.42 244.23 ;
      RECT 53.18 243.48 53.38 243.6 ;
      RECT 52.46 243.48 52.66 243.6 ;
      RECT 51.74 243.48 51.94 243.6 ;
      RECT 49.58 243.48 49.78 243.6 ;
      RECT 49.22 245.37 49.42 245.49 ;
      RECT 52.1 245.37 52.3 245.49 ;
      RECT 49.58 244.74 49.78 244.86 ;
      RECT 51.74 244.74 51.94 244.86 ;
      RECT 52.46 244.74 52.66 244.86 ;
      RECT 53.18 244.74 53.38 244.86 ;
      RECT 52.1 246.63 52.3 246.75 ;
      RECT 49.22 246.63 49.42 246.75 ;
      RECT 49.58 246 49.78 246.12 ;
      RECT 51.74 246 51.94 246.12 ;
      RECT 52.46 246 52.66 246.12 ;
      RECT 53.18 246 53.38 246.12 ;
      RECT 52.1 247.89 52.3 248.01 ;
      RECT 49.22 247.89 49.42 248.01 ;
      RECT 53.18 247.26 53.38 247.38 ;
      RECT 52.46 247.26 52.66 247.38 ;
      RECT 51.74 247.26 51.94 247.38 ;
      RECT 49.58 247.26 49.78 247.38 ;
      RECT 53.18 249.78 53.38 249.9 ;
      RECT 52.46 249.78 52.66 249.9 ;
      RECT 51.74 249.78 51.94 249.9 ;
      RECT 49.58 249.78 49.78 249.9 ;
      RECT 52.1 249.15 52.3 249.27 ;
      RECT 49.22 249.15 49.42 249.27 ;
      RECT 53.18 248.52 53.38 248.64 ;
      RECT 52.46 248.52 52.66 248.64 ;
      RECT 51.74 248.52 51.94 248.64 ;
      RECT 49.58 248.52 49.78 248.64 ;
      RECT 53.18 251.04 53.38 251.16 ;
      RECT 52.46 251.04 52.66 251.16 ;
      RECT 51.74 251.04 51.94 251.16 ;
      RECT 49.58 251.04 49.78 251.16 ;
      RECT 52.1 250.41 52.3 250.53 ;
      RECT 49.22 250.41 49.42 250.53 ;
      RECT 53.18 252.3 53.38 252.42 ;
      RECT 52.46 252.3 52.66 252.42 ;
      RECT 51.74 252.3 51.94 252.42 ;
      RECT 49.58 252.3 49.78 252.42 ;
      RECT 52.1 251.67 52.3 251.79 ;
      RECT 49.22 251.67 49.42 251.79 ;
      RECT 53.18 253.56 53.38 253.68 ;
      RECT 52.46 253.56 52.66 253.68 ;
      RECT 51.74 253.56 51.94 253.68 ;
      RECT 49.58 253.56 49.78 253.68 ;
      RECT 52.1 252.93 52.3 253.05 ;
      RECT 49.22 252.93 49.42 253.05 ;
      RECT 53.18 254.82 53.38 254.94 ;
      RECT 52.46 254.82 52.66 254.94 ;
      RECT 51.74 254.82 51.94 254.94 ;
      RECT 49.58 254.82 49.78 254.94 ;
      RECT 52.1 254.19 52.3 254.31 ;
      RECT 49.22 254.19 49.42 254.31 ;
      RECT 53.18 256.08 53.38 256.2 ;
      RECT 52.46 256.08 52.66 256.2 ;
      RECT 51.74 256.08 51.94 256.2 ;
      RECT 49.58 256.08 49.78 256.2 ;
      RECT 52.1 255.45 52.3 255.57 ;
      RECT 49.22 255.45 49.42 255.57 ;
      RECT 52.1 257.97 52.3 258.09 ;
      RECT 49.22 257.97 49.42 258.09 ;
      RECT 53.18 257.34 53.38 257.46 ;
      RECT 52.46 257.34 52.66 257.46 ;
      RECT 51.74 257.34 51.94 257.46 ;
      RECT 49.58 257.34 49.78 257.46 ;
      RECT 52.1 256.71 52.3 256.83 ;
      RECT 49.22 256.71 49.42 256.83 ;
      RECT 52.1 259.23 52.3 259.35 ;
      RECT 49.22 259.23 49.42 259.35 ;
      RECT 53.18 258.6 53.38 258.72 ;
      RECT 52.46 258.6 52.66 258.72 ;
      RECT 51.74 258.6 51.94 258.72 ;
      RECT 49.58 258.6 49.78 258.72 ;
      RECT 52.1 260.49 52.3 260.61 ;
      RECT 49.22 260.49 49.42 260.61 ;
      RECT 53.18 259.86 53.38 259.98 ;
      RECT 52.46 259.86 52.66 259.98 ;
      RECT 51.74 259.86 51.94 259.98 ;
      RECT 49.58 259.86 49.78 259.98 ;
      RECT 53.18 218.28 53.38 218.4 ;
      RECT 52.46 218.28 52.66 218.4 ;
      RECT 51.74 218.28 51.94 218.4 ;
      RECT 49.58 218.28 49.78 218.4 ;
      RECT 52.1 218.91 52.3 219.03 ;
      RECT 49.22 218.91 49.42 219.03 ;
      RECT 49.58 219.54 49.78 219.66 ;
      RECT 51.74 219.54 51.94 219.66 ;
      RECT 52.46 219.54 52.66 219.66 ;
      RECT 53.18 219.54 53.38 219.66 ;
      RECT 52.1 220.17 52.3 220.29 ;
      RECT 49.22 220.17 49.42 220.29 ;
      RECT 53.18 220.8 53.38 220.92 ;
      RECT 52.46 220.8 52.66 220.92 ;
      RECT 51.74 220.8 51.94 220.92 ;
      RECT 49.58 220.8 49.78 220.92 ;
      RECT 49.22 221.43 49.42 221.55 ;
      RECT 52.1 221.43 52.3 221.55 ;
      RECT 53.18 222.06 53.38 222.18 ;
      RECT 52.46 222.06 52.66 222.18 ;
      RECT 51.74 222.06 51.94 222.18 ;
      RECT 49.58 222.06 49.78 222.18 ;
      RECT 52.1 222.69 52.3 222.81 ;
      RECT 49.22 222.69 49.42 222.81 ;
      RECT 53.18 223.32 53.38 223.44 ;
      RECT 52.46 223.32 52.66 223.44 ;
      RECT 51.74 223.32 51.94 223.44 ;
      RECT 49.58 223.32 49.78 223.44 ;
      RECT 52.1 223.95 52.3 224.07 ;
      RECT 49.22 223.95 49.42 224.07 ;
      RECT 53.18 224.58 53.38 224.7 ;
      RECT 52.46 224.58 52.66 224.7 ;
      RECT 51.74 224.58 51.94 224.7 ;
      RECT 49.58 224.58 49.78 224.7 ;
      RECT 52.1 225.21 52.3 225.33 ;
      RECT 49.22 225.21 49.42 225.33 ;
      RECT 53.18 225.84 53.38 225.96 ;
      RECT 52.46 225.84 52.66 225.96 ;
      RECT 51.74 225.84 51.94 225.96 ;
      RECT 49.58 225.84 49.78 225.96 ;
      RECT 52.1 226.47 52.3 226.59 ;
      RECT 49.22 226.47 49.42 226.59 ;
      RECT 53.18 227.1 53.38 227.22 ;
      RECT 52.46 227.1 52.66 227.22 ;
      RECT 51.74 227.1 51.94 227.22 ;
      RECT 49.58 227.1 49.78 227.22 ;
      RECT 49.22 227.73 49.42 227.85 ;
      RECT 52.1 227.73 52.3 227.85 ;
      RECT 53.18 228.36 53.38 228.48 ;
      RECT 52.46 228.36 52.66 228.48 ;
      RECT 51.74 228.36 51.94 228.48 ;
      RECT 49.58 228.36 49.78 228.48 ;
      RECT 52.1 228.99 52.3 229.11 ;
      RECT 49.22 228.99 49.42 229.11 ;
      RECT 49.58 229.62 49.78 229.74 ;
      RECT 51.74 229.62 51.94 229.74 ;
      RECT 52.46 229.62 52.66 229.74 ;
      RECT 53.18 229.62 53.38 229.74 ;
      RECT 49.22 230.25 49.42 230.37 ;
      RECT 52.1 230.25 52.3 230.37 ;
      RECT 49.58 230.88 49.78 231 ;
      RECT 51.74 230.88 51.94 231 ;
      RECT 52.46 230.88 52.66 231 ;
      RECT 53.18 230.88 53.38 231 ;
      RECT 49.22 231.51 49.42 231.63 ;
      RECT 52.1 231.51 52.3 231.63 ;
      RECT 49.58 232.14 49.78 232.26 ;
      RECT 51.74 232.14 51.94 232.26 ;
      RECT 52.46 232.14 52.66 232.26 ;
      RECT 53.18 232.14 53.38 232.26 ;
      RECT 49.22 232.77 49.42 232.89 ;
      RECT 52.1 232.77 52.3 232.89 ;
      RECT 53.18 233.4 53.38 233.52 ;
      RECT 52.46 233.4 52.66 233.52 ;
      RECT 51.74 233.4 51.94 233.52 ;
      RECT 49.58 233.4 49.78 233.52 ;
      RECT 52.1 234.03 52.3 234.15 ;
      RECT 49.22 234.03 49.42 234.15 ;
      RECT 49.58 234.66 49.78 234.78 ;
      RECT 51.74 234.66 51.94 234.78 ;
      RECT 52.46 234.66 52.66 234.78 ;
      RECT 53.18 234.66 53.38 234.78 ;
      RECT 49.22 235.29 49.42 235.41 ;
      RECT 52.1 235.29 52.3 235.41 ;
      RECT 49.58 235.92 49.78 236.04 ;
      RECT 51.74 235.92 51.94 236.04 ;
      RECT 52.46 235.92 52.66 236.04 ;
      RECT 53.18 235.92 53.38 236.04 ;
      RECT 49.58 237.18 49.78 237.3 ;
      RECT 51.74 237.18 51.94 237.3 ;
      RECT 52.46 237.18 52.66 237.3 ;
      RECT 53.18 237.18 53.38 237.3 ;
      RECT 49.22 236.55 49.42 236.67 ;
      RECT 52.1 236.55 52.3 236.67 ;
      RECT 53.18 238.44 53.38 238.56 ;
      RECT 52.46 238.44 52.66 238.56 ;
      RECT 51.74 238.44 51.94 238.56 ;
      RECT 49.58 238.44 49.78 238.56 ;
      RECT 49.22 237.81 49.42 237.93 ;
      RECT 52.1 237.81 52.3 237.93 ;
      RECT 53.18 239.7 53.38 239.82 ;
      RECT 52.46 239.7 52.66 239.82 ;
      RECT 51.74 189.06 51.94 189.18 ;
      RECT 52.46 189.06 52.66 189.18 ;
      RECT 53.18 189.06 53.38 189.18 ;
      RECT 49.58 188.82 49.78 188.94 ;
      RECT 49.22 190.622 49.42 190.742 ;
      RECT 52.1 190.622 52.3 190.742 ;
      RECT 52.82 190.08 53.02 190.2 ;
      RECT 49.22 192.122 49.42 192.242 ;
      RECT 52.1 191.882 52.3 192.002 ;
      RECT 53.18 191.58 53.38 191.7 ;
      RECT 49.58 191.34 49.78 191.46 ;
      RECT 51.74 191.34 51.94 191.46 ;
      RECT 52.46 191.34 52.66 191.46 ;
      RECT 49.22 193.382 49.42 193.502 ;
      RECT 52.1 193.142 52.3 193.262 ;
      RECT 52.82 192.84 53.02 192.96 ;
      RECT 49.22 194.642 49.42 194.762 ;
      RECT 52.1 194.642 52.3 194.762 ;
      RECT 52.46 194.1 52.66 194.22 ;
      RECT 49.58 193.86 49.78 193.98 ;
      RECT 51.74 193.86 51.94 193.98 ;
      RECT 53.18 193.86 53.38 193.98 ;
      RECT 52.82 195.36 53.02 195.48 ;
      RECT 49.22 195.662 49.42 195.782 ;
      RECT 52.1 195.902 52.3 196.022 ;
      RECT 53.18 196.38 53.38 196.5 ;
      RECT 52.46 196.38 52.66 196.5 ;
      RECT 49.58 196.38 49.78 196.5 ;
      RECT 51.74 196.62 51.94 196.74 ;
      RECT 52.82 197.88 53.02 198 ;
      RECT 52.1 198.182 52.3 198.302 ;
      RECT 49.22 198.182 49.42 198.302 ;
      RECT 51.74 198.9 51.94 199.02 ;
      RECT 52.46 198.9 52.66 199.02 ;
      RECT 53.18 199.14 53.38 199.26 ;
      RECT 49.58 199.14 49.78 199.26 ;
      RECT 52.82 200.16 53.02 200.28 ;
      RECT 49.22 200.702 49.42 200.822 ;
      RECT 52.1 200.942 52.3 201.062 ;
      RECT 52.46 201.42 52.66 201.54 ;
      RECT 51.74 201.42 51.94 201.54 ;
      RECT 49.58 201.42 49.78 201.54 ;
      RECT 53.18 201.66 53.38 201.78 ;
      RECT 52.82 202.92 53.02 203.04 ;
      RECT 49.22 203.462 49.42 203.582 ;
      RECT 52.1 203.462 52.3 203.582 ;
      RECT 52.46 203.94 52.66 204.06 ;
      RECT 53.18 203.94 53.38 204.06 ;
      RECT 51.74 204.18 51.94 204.3 ;
      RECT 49.58 204.18 49.78 204.3 ;
      RECT 52.82 205.44 53.02 205.56 ;
      RECT 52.1 205.742 52.3 205.862 ;
      RECT 49.22 205.982 49.42 206.102 ;
      RECT 49.58 206.46 49.78 206.58 ;
      RECT 52.46 206.46 52.66 206.58 ;
      RECT 51.74 206.7 51.94 206.82 ;
      RECT 53.18 206.7 53.38 206.82 ;
      RECT 52.82 207.96 53.02 208.08 ;
      RECT 49.22 208.262 49.42 208.382 ;
      RECT 52.1 208.502 52.3 208.622 ;
      RECT 49.58 209.46 49.78 209.58 ;
      RECT 51.74 209.46 51.94 209.58 ;
      RECT 52.46 209.46 52.66 209.58 ;
      RECT 53.18 209.46 53.38 209.58 ;
      RECT 52.1 210.09 52.3 210.21 ;
      RECT 49.22 210.09 49.42 210.21 ;
      RECT 53.18 210.72 53.38 210.84 ;
      RECT 52.46 210.72 52.66 210.84 ;
      RECT 51.74 210.72 51.94 210.84 ;
      RECT 49.58 210.72 49.78 210.84 ;
      RECT 52.1 211.35 52.3 211.47 ;
      RECT 49.22 211.35 49.42 211.47 ;
      RECT 53.18 211.98 53.38 212.1 ;
      RECT 52.46 211.98 52.66 212.1 ;
      RECT 51.74 211.98 51.94 212.1 ;
      RECT 49.58 211.98 49.78 212.1 ;
      RECT 52.1 212.61 52.3 212.73 ;
      RECT 49.22 212.61 49.42 212.73 ;
      RECT 53.18 213.24 53.38 213.36 ;
      RECT 52.46 213.24 52.66 213.36 ;
      RECT 51.74 213.24 51.94 213.36 ;
      RECT 49.58 213.24 49.78 213.36 ;
      RECT 49.22 213.87 49.42 213.99 ;
      RECT 52.1 213.87 52.3 213.99 ;
      RECT 53.18 214.5 53.38 214.62 ;
      RECT 52.46 214.5 52.66 214.62 ;
      RECT 51.74 214.5 51.94 214.62 ;
      RECT 49.58 214.5 49.78 214.62 ;
      RECT 52.1 215.13 52.3 215.25 ;
      RECT 49.22 215.13 49.42 215.25 ;
      RECT 53.18 215.76 53.38 215.88 ;
      RECT 52.46 215.76 52.66 215.88 ;
      RECT 51.74 215.76 51.94 215.88 ;
      RECT 49.58 215.76 49.78 215.88 ;
      RECT 49.22 216.39 49.42 216.51 ;
      RECT 52.1 216.39 52.3 216.51 ;
      RECT 53.18 217.02 53.38 217.14 ;
      RECT 52.46 217.02 52.66 217.14 ;
      RECT 51.74 217.02 51.94 217.14 ;
      RECT 49.58 217.02 49.78 217.14 ;
      RECT 52.1 217.65 52.3 217.77 ;
      RECT 49.22 217.65 49.42 217.77 ;
      RECT 52.46 138.66 52.66 138.78 ;
      RECT 49.58 138.66 49.78 138.78 ;
      RECT 51.74 138.42 51.94 138.54 ;
      RECT 52.82 139.92 53.02 140.04 ;
      RECT 53.18 141.18 53.38 141.3 ;
      RECT 52.46 141.18 52.66 141.3 ;
      RECT 49.58 141.18 49.78 141.3 ;
      RECT 51.74 140.94 51.94 141.06 ;
      RECT 52.82 142.2 53.02 142.32 ;
      RECT 52.46 143.7 52.66 143.82 ;
      RECT 51.74 143.7 51.94 143.82 ;
      RECT 53.18 143.46 53.38 143.58 ;
      RECT 49.58 143.46 49.78 143.58 ;
      RECT 49.58 145.98 49.78 146.1 ;
      RECT 51.74 145.98 51.94 146.1 ;
      RECT 52.46 145.98 52.66 146.1 ;
      RECT 53.18 145.98 53.38 146.1 ;
      RECT 52.82 144.96 53.02 145.08 ;
      RECT 49.58 148.74 49.78 148.86 ;
      RECT 52.46 148.74 52.66 148.86 ;
      RECT 53.18 148.74 53.38 148.86 ;
      RECT 51.74 148.5 51.94 148.62 ;
      RECT 52.82 149.76 53.02 149.88 ;
      RECT 49.58 151.26 49.78 151.38 ;
      RECT 52.46 151.26 52.66 151.38 ;
      RECT 53.18 151.02 53.38 151.14 ;
      RECT 51.74 151.02 51.94 151.14 ;
      RECT 52.82 152.52 53.02 152.64 ;
      RECT 53.18 153.78 53.38 153.9 ;
      RECT 52.46 153.78 52.66 153.9 ;
      RECT 51.74 153.78 51.94 153.9 ;
      RECT 49.58 153.78 49.78 153.9 ;
      RECT 52.82 154.8 53.02 154.92 ;
      RECT 52.1 156.842 52.3 156.962 ;
      RECT 49.22 156.602 49.42 156.722 ;
      RECT 52.46 156.3 52.66 156.42 ;
      RECT 53.18 156.06 53.38 156.18 ;
      RECT 51.74 156.06 51.94 156.18 ;
      RECT 49.58 156.06 49.78 156.18 ;
      RECT 49.22 158.278 49.42 158.398 ;
      RECT 52.1 158.038 52.3 158.158 ;
      RECT 52.82 157.56 53.02 157.68 ;
      RECT 52.46 158.82 52.66 158.94 ;
      RECT 49.58 158.58 49.78 158.7 ;
      RECT 51.74 158.58 51.94 158.7 ;
      RECT 53.18 158.58 53.38 158.7 ;
      RECT 52.82 160.08 53.02 160.2 ;
      RECT 52.82 162.36 53.02 162.48 ;
      RECT 49.58 161.1 49.78 161.22 ;
      RECT 51.74 161.1 51.94 161.22 ;
      RECT 52.46 161.1 52.66 161.22 ;
      RECT 53.18 161.1 53.38 161.22 ;
      RECT 49.58 163.62 49.78 163.74 ;
      RECT 52.46 163.62 52.66 163.74 ;
      RECT 53.18 163.62 53.38 163.74 ;
      RECT 52.82 165.12 53.02 165.24 ;
      RECT 51.74 163.86 51.94 163.98 ;
      RECT 52.46 166.38 52.66 166.5 ;
      RECT 49.58 166.38 49.78 166.5 ;
      RECT 53.18 166.14 53.38 166.26 ;
      RECT 51.74 166.14 51.94 166.26 ;
      RECT 52.82 167.64 53.02 167.76 ;
      RECT 53.18 168.9 53.38 169.02 ;
      RECT 52.46 168.9 52.66 169.02 ;
      RECT 49.58 168.9 49.78 169.02 ;
      RECT 51.74 168.66 51.94 168.78 ;
      RECT 52.82 169.92 53.02 170.04 ;
      RECT 52.46 171.42 52.66 171.54 ;
      RECT 51.74 171.42 51.94 171.54 ;
      RECT 49.58 171.18 49.78 171.3 ;
      RECT 53.18 171.18 53.38 171.3 ;
      RECT 52.82 172.68 53.02 172.8 ;
      RECT 52.46 173.94 52.66 174.06 ;
      RECT 49.58 173.94 49.78 174.06 ;
      RECT 51.74 173.7 51.94 173.82 ;
      RECT 53.18 173.7 53.38 173.82 ;
      RECT 52.82 175.2 53.02 175.32 ;
      RECT 53.18 176.46 53.38 176.58 ;
      RECT 49.58 176.46 49.78 176.58 ;
      RECT 52.46 176.22 52.66 176.34 ;
      RECT 51.74 176.22 51.94 176.34 ;
      RECT 53.18 178.74 53.38 178.86 ;
      RECT 49.58 178.74 49.78 178.86 ;
      RECT 52.82 177.72 53.02 177.84 ;
      RECT 52.46 178.98 52.66 179.1 ;
      RECT 51.74 178.98 51.94 179.1 ;
      RECT 51.74 181.5 51.94 181.62 ;
      RECT 53.18 181.5 53.38 181.62 ;
      RECT 52.46 181.26 52.66 181.38 ;
      RECT 49.58 181.26 49.78 181.38 ;
      RECT 52.82 180.24 53.02 180.36 ;
      RECT 52.82 182.76 53.02 182.88 ;
      RECT 51.74 184.02 51.94 184.14 ;
      RECT 49.58 184.02 49.78 184.14 ;
      RECT 53.18 183.78 53.38 183.9 ;
      RECT 52.46 183.78 52.66 183.9 ;
      RECT 52.82 185.28 53.02 185.4 ;
      RECT 51.74 186.54 51.94 186.66 ;
      RECT 53.18 186.54 53.38 186.66 ;
      RECT 49.58 186.3 49.78 186.42 ;
      RECT 52.46 186.3 52.66 186.42 ;
      RECT 52.82 187.56 53.02 187.68 ;
      RECT 46.7 278.76 46.9 278.88 ;
      RECT 47.42 278.76 47.62 278.88 ;
      RECT 48.14 278.76 48.34 278.88 ;
      RECT 48.86 278.76 49.06 278.88 ;
      RECT 45.98 283.087 46.18 283.207 ;
      RECT 46.7 283.087 46.9 283.207 ;
      RECT 47.42 283.087 47.62 283.207 ;
      RECT 48.14 283.087 48.34 283.207 ;
      RECT 48.86 283.087 49.06 283.207 ;
      RECT 48.5 305.498 48.7 305.618 ;
      RECT 47.06 305.498 47.26 305.618 ;
      RECT 48.86 305.967 49.06 306.087 ;
      RECT 48.14 305.967 48.34 306.087 ;
      RECT 47.42 305.967 47.62 306.087 ;
      RECT 46.7 305.967 46.9 306.087 ;
      RECT 45.98 305.967 46.18 306.087 ;
      RECT 47.06 323.3835 47.26 323.5035 ;
      RECT 48.5 323.3835 48.7 323.5035 ;
      RECT 45.98 325.9425 46.18 326.0625 ;
      RECT 46.7 325.9425 46.9 326.0625 ;
      RECT 47.42 325.9425 47.62 326.0625 ;
      RECT 48.14 325.9425 48.34 326.0625 ;
      RECT 48.86 325.9425 49.06 326.0625 ;
      RECT 48.5 348.339 48.7 348.459 ;
      RECT 47.06 348.339 47.26 348.459 ;
      RECT 52.46 118.5 52.66 118.62 ;
      RECT 49.58 118.5 49.78 118.62 ;
      RECT 53.18 118.26 53.38 118.38 ;
      RECT 51.74 118.26 51.94 118.38 ;
      RECT 52.82 119.52 53.02 119.64 ;
      RECT 49.58 118.978 49.78 119.098 ;
      RECT 51.74 118.978 51.94 119.098 ;
      RECT 52.46 118.978 52.66 119.098 ;
      RECT 53.18 118.978 53.38 119.098 ;
      RECT 49.58 121.02 49.78 121.14 ;
      RECT 51.74 121.02 51.94 121.14 ;
      RECT 52.46 120.78 52.66 120.9 ;
      RECT 53.18 120.78 53.38 120.9 ;
      RECT 52.82 122.04 53.02 122.16 ;
      RECT 49.58 121.498 49.78 121.618 ;
      RECT 51.74 121.498 51.94 121.618 ;
      RECT 52.46 121.498 52.66 121.618 ;
      RECT 53.18 121.498 53.38 121.618 ;
      RECT 49.58 124.018 49.78 124.138 ;
      RECT 51.74 124.018 51.94 124.138 ;
      RECT 52.46 124.018 52.66 124.138 ;
      RECT 53.18 124.018 53.38 124.138 ;
      RECT 51.74 123.54 51.94 123.66 ;
      RECT 53.18 123.54 53.38 123.66 ;
      RECT 49.58 123.3 49.78 123.42 ;
      RECT 52.46 123.3 52.66 123.42 ;
      RECT 52.82 124.56 53.02 124.68 ;
      RECT 49.58 126.538 49.78 126.658 ;
      RECT 51.74 126.538 51.94 126.658 ;
      RECT 52.46 126.538 52.66 126.658 ;
      RECT 53.18 126.538 53.38 126.658 ;
      RECT 49.58 126.06 49.78 126.18 ;
      RECT 51.74 126.06 51.94 126.18 ;
      RECT 52.46 126.06 52.66 126.18 ;
      RECT 53.18 125.82 53.38 125.94 ;
      RECT 52.82 127.08 53.02 127.2 ;
      RECT 49.58 129.058 49.78 129.178 ;
      RECT 51.74 129.058 51.94 129.178 ;
      RECT 52.46 129.058 52.66 129.178 ;
      RECT 53.18 129.058 53.38 129.178 ;
      RECT 51.74 128.58 51.94 128.7 ;
      RECT 49.58 128.58 49.78 128.7 ;
      RECT 53.18 128.34 53.38 128.46 ;
      RECT 52.46 128.34 52.66 128.46 ;
      RECT 49.58 130.86 49.78 130.98 ;
      RECT 52.46 130.86 52.66 130.98 ;
      RECT 52.82 129.84 53.02 129.96 ;
      RECT 52.82 132.36 53.02 132.48 ;
      RECT 49.58 131.578 49.78 131.698 ;
      RECT 51.74 131.578 51.94 131.698 ;
      RECT 52.46 131.578 52.66 131.698 ;
      RECT 53.18 131.578 53.38 131.698 ;
      RECT 53.18 131.1 53.38 131.22 ;
      RECT 51.74 131.1 51.94 131.22 ;
      RECT 52.46 133.62 52.66 133.74 ;
      RECT 51.74 133.62 51.94 133.74 ;
      RECT 53.18 133.38 53.38 133.5 ;
      RECT 49.58 133.38 49.78 133.5 ;
      RECT 52.82 134.88 53.02 135 ;
      RECT 49.58 134.098 49.78 134.218 ;
      RECT 51.74 134.098 51.94 134.218 ;
      RECT 52.46 134.098 52.66 134.218 ;
      RECT 53.18 134.098 53.38 134.218 ;
      RECT 49.58 136.14 49.78 136.26 ;
      RECT 52.46 136.14 52.66 136.26 ;
      RECT 53.18 136.14 53.38 136.26 ;
      RECT 51.74 135.9 51.94 136.02 ;
      RECT 52.82 137.4 53.02 137.52 ;
      RECT 49.58 136.618 49.78 136.738 ;
      RECT 51.74 136.618 51.94 136.738 ;
      RECT 52.46 136.618 52.66 136.738 ;
      RECT 53.18 136.618 53.38 136.738 ;
      RECT 49.58 139.138 49.78 139.258 ;
      RECT 51.74 139.138 51.94 139.258 ;
      RECT 52.46 139.138 52.66 139.258 ;
      RECT 53.18 139.138 53.38 139.258 ;
      RECT 53.18 138.66 53.38 138.78 ;
      RECT 48.86 259.86 49.06 259.98 ;
      RECT 46.34 260.49 46.54 260.61 ;
      RECT 47.78 260.49 47.98 260.61 ;
      RECT 45.98 261.12 46.18 261.24 ;
      RECT 46.7 261.12 46.9 261.24 ;
      RECT 47.42 261.12 47.62 261.24 ;
      RECT 48.14 261.12 48.34 261.24 ;
      RECT 48.86 261.12 49.06 261.24 ;
      RECT 46.34 261.75 46.54 261.87 ;
      RECT 47.78 261.75 47.98 261.87 ;
      RECT 45.98 262.38 46.18 262.5 ;
      RECT 46.7 262.38 46.9 262.5 ;
      RECT 47.42 262.38 47.62 262.5 ;
      RECT 48.14 262.38 48.34 262.5 ;
      RECT 48.86 262.38 49.06 262.5 ;
      RECT 46.34 263.01 46.54 263.13 ;
      RECT 47.78 263.01 47.98 263.13 ;
      RECT 45.98 263.64 46.18 263.76 ;
      RECT 46.7 263.64 46.9 263.76 ;
      RECT 47.42 263.64 47.62 263.76 ;
      RECT 48.14 263.64 48.34 263.76 ;
      RECT 48.86 263.64 49.06 263.76 ;
      RECT 46.34 264.27 46.54 264.39 ;
      RECT 47.78 264.27 47.98 264.39 ;
      RECT 45.98 264.9 46.18 265.02 ;
      RECT 46.7 264.9 46.9 265.02 ;
      RECT 47.42 264.9 47.62 265.02 ;
      RECT 48.14 264.9 48.34 265.02 ;
      RECT 48.86 264.9 49.06 265.02 ;
      RECT 46.34 265.53 46.54 265.65 ;
      RECT 47.78 265.53 47.98 265.65 ;
      RECT 45.98 266.16 46.18 266.28 ;
      RECT 46.7 266.16 46.9 266.28 ;
      RECT 47.42 266.16 47.62 266.28 ;
      RECT 48.14 266.16 48.34 266.28 ;
      RECT 48.86 266.16 49.06 266.28 ;
      RECT 46.34 266.79 46.54 266.91 ;
      RECT 47.78 266.79 47.98 266.91 ;
      RECT 46.7 267.42 46.9 267.54 ;
      RECT 48.14 267.42 48.34 267.54 ;
      RECT 47.42 267.42 47.62 267.54 ;
      RECT 45.98 267.42 46.18 267.54 ;
      RECT 48.86 267.42 49.06 267.54 ;
      RECT 46.34 268.05 46.54 268.17 ;
      RECT 47.78 268.05 47.98 268.17 ;
      RECT 45.98 268.68 46.18 268.8 ;
      RECT 46.7 268.68 46.9 268.8 ;
      RECT 47.42 268.68 47.62 268.8 ;
      RECT 48.14 268.68 48.34 268.8 ;
      RECT 48.86 268.68 49.06 268.8 ;
      RECT 46.34 269.31 46.54 269.43 ;
      RECT 47.78 269.31 47.98 269.43 ;
      RECT 45.98 269.94 46.18 270.06 ;
      RECT 46.7 269.94 46.9 270.06 ;
      RECT 47.42 269.94 47.62 270.06 ;
      RECT 48.14 269.94 48.34 270.06 ;
      RECT 48.86 269.94 49.06 270.06 ;
      RECT 46.34 270.57 46.54 270.69 ;
      RECT 47.78 270.57 47.98 270.69 ;
      RECT 45.98 271.2 46.18 271.32 ;
      RECT 46.7 271.2 46.9 271.32 ;
      RECT 47.42 271.2 47.62 271.32 ;
      RECT 48.14 271.2 48.34 271.32 ;
      RECT 48.86 271.2 49.06 271.32 ;
      RECT 46.34 271.83 46.54 271.95 ;
      RECT 47.78 271.83 47.98 271.95 ;
      RECT 45.98 272.46 46.18 272.58 ;
      RECT 46.7 272.46 46.9 272.58 ;
      RECT 47.42 272.46 47.62 272.58 ;
      RECT 48.14 272.46 48.34 272.58 ;
      RECT 48.86 272.46 49.06 272.58 ;
      RECT 47.78 273.09 47.98 273.21 ;
      RECT 46.34 273.09 46.54 273.21 ;
      RECT 45.98 273.72 46.18 273.84 ;
      RECT 46.7 273.72 46.9 273.84 ;
      RECT 47.42 273.72 47.62 273.84 ;
      RECT 48.14 273.72 48.34 273.84 ;
      RECT 48.86 273.72 49.06 273.84 ;
      RECT 46.34 274.35 46.54 274.47 ;
      RECT 47.78 274.35 47.98 274.47 ;
      RECT 45.98 274.98 46.18 275.1 ;
      RECT 46.7 274.98 46.9 275.1 ;
      RECT 47.42 274.98 47.62 275.1 ;
      RECT 48.14 274.98 48.34 275.1 ;
      RECT 48.86 274.98 49.06 275.1 ;
      RECT 46.34 275.61 46.54 275.73 ;
      RECT 47.78 275.61 47.98 275.73 ;
      RECT 45.98 276.24 46.18 276.36 ;
      RECT 46.7 276.24 46.9 276.36 ;
      RECT 47.42 276.24 47.62 276.36 ;
      RECT 48.14 276.24 48.34 276.36 ;
      RECT 48.86 276.24 49.06 276.36 ;
      RECT 47.78 276.87 47.98 276.99 ;
      RECT 46.34 276.87 46.54 276.99 ;
      RECT 45.98 277.5 46.18 277.62 ;
      RECT 46.7 277.5 46.9 277.62 ;
      RECT 47.42 277.5 47.62 277.62 ;
      RECT 48.14 277.5 48.34 277.62 ;
      RECT 48.86 277.5 49.06 277.62 ;
      RECT 46.34 278.13 46.54 278.25 ;
      RECT 47.78 278.13 47.98 278.25 ;
      RECT 45.98 278.76 46.18 278.88 ;
      RECT 45.98 242.22 46.18 242.34 ;
      RECT 46.7 242.22 46.9 242.34 ;
      RECT 47.42 242.22 47.62 242.34 ;
      RECT 48.14 242.22 48.34 242.34 ;
      RECT 48.86 242.22 49.06 242.34 ;
      RECT 46.34 242.85 46.54 242.97 ;
      RECT 47.78 242.85 47.98 242.97 ;
      RECT 45.98 243.48 46.18 243.6 ;
      RECT 46.7 243.48 46.9 243.6 ;
      RECT 47.42 243.48 47.62 243.6 ;
      RECT 48.14 243.48 48.34 243.6 ;
      RECT 48.86 243.48 49.06 243.6 ;
      RECT 46.34 244.11 46.54 244.23 ;
      RECT 47.78 244.11 47.98 244.23 ;
      RECT 48.86 244.74 49.06 244.86 ;
      RECT 45.98 244.74 46.18 244.86 ;
      RECT 46.7 244.74 46.9 244.86 ;
      RECT 47.42 244.74 47.62 244.86 ;
      RECT 48.14 244.74 48.34 244.86 ;
      RECT 47.78 245.37 47.98 245.49 ;
      RECT 46.34 245.37 46.54 245.49 ;
      RECT 48.86 246 49.06 246.12 ;
      RECT 48.14 246 48.34 246.12 ;
      RECT 47.42 246 47.62 246.12 ;
      RECT 46.7 246 46.9 246.12 ;
      RECT 45.98 246 46.18 246.12 ;
      RECT 46.34 246.63 46.54 246.75 ;
      RECT 47.78 246.63 47.98 246.75 ;
      RECT 48.86 247.26 49.06 247.38 ;
      RECT 45.98 247.26 46.18 247.38 ;
      RECT 46.7 247.26 46.9 247.38 ;
      RECT 47.42 247.26 47.62 247.38 ;
      RECT 48.14 247.26 48.34 247.38 ;
      RECT 46.34 247.89 46.54 248.01 ;
      RECT 47.78 247.89 47.98 248.01 ;
      RECT 45.98 248.52 46.18 248.64 ;
      RECT 46.7 248.52 46.9 248.64 ;
      RECT 47.42 248.52 47.62 248.64 ;
      RECT 48.14 248.52 48.34 248.64 ;
      RECT 48.86 248.52 49.06 248.64 ;
      RECT 46.34 249.15 46.54 249.27 ;
      RECT 47.78 249.15 47.98 249.27 ;
      RECT 45.98 249.78 46.18 249.9 ;
      RECT 46.7 249.78 46.9 249.9 ;
      RECT 47.42 249.78 47.62 249.9 ;
      RECT 48.14 249.78 48.34 249.9 ;
      RECT 48.86 249.78 49.06 249.9 ;
      RECT 47.78 250.41 47.98 250.53 ;
      RECT 46.34 250.41 46.54 250.53 ;
      RECT 45.98 251.04 46.18 251.16 ;
      RECT 46.7 251.04 46.9 251.16 ;
      RECT 47.42 251.04 47.62 251.16 ;
      RECT 48.14 251.04 48.34 251.16 ;
      RECT 48.86 251.04 49.06 251.16 ;
      RECT 46.34 251.67 46.54 251.79 ;
      RECT 47.78 251.67 47.98 251.79 ;
      RECT 45.98 252.3 46.18 252.42 ;
      RECT 46.7 252.3 46.9 252.42 ;
      RECT 47.42 252.3 47.62 252.42 ;
      RECT 48.14 252.3 48.34 252.42 ;
      RECT 48.86 252.3 49.06 252.42 ;
      RECT 46.34 252.93 46.54 253.05 ;
      RECT 47.78 252.93 47.98 253.05 ;
      RECT 45.98 253.56 46.18 253.68 ;
      RECT 46.7 253.56 46.9 253.68 ;
      RECT 47.42 253.56 47.62 253.68 ;
      RECT 48.14 253.56 48.34 253.68 ;
      RECT 48.86 253.56 49.06 253.68 ;
      RECT 47.78 254.19 47.98 254.31 ;
      RECT 46.34 254.19 46.54 254.31 ;
      RECT 45.98 254.82 46.18 254.94 ;
      RECT 46.7 254.82 46.9 254.94 ;
      RECT 47.42 254.82 47.62 254.94 ;
      RECT 48.14 254.82 48.34 254.94 ;
      RECT 48.86 254.82 49.06 254.94 ;
      RECT 46.34 255.45 46.54 255.57 ;
      RECT 47.78 255.45 47.98 255.57 ;
      RECT 45.98 256.08 46.18 256.2 ;
      RECT 46.7 256.08 46.9 256.2 ;
      RECT 47.42 256.08 47.62 256.2 ;
      RECT 48.14 256.08 48.34 256.2 ;
      RECT 48.86 256.08 49.06 256.2 ;
      RECT 46.34 256.71 46.54 256.83 ;
      RECT 47.78 256.71 47.98 256.83 ;
      RECT 45.98 257.34 46.18 257.46 ;
      RECT 46.7 257.34 46.9 257.46 ;
      RECT 47.42 257.34 47.62 257.46 ;
      RECT 48.14 257.34 48.34 257.46 ;
      RECT 48.86 257.34 49.06 257.46 ;
      RECT 46.34 257.97 46.54 258.09 ;
      RECT 47.78 257.97 47.98 258.09 ;
      RECT 45.98 258.6 46.18 258.72 ;
      RECT 46.7 258.6 46.9 258.72 ;
      RECT 47.42 258.6 47.62 258.72 ;
      RECT 48.14 258.6 48.34 258.72 ;
      RECT 48.86 258.6 49.06 258.72 ;
      RECT 46.34 259.23 46.54 259.35 ;
      RECT 47.78 259.23 47.98 259.35 ;
      RECT 45.98 259.86 46.18 259.98 ;
      RECT 46.7 259.86 46.9 259.98 ;
      RECT 47.42 259.86 47.62 259.98 ;
      RECT 48.14 259.86 48.34 259.98 ;
      RECT 46.7 223.32 46.9 223.44 ;
      RECT 45.98 223.32 46.18 223.44 ;
      RECT 47.78 223.95 47.98 224.07 ;
      RECT 46.34 223.95 46.54 224.07 ;
      RECT 48.86 224.58 49.06 224.7 ;
      RECT 48.14 224.58 48.34 224.7 ;
      RECT 47.42 224.58 47.62 224.7 ;
      RECT 46.7 224.58 46.9 224.7 ;
      RECT 45.98 224.58 46.18 224.7 ;
      RECT 47.78 225.21 47.98 225.33 ;
      RECT 46.34 225.21 46.54 225.33 ;
      RECT 48.86 225.84 49.06 225.96 ;
      RECT 48.14 225.84 48.34 225.96 ;
      RECT 47.42 225.84 47.62 225.96 ;
      RECT 46.7 225.84 46.9 225.96 ;
      RECT 45.98 225.84 46.18 225.96 ;
      RECT 47.78 226.47 47.98 226.59 ;
      RECT 46.34 226.47 46.54 226.59 ;
      RECT 48.86 227.1 49.06 227.22 ;
      RECT 48.14 227.1 48.34 227.22 ;
      RECT 47.42 227.1 47.62 227.22 ;
      RECT 46.7 227.1 46.9 227.22 ;
      RECT 45.98 227.1 46.18 227.22 ;
      RECT 46.34 227.73 46.54 227.85 ;
      RECT 47.78 227.73 47.98 227.85 ;
      RECT 48.86 228.36 49.06 228.48 ;
      RECT 48.14 228.36 48.34 228.48 ;
      RECT 47.42 228.36 47.62 228.48 ;
      RECT 46.7 228.36 46.9 228.48 ;
      RECT 45.98 228.36 46.18 228.48 ;
      RECT 47.78 228.99 47.98 229.11 ;
      RECT 46.34 228.99 46.54 229.11 ;
      RECT 45.98 229.62 46.18 229.74 ;
      RECT 46.7 229.62 46.9 229.74 ;
      RECT 47.42 229.62 47.62 229.74 ;
      RECT 48.14 229.62 48.34 229.74 ;
      RECT 48.86 229.62 49.06 229.74 ;
      RECT 46.34 230.25 46.54 230.37 ;
      RECT 47.78 230.25 47.98 230.37 ;
      RECT 45.98 230.88 46.18 231 ;
      RECT 46.7 230.88 46.9 231 ;
      RECT 47.42 230.88 47.62 231 ;
      RECT 48.14 230.88 48.34 231 ;
      RECT 48.86 230.88 49.06 231 ;
      RECT 46.34 231.51 46.54 231.63 ;
      RECT 47.78 231.51 47.98 231.63 ;
      RECT 45.98 232.14 46.18 232.26 ;
      RECT 46.7 232.14 46.9 232.26 ;
      RECT 47.42 232.14 47.62 232.26 ;
      RECT 48.14 232.14 48.34 232.26 ;
      RECT 48.86 232.14 49.06 232.26 ;
      RECT 46.34 232.77 46.54 232.89 ;
      RECT 47.78 232.77 47.98 232.89 ;
      RECT 48.86 233.4 49.06 233.52 ;
      RECT 48.14 233.4 48.34 233.52 ;
      RECT 47.42 233.4 47.62 233.52 ;
      RECT 46.7 233.4 46.9 233.52 ;
      RECT 45.98 233.4 46.18 233.52 ;
      RECT 47.78 234.03 47.98 234.15 ;
      RECT 46.34 234.03 46.54 234.15 ;
      RECT 45.98 234.66 46.18 234.78 ;
      RECT 46.7 234.66 46.9 234.78 ;
      RECT 47.42 234.66 47.62 234.78 ;
      RECT 48.14 234.66 48.34 234.78 ;
      RECT 48.86 234.66 49.06 234.78 ;
      RECT 46.34 235.29 46.54 235.41 ;
      RECT 47.78 235.29 47.98 235.41 ;
      RECT 45.98 235.92 46.18 236.04 ;
      RECT 46.7 235.92 46.9 236.04 ;
      RECT 47.42 235.92 47.62 236.04 ;
      RECT 48.14 235.92 48.34 236.04 ;
      RECT 48.86 235.92 49.06 236.04 ;
      RECT 46.34 236.55 46.54 236.67 ;
      RECT 47.78 236.55 47.98 236.67 ;
      RECT 48.86 237.18 49.06 237.3 ;
      RECT 48.14 237.18 48.34 237.3 ;
      RECT 47.42 237.18 47.62 237.3 ;
      RECT 46.7 237.18 46.9 237.3 ;
      RECT 45.98 237.18 46.18 237.3 ;
      RECT 47.78 237.81 47.98 237.93 ;
      RECT 46.34 237.81 46.54 237.93 ;
      RECT 45.98 238.44 46.18 238.56 ;
      RECT 46.7 238.44 46.9 238.56 ;
      RECT 47.42 238.44 47.62 238.56 ;
      RECT 48.14 238.44 48.34 238.56 ;
      RECT 48.86 238.44 49.06 238.56 ;
      RECT 46.34 239.07 46.54 239.19 ;
      RECT 47.78 239.07 47.98 239.19 ;
      RECT 45.98 239.7 46.18 239.82 ;
      RECT 46.7 239.7 46.9 239.82 ;
      RECT 47.42 239.7 47.62 239.82 ;
      RECT 48.14 239.7 48.34 239.82 ;
      RECT 48.86 239.7 49.06 239.82 ;
      RECT 46.34 240.33 46.54 240.45 ;
      RECT 47.78 240.33 47.98 240.45 ;
      RECT 48.86 240.96 49.06 241.08 ;
      RECT 48.14 240.96 48.34 241.08 ;
      RECT 47.42 240.96 47.62 241.08 ;
      RECT 46.7 240.96 46.9 241.08 ;
      RECT 45.98 240.96 46.18 241.08 ;
      RECT 47.78 241.59 47.98 241.71 ;
      RECT 46.34 241.59 46.54 241.71 ;
      RECT 46.34 203.222 46.54 203.342 ;
      RECT 47.06 202.92 47.26 203.04 ;
      RECT 48.5 202.68 48.7 202.8 ;
      RECT 45.98 204.18 46.18 204.3 ;
      RECT 46.7 204.18 46.9 204.3 ;
      RECT 48.14 204.18 48.34 204.3 ;
      RECT 48.86 203.94 49.06 204.06 ;
      RECT 47.42 203.94 47.62 204.06 ;
      RECT 47.78 203.462 47.98 203.582 ;
      RECT 47.78 205.982 47.98 206.102 ;
      RECT 46.34 205.742 46.54 205.862 ;
      RECT 48.5 205.44 48.7 205.56 ;
      RECT 47.06 205.2 47.26 205.32 ;
      RECT 48.86 206.7 49.06 206.82 ;
      RECT 48.14 206.7 48.34 206.82 ;
      RECT 45.98 206.7 46.18 206.82 ;
      RECT 47.42 206.46 47.62 206.58 ;
      RECT 46.7 206.46 46.9 206.58 ;
      RECT 47.78 208.502 47.98 208.622 ;
      RECT 46.34 208.262 46.54 208.382 ;
      RECT 47.06 207.96 47.26 208.08 ;
      RECT 48.5 207.72 48.7 207.84 ;
      RECT 46.34 210.09 46.54 210.21 ;
      RECT 47.78 210.09 47.98 210.21 ;
      RECT 48.86 209.46 49.06 209.58 ;
      RECT 48.14 209.46 48.34 209.58 ;
      RECT 47.42 209.46 47.62 209.58 ;
      RECT 46.7 209.46 46.9 209.58 ;
      RECT 45.98 209.46 46.18 209.58 ;
      RECT 46.34 211.35 46.54 211.47 ;
      RECT 47.78 211.35 47.98 211.47 ;
      RECT 45.98 210.72 46.18 210.84 ;
      RECT 48.86 210.72 49.06 210.84 ;
      RECT 48.14 210.72 48.34 210.84 ;
      RECT 47.42 210.72 47.62 210.84 ;
      RECT 46.7 210.72 46.9 210.84 ;
      RECT 46.34 212.61 46.54 212.73 ;
      RECT 47.78 212.61 47.98 212.73 ;
      RECT 48.86 211.98 49.06 212.1 ;
      RECT 48.14 211.98 48.34 212.1 ;
      RECT 47.42 211.98 47.62 212.1 ;
      RECT 46.7 211.98 46.9 212.1 ;
      RECT 45.98 211.98 46.18 212.1 ;
      RECT 47.78 213.87 47.98 213.99 ;
      RECT 46.34 213.87 46.54 213.99 ;
      RECT 45.98 213.24 46.18 213.36 ;
      RECT 46.7 213.24 46.9 213.36 ;
      RECT 47.42 213.24 47.62 213.36 ;
      RECT 48.14 213.24 48.34 213.36 ;
      RECT 48.86 213.24 49.06 213.36 ;
      RECT 46.34 215.13 46.54 215.25 ;
      RECT 47.78 215.13 47.98 215.25 ;
      RECT 45.98 214.5 46.18 214.62 ;
      RECT 46.7 214.5 46.9 214.62 ;
      RECT 47.42 214.5 47.62 214.62 ;
      RECT 48.14 214.5 48.34 214.62 ;
      RECT 48.86 214.5 49.06 214.62 ;
      RECT 48.86 217.02 49.06 217.14 ;
      RECT 47.78 216.39 47.98 216.51 ;
      RECT 46.34 216.39 46.54 216.51 ;
      RECT 45.98 215.76 46.18 215.88 ;
      RECT 46.7 215.76 46.9 215.88 ;
      RECT 47.42 215.76 47.62 215.88 ;
      RECT 48.14 215.76 48.34 215.88 ;
      RECT 48.86 215.76 49.06 215.88 ;
      RECT 48.14 217.02 48.34 217.14 ;
      RECT 47.42 217.02 47.62 217.14 ;
      RECT 46.7 217.02 46.9 217.14 ;
      RECT 45.98 217.02 46.18 217.14 ;
      RECT 47.78 217.65 47.98 217.77 ;
      RECT 46.34 217.65 46.54 217.77 ;
      RECT 48.86 218.28 49.06 218.4 ;
      RECT 48.14 218.28 48.34 218.4 ;
      RECT 47.42 218.28 47.62 218.4 ;
      RECT 46.7 218.28 46.9 218.4 ;
      RECT 45.98 218.28 46.18 218.4 ;
      RECT 47.78 218.91 47.98 219.03 ;
      RECT 46.34 218.91 46.54 219.03 ;
      RECT 45.98 219.54 46.18 219.66 ;
      RECT 46.7 219.54 46.9 219.66 ;
      RECT 47.42 219.54 47.62 219.66 ;
      RECT 48.14 219.54 48.34 219.66 ;
      RECT 48.86 219.54 49.06 219.66 ;
      RECT 47.78 220.17 47.98 220.29 ;
      RECT 46.34 220.17 46.54 220.29 ;
      RECT 47.42 220.8 47.62 220.92 ;
      RECT 46.7 220.8 46.9 220.92 ;
      RECT 45.98 220.8 46.18 220.92 ;
      RECT 48.86 220.8 49.06 220.92 ;
      RECT 48.14 220.8 48.34 220.92 ;
      RECT 46.34 221.43 46.54 221.55 ;
      RECT 47.78 221.43 47.98 221.55 ;
      RECT 48.86 222.06 49.06 222.18 ;
      RECT 48.14 222.06 48.34 222.18 ;
      RECT 47.42 222.06 47.62 222.18 ;
      RECT 46.7 222.06 46.9 222.18 ;
      RECT 45.98 222.06 46.18 222.18 ;
      RECT 47.78 222.69 47.98 222.81 ;
      RECT 46.34 222.69 46.54 222.81 ;
      RECT 48.86 223.32 49.06 223.44 ;
      RECT 48.14 223.32 48.34 223.44 ;
      RECT 47.42 223.32 47.62 223.44 ;
      RECT 46.7 171.42 46.9 171.54 ;
      RECT 45.98 171.18 46.18 171.3 ;
      RECT 47.42 171.18 47.62 171.3 ;
      RECT 48.86 171.18 49.06 171.3 ;
      RECT 48.5 172.68 48.7 172.8 ;
      RECT 47.06 172.44 47.26 172.56 ;
      RECT 48.14 173.94 48.34 174.06 ;
      RECT 46.7 173.94 46.9 174.06 ;
      RECT 45.98 173.7 46.18 173.82 ;
      RECT 47.42 173.7 47.62 173.82 ;
      RECT 48.86 173.7 49.06 173.82 ;
      RECT 48.5 175.2 48.7 175.32 ;
      RECT 47.06 174.96 47.26 175.08 ;
      RECT 46.7 176.46 46.9 176.58 ;
      RECT 48.86 176.22 49.06 176.34 ;
      RECT 48.14 176.22 48.34 176.34 ;
      RECT 47.42 176.22 47.62 176.34 ;
      RECT 45.98 176.22 46.18 176.34 ;
      RECT 46.7 178.74 46.9 178.86 ;
      RECT 47.06 177.72 47.26 177.84 ;
      RECT 48.5 177.48 48.7 177.6 ;
      RECT 48.5 180 48.7 180.12 ;
      RECT 48.86 178.98 49.06 179.1 ;
      RECT 48.14 178.98 48.34 179.1 ;
      RECT 47.42 178.98 47.62 179.1 ;
      RECT 45.98 178.98 46.18 179.1 ;
      RECT 46.7 181.5 46.9 181.62 ;
      RECT 47.42 181.5 47.62 181.62 ;
      RECT 48.86 181.5 49.06 181.62 ;
      RECT 48.14 181.26 48.34 181.38 ;
      RECT 45.98 181.26 46.18 181.38 ;
      RECT 47.06 180.24 47.26 180.36 ;
      RECT 47.06 182.76 47.26 182.88 ;
      RECT 48.5 182.52 48.7 182.64 ;
      RECT 48.14 184.02 48.34 184.14 ;
      RECT 47.42 184.02 47.62 184.14 ;
      RECT 46.7 184.02 46.9 184.14 ;
      RECT 48.86 183.78 49.06 183.9 ;
      RECT 45.98 183.78 46.18 183.9 ;
      RECT 47.06 185.28 47.26 185.4 ;
      RECT 48.5 185.04 48.7 185.16 ;
      RECT 45.98 186.54 46.18 186.66 ;
      RECT 46.7 186.54 46.9 186.66 ;
      RECT 47.42 186.54 47.62 186.66 ;
      RECT 48.86 186.54 49.06 186.66 ;
      RECT 48.14 186.3 48.34 186.42 ;
      RECT 48.5 187.8 48.7 187.92 ;
      RECT 47.06 187.8 47.26 187.92 ;
      RECT 45.98 189.06 46.18 189.18 ;
      RECT 47.42 189.06 47.62 189.18 ;
      RECT 48.86 189.06 49.06 189.18 ;
      RECT 48.14 188.82 48.34 188.94 ;
      RECT 46.7 188.82 46.9 188.94 ;
      RECT 46.34 190.862 46.54 190.982 ;
      RECT 47.78 190.862 47.98 190.982 ;
      RECT 47.06 190.32 47.26 190.44 ;
      RECT 48.5 190.08 48.7 190.2 ;
      RECT 47.78 192.122 47.98 192.242 ;
      RECT 46.34 191.882 46.54 192.002 ;
      RECT 47.42 191.58 47.62 191.7 ;
      RECT 45.98 191.58 46.18 191.7 ;
      RECT 48.14 191.34 48.34 191.46 ;
      RECT 48.86 191.34 49.06 191.46 ;
      RECT 46.7 191.34 46.9 191.46 ;
      RECT 46.34 193.382 46.54 193.502 ;
      RECT 47.78 193.142 47.98 193.262 ;
      RECT 47.06 192.6 47.26 192.72 ;
      RECT 48.5 192.6 48.7 192.72 ;
      RECT 46.34 194.642 46.54 194.762 ;
      RECT 47.78 194.402 47.98 194.522 ;
      RECT 48.86 194.1 49.06 194.22 ;
      RECT 47.42 194.1 47.62 194.22 ;
      RECT 46.7 194.1 46.9 194.22 ;
      RECT 45.98 193.86 46.18 193.98 ;
      RECT 48.14 193.86 48.34 193.98 ;
      RECT 46.7 196.38 46.9 196.5 ;
      RECT 48.14 196.38 48.34 196.5 ;
      RECT 48.86 196.38 49.06 196.5 ;
      RECT 46.34 195.902 46.54 196.022 ;
      RECT 47.78 195.902 47.98 196.022 ;
      RECT 47.06 195.36 47.26 195.48 ;
      RECT 48.5 195.36 48.7 195.48 ;
      RECT 47.06 197.88 47.26 198 ;
      RECT 48.5 197.64 48.7 197.76 ;
      RECT 47.42 196.62 47.62 196.74 ;
      RECT 45.98 196.62 46.18 196.74 ;
      RECT 46.7 199.14 46.9 199.26 ;
      RECT 47.42 199.14 47.62 199.26 ;
      RECT 48.86 198.9 49.06 199.02 ;
      RECT 48.14 198.9 48.34 199.02 ;
      RECT 45.98 198.9 46.18 199.02 ;
      RECT 46.34 198.422 46.54 198.542 ;
      RECT 47.78 198.422 47.98 198.542 ;
      RECT 48.5 200.4 48.7 200.52 ;
      RECT 47.06 200.4 47.26 200.52 ;
      RECT 48.86 201.66 49.06 201.78 ;
      RECT 47.42 201.66 47.62 201.78 ;
      RECT 45.98 201.42 46.18 201.54 ;
      RECT 46.7 201.42 46.9 201.54 ;
      RECT 48.14 201.42 48.34 201.54 ;
      RECT 47.78 200.942 47.98 201.062 ;
      RECT 46.34 200.942 46.54 201.062 ;
      RECT 45.98 136.618 46.18 136.738 ;
      RECT 48.5 137.16 48.7 137.28 ;
      RECT 47.06 137.4 47.26 137.52 ;
      RECT 47.42 138.42 47.62 138.54 ;
      RECT 48.86 138.42 49.06 138.54 ;
      RECT 45.98 138.66 46.18 138.78 ;
      RECT 46.7 138.66 46.9 138.78 ;
      RECT 48.14 138.66 48.34 138.78 ;
      RECT 48.86 139.138 49.06 139.258 ;
      RECT 48.14 139.138 48.34 139.258 ;
      RECT 47.42 139.138 47.62 139.258 ;
      RECT 46.7 139.138 46.9 139.258 ;
      RECT 45.98 139.138 46.18 139.258 ;
      RECT 48.5 139.68 48.7 139.8 ;
      RECT 47.06 139.92 47.26 140.04 ;
      RECT 48.14 140.94 48.34 141.06 ;
      RECT 45.98 140.94 46.18 141.06 ;
      RECT 46.7 141.18 46.9 141.3 ;
      RECT 47.42 141.18 47.62 141.3 ;
      RECT 48.86 141.18 49.06 141.3 ;
      RECT 47.06 142.2 47.26 142.32 ;
      RECT 48.5 142.44 48.7 142.56 ;
      RECT 48.86 143.7 49.06 143.82 ;
      RECT 47.42 143.7 47.62 143.82 ;
      RECT 45.98 143.7 46.18 143.82 ;
      RECT 46.7 143.46 46.9 143.58 ;
      RECT 48.14 143.46 48.34 143.58 ;
      RECT 45.98 145.98 46.18 146.1 ;
      RECT 46.7 145.98 46.9 146.1 ;
      RECT 47.42 145.98 47.62 146.1 ;
      RECT 48.14 145.98 48.34 146.1 ;
      RECT 48.86 145.98 49.06 146.1 ;
      RECT 47.06 144.96 47.26 145.08 ;
      RECT 48.5 144.96 48.7 145.08 ;
      RECT 46.7 148.74 46.9 148.86 ;
      RECT 47.42 148.74 47.62 148.86 ;
      RECT 48.86 148.5 49.06 148.62 ;
      RECT 48.14 148.5 48.34 148.62 ;
      RECT 45.98 148.5 46.18 148.62 ;
      RECT 47.06 150 47.26 150.12 ;
      RECT 48.5 149.76 48.7 149.88 ;
      RECT 48.86 151.26 49.06 151.38 ;
      RECT 48.14 151.26 48.34 151.38 ;
      RECT 47.42 151.26 47.62 151.38 ;
      RECT 45.98 151.26 46.18 151.38 ;
      RECT 46.7 151.02 46.9 151.14 ;
      RECT 48.5 152.52 48.7 152.64 ;
      RECT 47.06 152.52 47.26 152.64 ;
      RECT 46.7 153.78 46.9 153.9 ;
      RECT 45.98 153.78 46.18 153.9 ;
      RECT 48.86 153.54 49.06 153.66 ;
      RECT 48.14 153.54 48.34 153.66 ;
      RECT 47.42 153.54 47.62 153.66 ;
      RECT 48.5 155.04 48.7 155.16 ;
      RECT 47.06 154.8 47.26 154.92 ;
      RECT 47.78 156.842 47.98 156.962 ;
      RECT 46.34 156.602 46.54 156.722 ;
      RECT 45.98 156.3 46.18 156.42 ;
      RECT 46.7 156.3 46.9 156.42 ;
      RECT 47.42 156.3 47.62 156.42 ;
      RECT 48.86 156.3 49.06 156.42 ;
      RECT 48.14 156.06 48.34 156.18 ;
      RECT 47.78 158.278 47.98 158.398 ;
      RECT 46.34 158.038 46.54 158.158 ;
      RECT 47.06 157.56 47.26 157.68 ;
      RECT 48.5 157.32 48.7 157.44 ;
      RECT 46.7 158.82 46.9 158.94 ;
      RECT 47.42 158.82 47.62 158.94 ;
      RECT 48.86 158.82 49.06 158.94 ;
      RECT 45.98 158.58 46.18 158.7 ;
      RECT 48.14 158.58 48.34 158.7 ;
      RECT 47.06 160.08 47.26 160.2 ;
      RECT 48.5 159.84 48.7 159.96 ;
      RECT 48.5 162.36 48.7 162.48 ;
      RECT 47.06 162.36 47.26 162.48 ;
      RECT 45.98 161.1 46.18 161.22 ;
      RECT 46.7 161.1 46.9 161.22 ;
      RECT 47.42 161.1 47.62 161.22 ;
      RECT 48.14 161.1 48.34 161.22 ;
      RECT 48.86 161.1 49.06 161.22 ;
      RECT 46.7 163.62 46.9 163.74 ;
      RECT 47.42 163.62 47.62 163.74 ;
      RECT 48.5 165.12 48.7 165.24 ;
      RECT 47.06 165.12 47.26 165.24 ;
      RECT 48.86 163.86 49.06 163.98 ;
      RECT 48.14 163.86 48.34 163.98 ;
      RECT 45.98 163.86 46.18 163.98 ;
      RECT 48.14 166.38 48.34 166.5 ;
      RECT 46.7 166.38 46.9 166.5 ;
      RECT 48.86 166.14 49.06 166.26 ;
      RECT 47.42 166.14 47.62 166.26 ;
      RECT 45.98 166.14 46.18 166.26 ;
      RECT 48.5 167.64 48.7 167.76 ;
      RECT 47.06 167.64 47.26 167.76 ;
      RECT 46.7 168.9 46.9 169.02 ;
      RECT 45.98 168.66 46.18 168.78 ;
      RECT 47.42 168.66 47.62 168.78 ;
      RECT 48.14 168.66 48.34 168.78 ;
      RECT 48.86 168.66 49.06 168.78 ;
      RECT 48.5 170.16 48.7 170.28 ;
      RECT 47.06 170.16 47.26 170.28 ;
      RECT 48.14 171.42 48.34 171.54 ;
      RECT 41.66 305.967 41.86 306.087 ;
      RECT 42.74 323.3835 42.94 323.5035 ;
      RECT 41.3 323.3835 41.5 323.5035 ;
      RECT 43.82 325.9425 44.02 326.0625 ;
      RECT 43.1 325.9425 43.3 326.0625 ;
      RECT 42.38 325.9425 42.58 326.0625 ;
      RECT 41.66 325.9425 41.86 326.0625 ;
      RECT 42.74 348.339 42.94 348.459 ;
      RECT 41.3 348.339 41.5 348.459 ;
      RECT 47.42 118.26 47.62 118.38 ;
      RECT 48.14 118.26 48.34 118.38 ;
      RECT 45.98 118.5 46.18 118.62 ;
      RECT 46.7 118.5 46.9 118.62 ;
      RECT 48.86 118.5 49.06 118.62 ;
      RECT 48.86 118.978 49.06 119.098 ;
      RECT 48.14 118.978 48.34 119.098 ;
      RECT 47.42 118.978 47.62 119.098 ;
      RECT 46.7 118.978 46.9 119.098 ;
      RECT 45.98 118.978 46.18 119.098 ;
      RECT 47.06 119.52 47.26 119.64 ;
      RECT 48.5 119.76 48.7 119.88 ;
      RECT 48.86 120.78 49.06 120.9 ;
      RECT 48.14 120.78 48.34 120.9 ;
      RECT 45.98 120.78 46.18 120.9 ;
      RECT 47.42 121.02 47.62 121.14 ;
      RECT 46.7 121.02 46.9 121.14 ;
      RECT 48.86 121.498 49.06 121.618 ;
      RECT 48.14 121.498 48.34 121.618 ;
      RECT 47.42 121.498 47.62 121.618 ;
      RECT 46.7 121.498 46.9 121.618 ;
      RECT 45.98 121.498 46.18 121.618 ;
      RECT 48.5 122.04 48.7 122.16 ;
      RECT 47.06 122.04 47.26 122.16 ;
      RECT 48.14 123.3 48.34 123.42 ;
      RECT 46.7 123.3 46.9 123.42 ;
      RECT 48.86 123.54 49.06 123.66 ;
      RECT 47.42 123.54 47.62 123.66 ;
      RECT 45.98 123.54 46.18 123.66 ;
      RECT 48.86 124.018 49.06 124.138 ;
      RECT 48.14 124.018 48.34 124.138 ;
      RECT 47.42 124.018 47.62 124.138 ;
      RECT 46.7 124.018 46.9 124.138 ;
      RECT 45.98 124.018 46.18 124.138 ;
      RECT 47.06 124.8 47.26 124.92 ;
      RECT 48.5 124.8 48.7 124.92 ;
      RECT 48.86 125.82 49.06 125.94 ;
      RECT 47.42 125.82 47.62 125.94 ;
      RECT 45.98 125.82 46.18 125.94 ;
      RECT 48.14 126.06 48.34 126.18 ;
      RECT 46.7 126.06 46.9 126.18 ;
      RECT 48.86 126.538 49.06 126.658 ;
      RECT 48.14 126.538 48.34 126.658 ;
      RECT 47.42 126.538 47.62 126.658 ;
      RECT 46.7 126.538 46.9 126.658 ;
      RECT 45.98 126.538 46.18 126.658 ;
      RECT 47.06 127.32 47.26 127.44 ;
      RECT 48.5 127.32 48.7 127.44 ;
      RECT 47.42 128.34 47.62 128.46 ;
      RECT 48.86 128.34 49.06 128.46 ;
      RECT 45.98 128.58 46.18 128.7 ;
      RECT 46.7 128.58 46.9 128.7 ;
      RECT 48.14 128.58 48.34 128.7 ;
      RECT 48.86 129.058 49.06 129.178 ;
      RECT 48.14 129.058 48.34 129.178 ;
      RECT 47.42 129.058 47.62 129.178 ;
      RECT 46.7 129.058 46.9 129.178 ;
      RECT 45.98 129.058 46.18 129.178 ;
      RECT 48.5 129.6 48.7 129.72 ;
      RECT 47.06 129.84 47.26 129.96 ;
      RECT 48.86 130.86 49.06 130.98 ;
      RECT 46.7 130.86 46.9 130.98 ;
      RECT 45.98 131.1 46.18 131.22 ;
      RECT 47.42 131.1 47.62 131.22 ;
      RECT 48.14 131.1 48.34 131.22 ;
      RECT 48.86 131.578 49.06 131.698 ;
      RECT 48.14 131.578 48.34 131.698 ;
      RECT 47.42 131.578 47.62 131.698 ;
      RECT 46.7 131.578 46.9 131.698 ;
      RECT 45.98 131.578 46.18 131.698 ;
      RECT 47.06 132.12 47.26 132.24 ;
      RECT 48.5 132.12 48.7 132.24 ;
      RECT 48.14 133.38 48.34 133.5 ;
      RECT 48.86 133.62 49.06 133.74 ;
      RECT 47.42 133.62 47.62 133.74 ;
      RECT 46.7 133.62 46.9 133.74 ;
      RECT 45.98 133.62 46.18 133.74 ;
      RECT 48.86 134.098 49.06 134.218 ;
      RECT 48.14 134.098 48.34 134.218 ;
      RECT 47.42 134.098 47.62 134.218 ;
      RECT 46.7 134.098 46.9 134.218 ;
      RECT 45.98 134.098 46.18 134.218 ;
      RECT 47.06 134.64 47.26 134.76 ;
      RECT 48.5 134.88 48.7 135 ;
      RECT 45.98 135.9 46.18 136.02 ;
      RECT 47.42 135.9 47.62 136.02 ;
      RECT 48.86 135.9 49.06 136.02 ;
      RECT 48.14 136.14 48.34 136.26 ;
      RECT 46.7 136.14 46.9 136.26 ;
      RECT 48.86 136.618 49.06 136.738 ;
      RECT 48.14 136.618 48.34 136.738 ;
      RECT 47.42 136.618 47.62 136.738 ;
      RECT 46.7 136.618 46.9 136.738 ;
      RECT 42.02 260.49 42.22 260.61 ;
      RECT 43.82 259.86 44.02 259.98 ;
      RECT 43.1 259.86 43.3 259.98 ;
      RECT 42.38 259.86 42.58 259.98 ;
      RECT 41.66 259.86 41.86 259.98 ;
      RECT 43.46 261.75 43.66 261.87 ;
      RECT 42.02 261.75 42.22 261.87 ;
      RECT 42.38 261.12 42.58 261.24 ;
      RECT 41.66 261.12 41.86 261.24 ;
      RECT 43.82 261.12 44.02 261.24 ;
      RECT 43.1 261.12 43.3 261.24 ;
      RECT 43.46 263.01 43.66 263.13 ;
      RECT 42.02 263.01 42.22 263.13 ;
      RECT 43.82 262.38 44.02 262.5 ;
      RECT 43.1 262.38 43.3 262.5 ;
      RECT 42.38 262.38 42.58 262.5 ;
      RECT 41.66 262.38 41.86 262.5 ;
      RECT 43.46 264.27 43.66 264.39 ;
      RECT 42.02 264.27 42.22 264.39 ;
      RECT 43.82 263.64 44.02 263.76 ;
      RECT 43.1 263.64 43.3 263.76 ;
      RECT 42.38 263.64 42.58 263.76 ;
      RECT 41.66 263.64 41.86 263.76 ;
      RECT 43.82 266.16 44.02 266.28 ;
      RECT 43.1 266.16 43.3 266.28 ;
      RECT 42.38 266.16 42.58 266.28 ;
      RECT 41.66 266.16 41.86 266.28 ;
      RECT 43.46 265.53 43.66 265.65 ;
      RECT 42.02 265.53 42.22 265.65 ;
      RECT 43.82 264.9 44.02 265.02 ;
      RECT 43.1 264.9 43.3 265.02 ;
      RECT 42.38 264.9 42.58 265.02 ;
      RECT 41.66 264.9 41.86 265.02 ;
      RECT 43.82 267.42 44.02 267.54 ;
      RECT 43.1 267.42 43.3 267.54 ;
      RECT 42.38 267.42 42.58 267.54 ;
      RECT 41.66 267.42 41.86 267.54 ;
      RECT 43.46 266.79 43.66 266.91 ;
      RECT 42.02 266.79 42.22 266.91 ;
      RECT 43.82 268.68 44.02 268.8 ;
      RECT 43.1 268.68 43.3 268.8 ;
      RECT 42.38 268.68 42.58 268.8 ;
      RECT 41.66 268.68 41.86 268.8 ;
      RECT 43.46 268.05 43.66 268.17 ;
      RECT 42.02 268.05 42.22 268.17 ;
      RECT 43.82 269.94 44.02 270.06 ;
      RECT 43.1 269.94 43.3 270.06 ;
      RECT 42.38 269.94 42.58 270.06 ;
      RECT 41.66 269.94 41.86 270.06 ;
      RECT 43.46 269.31 43.66 269.43 ;
      RECT 42.02 269.31 42.22 269.43 ;
      RECT 43.82 271.2 44.02 271.32 ;
      RECT 43.1 271.2 43.3 271.32 ;
      RECT 42.38 271.2 42.58 271.32 ;
      RECT 41.66 271.2 41.86 271.32 ;
      RECT 43.46 270.57 43.66 270.69 ;
      RECT 42.02 270.57 42.22 270.69 ;
      RECT 42.02 271.83 42.22 271.95 ;
      RECT 43.46 271.83 43.66 271.95 ;
      RECT 41.66 272.46 41.86 272.58 ;
      RECT 42.38 272.46 42.58 272.58 ;
      RECT 43.1 272.46 43.3 272.58 ;
      RECT 43.82 272.46 44.02 272.58 ;
      RECT 43.46 273.09 43.66 273.21 ;
      RECT 42.02 273.09 42.22 273.21 ;
      RECT 41.66 273.72 41.86 273.84 ;
      RECT 42.38 273.72 42.58 273.84 ;
      RECT 43.1 273.72 43.3 273.84 ;
      RECT 43.82 273.72 44.02 273.84 ;
      RECT 42.02 274.35 42.22 274.47 ;
      RECT 43.46 274.35 43.66 274.47 ;
      RECT 43.1 274.98 43.3 275.1 ;
      RECT 43.82 274.98 44.02 275.1 ;
      RECT 41.66 274.98 41.86 275.1 ;
      RECT 42.38 274.98 42.58 275.1 ;
      RECT 42.02 275.61 42.22 275.73 ;
      RECT 43.46 275.61 43.66 275.73 ;
      RECT 41.66 276.24 41.86 276.36 ;
      RECT 42.38 276.24 42.58 276.36 ;
      RECT 43.1 276.24 43.3 276.36 ;
      RECT 43.82 276.24 44.02 276.36 ;
      RECT 42.02 276.87 42.22 276.99 ;
      RECT 43.46 276.87 43.66 276.99 ;
      RECT 41.66 277.5 41.86 277.62 ;
      RECT 42.38 277.5 42.58 277.62 ;
      RECT 43.1 277.5 43.3 277.62 ;
      RECT 43.82 277.5 44.02 277.62 ;
      RECT 42.02 278.13 42.22 278.25 ;
      RECT 43.46 278.13 43.66 278.25 ;
      RECT 41.66 278.76 41.86 278.88 ;
      RECT 42.38 278.76 42.58 278.88 ;
      RECT 43.1 278.76 43.3 278.88 ;
      RECT 43.82 278.76 44.02 278.88 ;
      RECT 41.66 283.087 41.86 283.207 ;
      RECT 42.38 283.087 42.58 283.207 ;
      RECT 43.1 283.087 43.3 283.207 ;
      RECT 43.82 283.087 44.02 283.207 ;
      RECT 42.74 305.498 42.94 305.618 ;
      RECT 41.3 305.498 41.5 305.618 ;
      RECT 43.82 305.967 44.02 306.087 ;
      RECT 43.1 305.967 43.3 306.087 ;
      RECT 42.38 305.967 42.58 306.087 ;
      RECT 41.66 238.44 41.86 238.56 ;
      RECT 42.02 237.81 42.22 237.93 ;
      RECT 43.46 237.81 43.66 237.93 ;
      RECT 43.82 239.7 44.02 239.82 ;
      RECT 43.1 239.7 43.3 239.82 ;
      RECT 42.38 239.7 42.58 239.82 ;
      RECT 41.66 239.7 41.86 239.82 ;
      RECT 43.46 239.07 43.66 239.19 ;
      RECT 42.02 239.07 42.22 239.19 ;
      RECT 42.02 241.59 42.22 241.71 ;
      RECT 43.46 241.59 43.66 241.71 ;
      RECT 41.66 240.96 41.86 241.08 ;
      RECT 42.38 240.96 42.58 241.08 ;
      RECT 43.1 240.96 43.3 241.08 ;
      RECT 43.82 240.96 44.02 241.08 ;
      RECT 42.02 240.33 42.22 240.45 ;
      RECT 43.46 240.33 43.66 240.45 ;
      RECT 43.46 242.85 43.66 242.97 ;
      RECT 42.02 242.85 42.22 242.97 ;
      RECT 43.82 242.22 44.02 242.34 ;
      RECT 43.1 242.22 43.3 242.34 ;
      RECT 42.38 242.22 42.58 242.34 ;
      RECT 41.66 242.22 41.86 242.34 ;
      RECT 43.46 244.11 43.66 244.23 ;
      RECT 42.02 244.11 42.22 244.23 ;
      RECT 43.82 243.48 44.02 243.6 ;
      RECT 43.1 243.48 43.3 243.6 ;
      RECT 42.38 243.48 42.58 243.6 ;
      RECT 41.66 243.48 41.86 243.6 ;
      RECT 42.02 245.37 42.22 245.49 ;
      RECT 43.46 245.37 43.66 245.49 ;
      RECT 41.66 244.74 41.86 244.86 ;
      RECT 42.38 244.74 42.58 244.86 ;
      RECT 43.1 244.74 43.3 244.86 ;
      RECT 43.82 244.74 44.02 244.86 ;
      RECT 41.66 246 41.86 246.12 ;
      RECT 42.38 246 42.58 246.12 ;
      RECT 43.1 246 43.3 246.12 ;
      RECT 43.82 246 44.02 246.12 ;
      RECT 42.02 246.63 42.22 246.75 ;
      RECT 43.46 246.63 43.66 246.75 ;
      RECT 41.66 247.26 41.86 247.38 ;
      RECT 42.38 247.26 42.58 247.38 ;
      RECT 43.1 247.26 43.3 247.38 ;
      RECT 43.82 247.26 44.02 247.38 ;
      RECT 42.02 247.89 42.22 248.01 ;
      RECT 43.46 247.89 43.66 248.01 ;
      RECT 43.82 249.78 44.02 249.9 ;
      RECT 43.1 249.78 43.3 249.9 ;
      RECT 42.38 249.78 42.58 249.9 ;
      RECT 41.66 249.78 41.86 249.9 ;
      RECT 43.46 249.15 43.66 249.27 ;
      RECT 42.02 249.15 42.22 249.27 ;
      RECT 42.38 248.52 42.58 248.64 ;
      RECT 41.66 248.52 41.86 248.64 ;
      RECT 43.82 248.52 44.02 248.64 ;
      RECT 43.1 248.52 43.3 248.64 ;
      RECT 43.82 251.04 44.02 251.16 ;
      RECT 43.1 251.04 43.3 251.16 ;
      RECT 42.38 251.04 42.58 251.16 ;
      RECT 41.66 251.04 41.86 251.16 ;
      RECT 42.02 250.41 42.22 250.53 ;
      RECT 43.46 250.41 43.66 250.53 ;
      RECT 43.82 252.3 44.02 252.42 ;
      RECT 43.1 252.3 43.3 252.42 ;
      RECT 42.38 252.3 42.58 252.42 ;
      RECT 41.66 252.3 41.86 252.42 ;
      RECT 43.46 251.67 43.66 251.79 ;
      RECT 42.02 251.67 42.22 251.79 ;
      RECT 43.82 253.56 44.02 253.68 ;
      RECT 43.1 253.56 43.3 253.68 ;
      RECT 42.38 253.56 42.58 253.68 ;
      RECT 41.66 253.56 41.86 253.68 ;
      RECT 43.46 252.93 43.66 253.05 ;
      RECT 42.02 252.93 42.22 253.05 ;
      RECT 43.82 254.82 44.02 254.94 ;
      RECT 43.1 254.82 43.3 254.94 ;
      RECT 42.38 254.82 42.58 254.94 ;
      RECT 41.66 254.82 41.86 254.94 ;
      RECT 42.02 254.19 42.22 254.31 ;
      RECT 43.46 254.19 43.66 254.31 ;
      RECT 43.82 256.08 44.02 256.2 ;
      RECT 43.1 256.08 43.3 256.2 ;
      RECT 42.38 256.08 42.58 256.2 ;
      RECT 41.66 256.08 41.86 256.2 ;
      RECT 43.46 255.45 43.66 255.57 ;
      RECT 42.02 255.45 42.22 255.57 ;
      RECT 43.46 257.97 43.66 258.09 ;
      RECT 42.02 257.97 42.22 258.09 ;
      RECT 43.82 257.34 44.02 257.46 ;
      RECT 43.1 257.34 43.3 257.46 ;
      RECT 42.38 257.34 42.58 257.46 ;
      RECT 41.66 257.34 41.86 257.46 ;
      RECT 43.46 256.71 43.66 256.83 ;
      RECT 42.02 256.71 42.22 256.83 ;
      RECT 43.46 259.23 43.66 259.35 ;
      RECT 42.02 259.23 42.22 259.35 ;
      RECT 43.82 258.6 44.02 258.72 ;
      RECT 43.1 258.6 43.3 258.72 ;
      RECT 42.38 258.6 42.58 258.72 ;
      RECT 41.66 258.6 41.86 258.72 ;
      RECT 43.46 260.49 43.66 260.61 ;
      RECT 43.82 215.76 44.02 215.88 ;
      RECT 41.66 215.76 41.86 215.88 ;
      RECT 42.38 215.76 42.58 215.88 ;
      RECT 41.66 218.28 41.86 218.4 ;
      RECT 42.38 218.28 42.58 218.4 ;
      RECT 43.1 218.28 43.3 218.4 ;
      RECT 43.82 218.28 44.02 218.4 ;
      RECT 42.02 217.65 42.22 217.77 ;
      RECT 43.46 217.65 43.66 217.77 ;
      RECT 43.82 219.54 44.02 219.66 ;
      RECT 43.1 219.54 43.3 219.66 ;
      RECT 42.38 219.54 42.58 219.66 ;
      RECT 41.66 219.54 41.86 219.66 ;
      RECT 42.02 218.91 42.22 219.03 ;
      RECT 43.46 218.91 43.66 219.03 ;
      RECT 42.02 220.17 42.22 220.29 ;
      RECT 43.46 220.17 43.66 220.29 ;
      RECT 41.66 220.8 41.86 220.92 ;
      RECT 42.38 220.8 42.58 220.92 ;
      RECT 43.1 220.8 43.3 220.92 ;
      RECT 43.82 220.8 44.02 220.92 ;
      RECT 41.66 222.06 41.86 222.18 ;
      RECT 42.38 222.06 42.58 222.18 ;
      RECT 43.1 222.06 43.3 222.18 ;
      RECT 43.82 222.06 44.02 222.18 ;
      RECT 42.02 221.43 42.22 221.55 ;
      RECT 43.46 221.43 43.66 221.55 ;
      RECT 41.66 223.32 41.86 223.44 ;
      RECT 42.38 223.32 42.58 223.44 ;
      RECT 43.1 223.32 43.3 223.44 ;
      RECT 43.82 223.32 44.02 223.44 ;
      RECT 42.02 222.69 42.22 222.81 ;
      RECT 43.46 222.69 43.66 222.81 ;
      RECT 42.02 225.21 42.22 225.33 ;
      RECT 43.46 225.21 43.66 225.33 ;
      RECT 41.66 224.58 41.86 224.7 ;
      RECT 42.38 224.58 42.58 224.7 ;
      RECT 43.1 224.58 43.3 224.7 ;
      RECT 43.82 224.58 44.02 224.7 ;
      RECT 42.02 223.95 42.22 224.07 ;
      RECT 43.46 223.95 43.66 224.07 ;
      RECT 42.02 226.47 42.22 226.59 ;
      RECT 43.46 226.47 43.66 226.59 ;
      RECT 41.66 225.84 41.86 225.96 ;
      RECT 42.38 225.84 42.58 225.96 ;
      RECT 43.1 225.84 43.3 225.96 ;
      RECT 43.82 225.84 44.02 225.96 ;
      RECT 43.46 227.73 43.66 227.85 ;
      RECT 42.02 227.73 42.22 227.85 ;
      RECT 41.66 227.1 41.86 227.22 ;
      RECT 42.38 227.1 42.58 227.22 ;
      RECT 43.1 227.1 43.3 227.22 ;
      RECT 43.82 227.1 44.02 227.22 ;
      RECT 42.02 228.99 42.22 229.11 ;
      RECT 43.46 228.99 43.66 229.11 ;
      RECT 43.82 228.36 44.02 228.48 ;
      RECT 41.66 228.36 41.86 228.48 ;
      RECT 42.38 228.36 42.58 228.48 ;
      RECT 43.1 228.36 43.3 228.48 ;
      RECT 43.46 230.25 43.66 230.37 ;
      RECT 42.02 230.25 42.22 230.37 ;
      RECT 41.66 229.62 41.86 229.74 ;
      RECT 42.38 229.62 42.58 229.74 ;
      RECT 43.82 229.62 44.02 229.74 ;
      RECT 43.1 229.62 43.3 229.74 ;
      RECT 43.46 231.51 43.66 231.63 ;
      RECT 42.02 231.51 42.22 231.63 ;
      RECT 43.82 230.88 44.02 231 ;
      RECT 43.1 230.88 43.3 231 ;
      RECT 42.38 230.88 42.58 231 ;
      RECT 41.66 230.88 41.86 231 ;
      RECT 43.1 233.4 43.3 233.52 ;
      RECT 43.82 233.4 44.02 233.52 ;
      RECT 41.66 233.4 41.86 233.52 ;
      RECT 42.38 233.4 42.58 233.52 ;
      RECT 43.46 232.77 43.66 232.89 ;
      RECT 42.02 232.77 42.22 232.89 ;
      RECT 43.82 232.14 44.02 232.26 ;
      RECT 43.1 232.14 43.3 232.26 ;
      RECT 42.38 232.14 42.58 232.26 ;
      RECT 41.66 232.14 41.86 232.26 ;
      RECT 43.82 234.66 44.02 234.78 ;
      RECT 43.1 234.66 43.3 234.78 ;
      RECT 42.38 234.66 42.58 234.78 ;
      RECT 41.66 234.66 41.86 234.78 ;
      RECT 42.02 234.03 42.22 234.15 ;
      RECT 43.46 234.03 43.66 234.15 ;
      RECT 43.82 235.92 44.02 236.04 ;
      RECT 43.1 235.92 43.3 236.04 ;
      RECT 42.38 235.92 42.58 236.04 ;
      RECT 41.66 235.92 41.86 236.04 ;
      RECT 43.46 235.29 43.66 235.41 ;
      RECT 42.02 235.29 42.22 235.41 ;
      RECT 41.66 237.18 41.86 237.3 ;
      RECT 42.38 237.18 42.58 237.3 ;
      RECT 43.1 237.18 43.3 237.3 ;
      RECT 43.82 237.18 44.02 237.3 ;
      RECT 43.46 236.55 43.66 236.67 ;
      RECT 42.02 236.55 42.22 236.67 ;
      RECT 43.82 238.44 44.02 238.56 ;
      RECT 43.1 238.44 43.3 238.56 ;
      RECT 42.38 238.44 42.58 238.56 ;
      RECT 41.66 188.82 41.86 188.94 ;
      RECT 42.02 190.862 42.22 190.982 ;
      RECT 43.46 190.622 43.66 190.742 ;
      RECT 42.74 190.32 42.94 190.44 ;
      RECT 41.3 190.32 41.5 190.44 ;
      RECT 43.46 192.122 43.66 192.242 ;
      RECT 42.02 191.882 42.22 192.002 ;
      RECT 43.1 191.58 43.3 191.7 ;
      RECT 41.66 191.58 41.86 191.7 ;
      RECT 42.38 191.34 42.58 191.46 ;
      RECT 43.82 191.34 44.02 191.46 ;
      RECT 42.02 193.382 42.22 193.502 ;
      RECT 43.46 193.142 43.66 193.262 ;
      RECT 42.74 192.84 42.94 192.96 ;
      RECT 41.3 192.84 41.5 192.96 ;
      RECT 42.74 195.12 42.94 195.24 ;
      RECT 42.02 194.642 42.22 194.762 ;
      RECT 43.46 194.402 43.66 194.522 ;
      RECT 43.1 194.1 43.3 194.22 ;
      RECT 42.38 194.1 42.58 194.22 ;
      RECT 41.66 193.86 41.86 193.98 ;
      RECT 43.82 193.86 44.02 193.98 ;
      RECT 41.66 196.38 41.86 196.5 ;
      RECT 43.82 196.38 44.02 196.5 ;
      RECT 43.46 195.902 43.66 196.022 ;
      RECT 42.02 195.662 42.22 195.782 ;
      RECT 41.3 195.36 41.5 195.48 ;
      RECT 41.3 197.88 41.5 198 ;
      RECT 42.74 197.64 42.94 197.76 ;
      RECT 43.1 196.62 43.3 196.74 ;
      RECT 42.38 196.62 42.58 196.74 ;
      RECT 41.66 199.14 41.86 199.26 ;
      RECT 42.38 199.14 42.58 199.26 ;
      RECT 43.82 198.9 44.02 199.02 ;
      RECT 43.1 198.9 43.3 199.02 ;
      RECT 42.02 198.422 42.22 198.542 ;
      RECT 43.46 198.182 43.66 198.302 ;
      RECT 42.74 200.4 42.94 200.52 ;
      RECT 41.3 200.4 41.5 200.52 ;
      RECT 43.82 201.66 44.02 201.78 ;
      RECT 42.38 201.66 42.58 201.78 ;
      RECT 41.66 201.42 41.86 201.54 ;
      RECT 43.1 201.42 43.3 201.54 ;
      RECT 43.46 200.942 43.66 201.062 ;
      RECT 42.02 200.702 42.22 200.822 ;
      RECT 42.02 203.222 42.22 203.342 ;
      RECT 41.3 202.92 41.5 203.04 ;
      RECT 42.74 202.68 42.94 202.8 ;
      RECT 41.66 204.18 41.86 204.3 ;
      RECT 42.38 204.18 42.58 204.3 ;
      RECT 43.82 203.94 44.02 204.06 ;
      RECT 43.1 203.94 43.3 204.06 ;
      RECT 43.46 203.462 43.66 203.582 ;
      RECT 43.46 205.982 43.66 206.102 ;
      RECT 42.02 205.742 42.22 205.862 ;
      RECT 41.3 205.44 41.5 205.56 ;
      RECT 42.74 205.2 42.94 205.32 ;
      RECT 43.82 206.7 44.02 206.82 ;
      RECT 42.38 206.7 42.58 206.82 ;
      RECT 43.1 206.46 43.3 206.58 ;
      RECT 41.66 206.46 41.86 206.58 ;
      RECT 43.46 208.502 43.66 208.622 ;
      RECT 42.02 208.262 42.22 208.382 ;
      RECT 42.74 207.96 42.94 208.08 ;
      RECT 41.3 207.72 41.5 207.84 ;
      RECT 42.02 210.09 42.22 210.21 ;
      RECT 43.46 210.09 43.66 210.21 ;
      RECT 43.82 209.46 44.02 209.58 ;
      RECT 43.1 209.46 43.3 209.58 ;
      RECT 42.38 209.46 42.58 209.58 ;
      RECT 41.66 209.46 41.86 209.58 ;
      RECT 42.02 211.35 42.22 211.47 ;
      RECT 43.46 211.35 43.66 211.47 ;
      RECT 41.66 210.72 41.86 210.84 ;
      RECT 42.38 210.72 42.58 210.84 ;
      RECT 43.1 210.72 43.3 210.84 ;
      RECT 43.82 210.72 44.02 210.84 ;
      RECT 42.02 212.61 42.22 212.73 ;
      RECT 43.46 212.61 43.66 212.73 ;
      RECT 43.82 211.98 44.02 212.1 ;
      RECT 43.1 211.98 43.3 212.1 ;
      RECT 42.38 211.98 42.58 212.1 ;
      RECT 41.66 211.98 41.86 212.1 ;
      RECT 42.02 213.87 42.22 213.99 ;
      RECT 43.46 213.87 43.66 213.99 ;
      RECT 41.66 213.24 41.86 213.36 ;
      RECT 42.38 213.24 42.58 213.36 ;
      RECT 43.1 213.24 43.3 213.36 ;
      RECT 43.82 213.24 44.02 213.36 ;
      RECT 42.02 215.13 42.22 215.25 ;
      RECT 43.46 215.13 43.66 215.25 ;
      RECT 41.66 214.5 41.86 214.62 ;
      RECT 42.38 214.5 42.58 214.62 ;
      RECT 43.1 214.5 43.3 214.62 ;
      RECT 43.82 214.5 44.02 214.62 ;
      RECT 41.66 217.02 41.86 217.14 ;
      RECT 42.38 217.02 42.58 217.14 ;
      RECT 43.1 217.02 43.3 217.14 ;
      RECT 43.82 217.02 44.02 217.14 ;
      RECT 43.46 216.39 43.66 216.51 ;
      RECT 42.02 216.39 42.22 216.51 ;
      RECT 43.1 215.76 43.3 215.88 ;
      RECT 42.38 148.74 42.58 148.86 ;
      RECT 43.82 148.5 44.02 148.62 ;
      RECT 43.1 148.5 43.3 148.62 ;
      RECT 42.74 150 42.94 150.12 ;
      RECT 41.3 150 41.5 150.12 ;
      RECT 43.1 151.26 43.3 151.38 ;
      RECT 43.82 151.02 44.02 151.14 ;
      RECT 42.38 151.02 42.58 151.14 ;
      RECT 41.66 151.02 41.86 151.14 ;
      RECT 41.3 152.52 41.5 152.64 ;
      RECT 42.74 152.52 42.94 152.64 ;
      RECT 43.82 153.78 44.02 153.9 ;
      RECT 42.38 153.78 42.58 153.9 ;
      RECT 43.1 153.54 43.3 153.66 ;
      RECT 41.66 153.54 41.86 153.66 ;
      RECT 42.74 155.04 42.94 155.16 ;
      RECT 41.3 154.8 41.5 154.92 ;
      RECT 43.46 156.842 43.66 156.962 ;
      RECT 42.02 156.602 42.22 156.722 ;
      RECT 43.1 156.3 43.3 156.42 ;
      RECT 42.38 156.3 42.58 156.42 ;
      RECT 43.82 156.06 44.02 156.18 ;
      RECT 41.66 156.06 41.86 156.18 ;
      RECT 43.46 158.278 43.66 158.398 ;
      RECT 42.02 158.038 42.22 158.158 ;
      RECT 41.3 157.56 41.5 157.68 ;
      RECT 42.74 157.32 42.94 157.44 ;
      RECT 42.38 158.82 42.58 158.94 ;
      RECT 41.66 158.82 41.86 158.94 ;
      RECT 43.82 158.82 44.02 158.94 ;
      RECT 43.1 158.58 43.3 158.7 ;
      RECT 41.3 160.08 41.5 160.2 ;
      RECT 42.74 159.84 42.94 159.96 ;
      RECT 41.66 161.1 41.86 161.22 ;
      RECT 42.38 161.1 42.58 161.22 ;
      RECT 43.1 161.1 43.3 161.22 ;
      RECT 43.82 161.1 44.02 161.22 ;
      RECT 41.66 163.62 41.86 163.74 ;
      RECT 43.82 163.62 44.02 163.74 ;
      RECT 42.74 162.6 42.94 162.72 ;
      RECT 41.3 162.6 41.5 162.72 ;
      RECT 41.3 165.12 41.5 165.24 ;
      RECT 42.74 164.88 42.94 165 ;
      RECT 43.1 163.86 43.3 163.98 ;
      RECT 42.38 163.86 42.58 163.98 ;
      RECT 42.38 166.38 42.58 166.5 ;
      RECT 41.66 166.38 41.86 166.5 ;
      RECT 43.82 166.14 44.02 166.26 ;
      RECT 43.1 166.14 43.3 166.26 ;
      RECT 42.74 167.64 42.94 167.76 ;
      RECT 41.3 167.64 41.5 167.76 ;
      RECT 43.82 168.9 44.02 169.02 ;
      RECT 42.38 168.9 42.58 169.02 ;
      RECT 41.66 168.66 41.86 168.78 ;
      RECT 43.1 168.66 43.3 168.78 ;
      RECT 42.74 169.92 42.94 170.04 ;
      RECT 41.3 169.92 41.5 170.04 ;
      RECT 43.1 171.42 43.3 171.54 ;
      RECT 41.66 171.42 41.86 171.54 ;
      RECT 42.38 171.18 42.58 171.3 ;
      RECT 43.82 171.18 44.02 171.3 ;
      RECT 42.74 172.68 42.94 172.8 ;
      RECT 41.3 172.44 41.5 172.56 ;
      RECT 43.82 173.94 44.02 174.06 ;
      RECT 41.66 173.94 41.86 174.06 ;
      RECT 42.38 173.7 42.58 173.82 ;
      RECT 43.1 173.7 43.3 173.82 ;
      RECT 41.3 175.2 41.5 175.32 ;
      RECT 42.74 174.96 42.94 175.08 ;
      RECT 43.1 176.46 43.3 176.58 ;
      RECT 42.38 176.46 42.58 176.58 ;
      RECT 41.66 176.46 41.86 176.58 ;
      RECT 43.82 176.22 44.02 176.34 ;
      RECT 43.1 178.74 43.3 178.86 ;
      RECT 41.66 178.74 41.86 178.86 ;
      RECT 42.74 177.72 42.94 177.84 ;
      RECT 41.3 177.72 41.5 177.84 ;
      RECT 43.82 178.98 44.02 179.1 ;
      RECT 42.38 178.98 42.58 179.1 ;
      RECT 42.38 181.5 42.58 181.62 ;
      RECT 43.82 181.5 44.02 181.62 ;
      RECT 43.1 181.26 43.3 181.38 ;
      RECT 41.66 181.26 41.86 181.38 ;
      RECT 42.74 180.24 42.94 180.36 ;
      RECT 41.3 180.24 41.5 180.36 ;
      RECT 42.74 182.52 42.94 182.64 ;
      RECT 41.3 182.52 41.5 182.64 ;
      RECT 43.82 184.02 44.02 184.14 ;
      RECT 43.1 184.02 43.3 184.14 ;
      RECT 41.66 184.02 41.86 184.14 ;
      RECT 42.38 183.78 42.58 183.9 ;
      RECT 41.3 185.28 41.5 185.4 ;
      RECT 42.74 185.04 42.94 185.16 ;
      RECT 41.66 186.54 41.86 186.66 ;
      RECT 42.38 186.54 42.58 186.66 ;
      RECT 43.82 186.54 44.02 186.66 ;
      RECT 43.1 186.3 43.3 186.42 ;
      RECT 41.3 187.8 41.5 187.92 ;
      RECT 42.74 187.56 42.94 187.68 ;
      RECT 42.38 189.06 42.58 189.18 ;
      RECT 43.82 189.06 44.02 189.18 ;
      RECT 43.1 188.82 43.3 188.94 ;
      RECT 43.1 118.978 43.3 119.098 ;
      RECT 42.38 118.978 42.58 119.098 ;
      RECT 41.66 118.978 41.86 119.098 ;
      RECT 42.74 119.76 42.94 119.88 ;
      RECT 41.3 119.76 41.5 119.88 ;
      RECT 43.1 120.78 43.3 120.9 ;
      RECT 41.66 120.78 41.86 120.9 ;
      RECT 43.82 121.02 44.02 121.14 ;
      RECT 42.38 121.02 42.58 121.14 ;
      RECT 43.82 121.498 44.02 121.618 ;
      RECT 43.1 121.498 43.3 121.618 ;
      RECT 42.38 121.498 42.58 121.618 ;
      RECT 41.66 121.498 41.86 121.618 ;
      RECT 42.74 122.28 42.94 122.4 ;
      RECT 41.3 122.28 41.5 122.4 ;
      RECT 43.82 123.3 44.02 123.42 ;
      RECT 43.1 123.3 43.3 123.42 ;
      RECT 42.38 123.54 42.58 123.66 ;
      RECT 41.66 123.54 41.86 123.66 ;
      RECT 43.82 124.018 44.02 124.138 ;
      RECT 43.1 124.018 43.3 124.138 ;
      RECT 42.38 124.018 42.58 124.138 ;
      RECT 41.66 124.018 41.86 124.138 ;
      RECT 42.74 124.56 42.94 124.68 ;
      RECT 41.3 124.56 41.5 124.68 ;
      RECT 43.1 125.82 43.3 125.94 ;
      RECT 42.38 125.82 42.58 125.94 ;
      RECT 41.66 125.82 41.86 125.94 ;
      RECT 43.82 126.06 44.02 126.18 ;
      RECT 43.82 126.538 44.02 126.658 ;
      RECT 43.1 126.538 43.3 126.658 ;
      RECT 42.38 126.538 42.58 126.658 ;
      RECT 41.66 126.538 41.86 126.658 ;
      RECT 42.74 127.08 42.94 127.2 ;
      RECT 41.3 127.32 41.5 127.44 ;
      RECT 42.38 128.34 42.58 128.46 ;
      RECT 43.1 128.34 43.3 128.46 ;
      RECT 41.66 128.58 41.86 128.7 ;
      RECT 43.82 128.58 44.02 128.7 ;
      RECT 43.82 129.058 44.02 129.178 ;
      RECT 43.1 129.058 43.3 129.178 ;
      RECT 42.38 129.058 42.58 129.178 ;
      RECT 41.66 129.058 41.86 129.178 ;
      RECT 42.74 129.6 42.94 129.72 ;
      RECT 41.3 129.84 41.5 129.96 ;
      RECT 43.82 130.86 44.02 130.98 ;
      RECT 43.1 130.86 43.3 130.98 ;
      RECT 42.38 130.86 42.58 130.98 ;
      RECT 41.66 131.1 41.86 131.22 ;
      RECT 43.82 131.578 44.02 131.698 ;
      RECT 43.1 131.578 43.3 131.698 ;
      RECT 42.38 131.578 42.58 131.698 ;
      RECT 41.66 131.578 41.86 131.698 ;
      RECT 41.3 132.36 41.5 132.48 ;
      RECT 42.74 132.36 42.94 132.48 ;
      RECT 42.38 133.38 42.58 133.5 ;
      RECT 43.82 133.38 44.02 133.5 ;
      RECT 43.1 133.62 43.3 133.74 ;
      RECT 41.66 133.62 41.86 133.74 ;
      RECT 43.82 134.098 44.02 134.218 ;
      RECT 43.1 134.098 43.3 134.218 ;
      RECT 42.38 134.098 42.58 134.218 ;
      RECT 41.66 134.098 41.86 134.218 ;
      RECT 42.74 134.64 42.94 134.76 ;
      RECT 41.3 134.88 41.5 135 ;
      RECT 41.66 135.9 41.86 136.02 ;
      RECT 43.82 135.9 44.02 136.02 ;
      RECT 42.38 136.14 42.58 136.26 ;
      RECT 43.1 136.14 43.3 136.26 ;
      RECT 43.82 136.618 44.02 136.738 ;
      RECT 43.1 136.618 43.3 136.738 ;
      RECT 42.38 136.618 42.58 136.738 ;
      RECT 41.66 136.618 41.86 136.738 ;
      RECT 42.74 137.16 42.94 137.28 ;
      RECT 41.3 137.4 41.5 137.52 ;
      RECT 43.1 138.42 43.3 138.54 ;
      RECT 41.66 138.42 41.86 138.54 ;
      RECT 42.38 138.66 42.58 138.78 ;
      RECT 43.82 138.66 44.02 138.78 ;
      RECT 43.82 139.138 44.02 139.258 ;
      RECT 43.1 139.138 43.3 139.258 ;
      RECT 42.38 139.138 42.58 139.258 ;
      RECT 41.66 139.138 41.86 139.258 ;
      RECT 42.74 139.68 42.94 139.8 ;
      RECT 41.3 139.92 41.5 140.04 ;
      RECT 43.1 140.94 43.3 141.06 ;
      RECT 41.66 141.18 41.86 141.3 ;
      RECT 42.38 141.18 42.58 141.3 ;
      RECT 43.82 141.18 44.02 141.3 ;
      RECT 41.3 142.44 41.5 142.56 ;
      RECT 42.74 142.44 42.94 142.56 ;
      RECT 43.1 143.7 43.3 143.82 ;
      RECT 41.66 143.7 41.86 143.82 ;
      RECT 42.38 143.46 42.58 143.58 ;
      RECT 43.82 143.46 44.02 143.58 ;
      RECT 41.66 145.98 41.86 146.1 ;
      RECT 42.38 145.98 42.58 146.1 ;
      RECT 43.1 145.98 43.3 146.1 ;
      RECT 43.82 145.98 44.02 146.1 ;
      RECT 42.74 144.96 42.94 145.08 ;
      RECT 41.3 144.72 41.5 144.84 ;
      RECT 41.66 148.74 41.86 148.86 ;
      RECT 40.58 263.01 40.78 263.13 ;
      RECT 37.7 263.01 37.9 263.13 ;
      RECT 40.94 262.38 41.14 262.5 ;
      RECT 40.22 262.38 40.42 262.5 ;
      RECT 38.06 262.38 38.26 262.5 ;
      RECT 37.34 262.38 37.54 262.5 ;
      RECT 40.58 264.27 40.78 264.39 ;
      RECT 37.7 264.27 37.9 264.39 ;
      RECT 40.94 263.64 41.14 263.76 ;
      RECT 40.22 263.64 40.42 263.76 ;
      RECT 38.06 263.64 38.26 263.76 ;
      RECT 37.34 263.64 37.54 263.76 ;
      RECT 40.94 266.16 41.14 266.28 ;
      RECT 40.22 266.16 40.42 266.28 ;
      RECT 38.06 266.16 38.26 266.28 ;
      RECT 37.34 266.16 37.54 266.28 ;
      RECT 40.58 265.53 40.78 265.65 ;
      RECT 37.7 265.53 37.9 265.65 ;
      RECT 40.94 264.9 41.14 265.02 ;
      RECT 40.22 264.9 40.42 265.02 ;
      RECT 38.06 264.9 38.26 265.02 ;
      RECT 37.34 264.9 37.54 265.02 ;
      RECT 40.94 267.42 41.14 267.54 ;
      RECT 40.22 267.42 40.42 267.54 ;
      RECT 38.06 267.42 38.26 267.54 ;
      RECT 37.34 267.42 37.54 267.54 ;
      RECT 40.58 266.79 40.78 266.91 ;
      RECT 37.7 266.79 37.9 266.91 ;
      RECT 40.94 268.68 41.14 268.8 ;
      RECT 40.22 268.68 40.42 268.8 ;
      RECT 38.06 268.68 38.26 268.8 ;
      RECT 37.34 268.68 37.54 268.8 ;
      RECT 40.58 268.05 40.78 268.17 ;
      RECT 37.7 268.05 37.9 268.17 ;
      RECT 40.94 269.94 41.14 270.06 ;
      RECT 40.22 269.94 40.42 270.06 ;
      RECT 38.06 269.94 38.26 270.06 ;
      RECT 37.34 269.94 37.54 270.06 ;
      RECT 40.58 269.31 40.78 269.43 ;
      RECT 37.7 269.31 37.9 269.43 ;
      RECT 40.94 271.2 41.14 271.32 ;
      RECT 40.22 271.2 40.42 271.32 ;
      RECT 38.06 271.2 38.26 271.32 ;
      RECT 37.34 271.2 37.54 271.32 ;
      RECT 40.58 270.57 40.78 270.69 ;
      RECT 37.7 270.57 37.9 270.69 ;
      RECT 37.7 271.83 37.9 271.95 ;
      RECT 40.58 271.83 40.78 271.95 ;
      RECT 37.34 272.46 37.54 272.58 ;
      RECT 38.06 272.46 38.26 272.58 ;
      RECT 40.22 272.46 40.42 272.58 ;
      RECT 40.94 272.46 41.14 272.58 ;
      RECT 37.7 273.09 37.9 273.21 ;
      RECT 40.58 273.09 40.78 273.21 ;
      RECT 40.94 273.72 41.14 273.84 ;
      RECT 37.34 273.72 37.54 273.84 ;
      RECT 38.06 273.72 38.26 273.84 ;
      RECT 40.22 273.72 40.42 273.84 ;
      RECT 37.7 274.35 37.9 274.47 ;
      RECT 40.58 274.35 40.78 274.47 ;
      RECT 37.34 274.98 37.54 275.1 ;
      RECT 38.06 274.98 38.26 275.1 ;
      RECT 40.22 274.98 40.42 275.1 ;
      RECT 40.94 274.98 41.14 275.1 ;
      RECT 37.7 275.61 37.9 275.73 ;
      RECT 40.58 275.61 40.78 275.73 ;
      RECT 37.34 276.24 37.54 276.36 ;
      RECT 38.06 276.24 38.26 276.36 ;
      RECT 40.22 276.24 40.42 276.36 ;
      RECT 40.94 276.24 41.14 276.36 ;
      RECT 37.7 276.87 37.9 276.99 ;
      RECT 40.58 276.87 40.78 276.99 ;
      RECT 37.34 277.5 37.54 277.62 ;
      RECT 38.06 277.5 38.26 277.62 ;
      RECT 40.22 277.5 40.42 277.62 ;
      RECT 40.94 277.5 41.14 277.62 ;
      RECT 37.7 278.13 37.9 278.25 ;
      RECT 40.58 278.13 40.78 278.25 ;
      RECT 37.34 278.76 37.54 278.88 ;
      RECT 38.06 278.76 38.26 278.88 ;
      RECT 40.22 278.76 40.42 278.88 ;
      RECT 40.94 278.76 41.14 278.88 ;
      RECT 37.34 283.087 37.54 283.207 ;
      RECT 38.06 283.087 38.26 283.207 ;
      RECT 40.22 283.087 40.42 283.207 ;
      RECT 40.94 283.087 41.14 283.207 ;
      RECT 36.98 305.498 37.18 305.618 ;
      RECT 40.94 305.967 41.14 306.087 ;
      RECT 40.22 305.967 40.42 306.087 ;
      RECT 38.06 305.967 38.26 306.087 ;
      RECT 37.34 305.967 37.54 306.087 ;
      RECT 36.98 323.3835 37.18 323.5035 ;
      RECT 40.94 325.9425 41.14 326.0625 ;
      RECT 40.22 325.9425 40.42 326.0625 ;
      RECT 38.06 325.9425 38.26 326.0625 ;
      RECT 37.34 325.9425 37.54 326.0625 ;
      RECT 36.98 348.339 37.18 348.459 ;
      RECT 43.82 118.26 44.02 118.38 ;
      RECT 41.66 118.5 41.86 118.62 ;
      RECT 42.38 118.5 42.58 118.62 ;
      RECT 43.1 118.5 43.3 118.62 ;
      RECT 43.82 118.978 44.02 119.098 ;
      RECT 37.34 240.96 37.54 241.08 ;
      RECT 38.06 240.96 38.26 241.08 ;
      RECT 40.22 240.96 40.42 241.08 ;
      RECT 40.94 240.96 41.14 241.08 ;
      RECT 37.7 240.33 37.9 240.45 ;
      RECT 40.58 240.33 40.78 240.45 ;
      RECT 40.58 242.85 40.78 242.97 ;
      RECT 37.7 242.85 37.9 242.97 ;
      RECT 40.22 242.22 40.42 242.34 ;
      RECT 38.06 242.22 38.26 242.34 ;
      RECT 37.34 242.22 37.54 242.34 ;
      RECT 40.94 242.22 41.14 242.34 ;
      RECT 40.58 244.11 40.78 244.23 ;
      RECT 37.7 244.11 37.9 244.23 ;
      RECT 40.94 243.48 41.14 243.6 ;
      RECT 40.22 243.48 40.42 243.6 ;
      RECT 38.06 243.48 38.26 243.6 ;
      RECT 37.34 243.48 37.54 243.6 ;
      RECT 37.7 245.37 37.9 245.49 ;
      RECT 40.58 245.37 40.78 245.49 ;
      RECT 37.34 244.74 37.54 244.86 ;
      RECT 38.06 244.74 38.26 244.86 ;
      RECT 40.22 244.74 40.42 244.86 ;
      RECT 40.94 244.74 41.14 244.86 ;
      RECT 37.34 246 37.54 246.12 ;
      RECT 38.06 246 38.26 246.12 ;
      RECT 40.22 246 40.42 246.12 ;
      RECT 40.94 246 41.14 246.12 ;
      RECT 37.7 246.63 37.9 246.75 ;
      RECT 40.58 246.63 40.78 246.75 ;
      RECT 37.34 247.26 37.54 247.38 ;
      RECT 38.06 247.26 38.26 247.38 ;
      RECT 40.22 247.26 40.42 247.38 ;
      RECT 40.94 247.26 41.14 247.38 ;
      RECT 37.7 247.89 37.9 248.01 ;
      RECT 40.58 247.89 40.78 248.01 ;
      RECT 37.34 248.52 37.54 248.64 ;
      RECT 38.06 248.52 38.26 248.64 ;
      RECT 40.22 248.52 40.42 248.64 ;
      RECT 40.94 248.52 41.14 248.64 ;
      RECT 37.7 249.15 37.9 249.27 ;
      RECT 40.58 249.15 40.78 249.27 ;
      RECT 37.34 249.78 37.54 249.9 ;
      RECT 38.06 249.78 38.26 249.9 ;
      RECT 40.22 249.78 40.42 249.9 ;
      RECT 40.94 249.78 41.14 249.9 ;
      RECT 37.7 250.41 37.9 250.53 ;
      RECT 40.58 250.41 40.78 250.53 ;
      RECT 37.34 251.04 37.54 251.16 ;
      RECT 38.06 251.04 38.26 251.16 ;
      RECT 40.22 251.04 40.42 251.16 ;
      RECT 40.94 251.04 41.14 251.16 ;
      RECT 37.7 251.67 37.9 251.79 ;
      RECT 40.58 251.67 40.78 251.79 ;
      RECT 37.34 252.3 37.54 252.42 ;
      RECT 38.06 252.3 38.26 252.42 ;
      RECT 40.22 252.3 40.42 252.42 ;
      RECT 40.94 252.3 41.14 252.42 ;
      RECT 37.7 252.93 37.9 253.05 ;
      RECT 40.58 252.93 40.78 253.05 ;
      RECT 37.34 253.56 37.54 253.68 ;
      RECT 38.06 253.56 38.26 253.68 ;
      RECT 40.22 253.56 40.42 253.68 ;
      RECT 40.94 253.56 41.14 253.68 ;
      RECT 37.7 254.19 37.9 254.31 ;
      RECT 40.58 254.19 40.78 254.31 ;
      RECT 37.34 254.82 37.54 254.94 ;
      RECT 38.06 254.82 38.26 254.94 ;
      RECT 40.22 254.82 40.42 254.94 ;
      RECT 40.94 254.82 41.14 254.94 ;
      RECT 37.7 255.45 37.9 255.57 ;
      RECT 40.58 255.45 40.78 255.57 ;
      RECT 37.34 256.08 37.54 256.2 ;
      RECT 38.06 256.08 38.26 256.2 ;
      RECT 40.22 256.08 40.42 256.2 ;
      RECT 40.94 256.08 41.14 256.2 ;
      RECT 37.7 256.71 37.9 256.83 ;
      RECT 40.58 256.71 40.78 256.83 ;
      RECT 37.34 257.34 37.54 257.46 ;
      RECT 38.06 257.34 38.26 257.46 ;
      RECT 40.22 257.34 40.42 257.46 ;
      RECT 40.94 257.34 41.14 257.46 ;
      RECT 37.7 257.97 37.9 258.09 ;
      RECT 40.58 257.97 40.78 258.09 ;
      RECT 40.58 259.23 40.78 259.35 ;
      RECT 37.7 259.23 37.9 259.35 ;
      RECT 37.34 258.6 37.54 258.72 ;
      RECT 38.06 258.6 38.26 258.72 ;
      RECT 40.22 258.6 40.42 258.72 ;
      RECT 40.94 258.6 41.14 258.72 ;
      RECT 40.58 260.49 40.78 260.61 ;
      RECT 37.7 260.49 37.9 260.61 ;
      RECT 40.94 259.86 41.14 259.98 ;
      RECT 40.22 259.86 40.42 259.98 ;
      RECT 38.06 259.86 38.26 259.98 ;
      RECT 37.34 259.86 37.54 259.98 ;
      RECT 40.58 261.75 40.78 261.87 ;
      RECT 37.7 261.75 37.9 261.87 ;
      RECT 40.94 261.12 41.14 261.24 ;
      RECT 40.22 261.12 40.42 261.24 ;
      RECT 38.06 261.12 38.26 261.24 ;
      RECT 37.34 261.12 37.54 261.24 ;
      RECT 38.06 219.54 38.26 219.66 ;
      RECT 37.34 219.54 37.54 219.66 ;
      RECT 37.7 218.91 37.9 219.03 ;
      RECT 40.58 218.91 40.78 219.03 ;
      RECT 37.7 220.17 37.9 220.29 ;
      RECT 40.58 220.17 40.78 220.29 ;
      RECT 37.34 220.8 37.54 220.92 ;
      RECT 38.06 220.8 38.26 220.92 ;
      RECT 40.22 220.8 40.42 220.92 ;
      RECT 40.94 220.8 41.14 220.92 ;
      RECT 37.34 222.06 37.54 222.18 ;
      RECT 38.06 222.06 38.26 222.18 ;
      RECT 40.22 222.06 40.42 222.18 ;
      RECT 40.94 222.06 41.14 222.18 ;
      RECT 40.58 221.43 40.78 221.55 ;
      RECT 37.7 221.43 37.9 221.55 ;
      RECT 37.34 223.32 37.54 223.44 ;
      RECT 38.06 223.32 38.26 223.44 ;
      RECT 40.22 223.32 40.42 223.44 ;
      RECT 40.94 223.32 41.14 223.44 ;
      RECT 37.7 222.69 37.9 222.81 ;
      RECT 40.58 222.69 40.78 222.81 ;
      RECT 37.7 225.21 37.9 225.33 ;
      RECT 40.58 225.21 40.78 225.33 ;
      RECT 37.34 224.58 37.54 224.7 ;
      RECT 38.06 224.58 38.26 224.7 ;
      RECT 40.22 224.58 40.42 224.7 ;
      RECT 40.94 224.58 41.14 224.7 ;
      RECT 37.7 223.95 37.9 224.07 ;
      RECT 40.58 223.95 40.78 224.07 ;
      RECT 37.7 226.47 37.9 226.59 ;
      RECT 40.58 226.47 40.78 226.59 ;
      RECT 37.34 225.84 37.54 225.96 ;
      RECT 38.06 225.84 38.26 225.96 ;
      RECT 40.22 225.84 40.42 225.96 ;
      RECT 40.94 225.84 41.14 225.96 ;
      RECT 37.7 227.73 37.9 227.85 ;
      RECT 40.58 227.73 40.78 227.85 ;
      RECT 37.34 227.1 37.54 227.22 ;
      RECT 38.06 227.1 38.26 227.22 ;
      RECT 40.22 227.1 40.42 227.22 ;
      RECT 40.94 227.1 41.14 227.22 ;
      RECT 37.7 228.99 37.9 229.11 ;
      RECT 40.58 228.99 40.78 229.11 ;
      RECT 37.34 228.36 37.54 228.48 ;
      RECT 38.06 228.36 38.26 228.48 ;
      RECT 40.22 228.36 40.42 228.48 ;
      RECT 40.94 228.36 41.14 228.48 ;
      RECT 40.58 230.25 40.78 230.37 ;
      RECT 37.7 230.25 37.9 230.37 ;
      RECT 37.34 229.62 37.54 229.74 ;
      RECT 38.06 229.62 38.26 229.74 ;
      RECT 40.22 229.62 40.42 229.74 ;
      RECT 40.94 229.62 41.14 229.74 ;
      RECT 40.58 231.51 40.78 231.63 ;
      RECT 37.7 231.51 37.9 231.63 ;
      RECT 40.94 230.88 41.14 231 ;
      RECT 40.22 230.88 40.42 231 ;
      RECT 38.06 230.88 38.26 231 ;
      RECT 37.34 230.88 37.54 231 ;
      RECT 37.34 233.4 37.54 233.52 ;
      RECT 38.06 233.4 38.26 233.52 ;
      RECT 40.22 233.4 40.42 233.52 ;
      RECT 40.94 233.4 41.14 233.52 ;
      RECT 40.58 232.77 40.78 232.89 ;
      RECT 37.7 232.77 37.9 232.89 ;
      RECT 40.94 232.14 41.14 232.26 ;
      RECT 40.22 232.14 40.42 232.26 ;
      RECT 38.06 232.14 38.26 232.26 ;
      RECT 37.34 232.14 37.54 232.26 ;
      RECT 40.94 234.66 41.14 234.78 ;
      RECT 40.22 234.66 40.42 234.78 ;
      RECT 38.06 234.66 38.26 234.78 ;
      RECT 37.34 234.66 37.54 234.78 ;
      RECT 37.7 234.03 37.9 234.15 ;
      RECT 40.58 234.03 40.78 234.15 ;
      RECT 40.94 235.92 41.14 236.04 ;
      RECT 40.22 235.92 40.42 236.04 ;
      RECT 38.06 235.92 38.26 236.04 ;
      RECT 37.34 235.92 37.54 236.04 ;
      RECT 40.58 235.29 40.78 235.41 ;
      RECT 37.7 235.29 37.9 235.41 ;
      RECT 37.34 237.18 37.54 237.3 ;
      RECT 38.06 237.18 38.26 237.3 ;
      RECT 40.22 237.18 40.42 237.3 ;
      RECT 40.94 237.18 41.14 237.3 ;
      RECT 40.58 236.55 40.78 236.67 ;
      RECT 37.7 236.55 37.9 236.67 ;
      RECT 40.94 238.44 41.14 238.56 ;
      RECT 40.22 238.44 40.42 238.56 ;
      RECT 38.06 238.44 38.26 238.56 ;
      RECT 37.34 238.44 37.54 238.56 ;
      RECT 37.7 237.81 37.9 237.93 ;
      RECT 40.58 237.81 40.78 237.93 ;
      RECT 40.94 239.7 41.14 239.82 ;
      RECT 40.22 239.7 40.42 239.82 ;
      RECT 38.06 239.7 38.26 239.82 ;
      RECT 37.34 239.7 37.54 239.82 ;
      RECT 40.58 239.07 40.78 239.19 ;
      RECT 37.7 239.07 37.9 239.19 ;
      RECT 37.7 241.59 37.9 241.71 ;
      RECT 40.58 241.59 40.78 241.71 ;
      RECT 36.98 190.08 37.18 190.2 ;
      RECT 37.7 192.122 37.9 192.242 ;
      RECT 40.58 192.122 40.78 192.242 ;
      RECT 38.06 191.58 38.26 191.7 ;
      RECT 37.34 191.58 37.54 191.7 ;
      RECT 40.22 191.34 40.42 191.46 ;
      RECT 40.94 191.34 41.14 191.46 ;
      RECT 37.7 193.382 37.9 193.502 ;
      RECT 40.58 193.142 40.78 193.262 ;
      RECT 36.98 192.84 37.18 192.96 ;
      RECT 37.7 194.642 37.9 194.762 ;
      RECT 40.58 194.402 40.78 194.522 ;
      RECT 38.06 194.1 38.26 194.22 ;
      RECT 37.34 194.1 37.54 194.22 ;
      RECT 40.22 193.86 40.42 193.98 ;
      RECT 40.94 193.86 41.14 193.98 ;
      RECT 37.34 196.38 37.54 196.5 ;
      RECT 40.22 196.38 40.42 196.5 ;
      RECT 40.58 195.902 40.78 196.022 ;
      RECT 37.7 195.662 37.9 195.782 ;
      RECT 36.98 195.36 37.18 195.48 ;
      RECT 36.98 197.64 37.18 197.76 ;
      RECT 40.94 196.62 41.14 196.74 ;
      RECT 38.06 196.62 38.26 196.74 ;
      RECT 37.34 199.14 37.54 199.26 ;
      RECT 38.06 199.14 38.26 199.26 ;
      RECT 40.94 198.9 41.14 199.02 ;
      RECT 40.22 198.9 40.42 199.02 ;
      RECT 37.7 198.422 37.9 198.542 ;
      RECT 40.58 198.422 40.78 198.542 ;
      RECT 36.98 200.16 37.18 200.28 ;
      RECT 40.94 201.66 41.14 201.78 ;
      RECT 38.06 201.66 38.26 201.78 ;
      RECT 37.34 201.42 37.54 201.54 ;
      RECT 40.22 201.42 40.42 201.54 ;
      RECT 40.58 200.942 40.78 201.062 ;
      RECT 37.7 200.702 37.9 200.822 ;
      RECT 37.7 203.222 37.9 203.342 ;
      RECT 36.98 202.92 37.18 203.04 ;
      RECT 37.34 204.18 37.54 204.3 ;
      RECT 40.94 204.18 41.14 204.3 ;
      RECT 40.22 203.94 40.42 204.06 ;
      RECT 38.06 203.94 38.26 204.06 ;
      RECT 40.58 203.462 40.78 203.582 ;
      RECT 40.58 205.982 40.78 206.102 ;
      RECT 37.7 205.742 37.9 205.862 ;
      RECT 36.98 205.2 37.18 205.32 ;
      RECT 40.94 206.7 41.14 206.82 ;
      RECT 38.06 206.7 38.26 206.82 ;
      RECT 40.22 206.46 40.42 206.58 ;
      RECT 37.34 206.46 37.54 206.58 ;
      RECT 40.58 208.502 40.78 208.622 ;
      RECT 37.7 208.262 37.9 208.382 ;
      RECT 36.98 207.72 37.18 207.84 ;
      RECT 37.7 210.09 37.9 210.21 ;
      RECT 40.58 210.09 40.78 210.21 ;
      RECT 40.94 209.46 41.14 209.58 ;
      RECT 40.22 209.46 40.42 209.58 ;
      RECT 38.06 209.46 38.26 209.58 ;
      RECT 37.34 209.46 37.54 209.58 ;
      RECT 37.7 211.35 37.9 211.47 ;
      RECT 40.58 211.35 40.78 211.47 ;
      RECT 37.34 210.72 37.54 210.84 ;
      RECT 38.06 210.72 38.26 210.84 ;
      RECT 40.22 210.72 40.42 210.84 ;
      RECT 40.94 210.72 41.14 210.84 ;
      RECT 37.7 212.61 37.9 212.73 ;
      RECT 40.58 212.61 40.78 212.73 ;
      RECT 40.94 211.98 41.14 212.1 ;
      RECT 40.22 211.98 40.42 212.1 ;
      RECT 38.06 211.98 38.26 212.1 ;
      RECT 37.34 211.98 37.54 212.1 ;
      RECT 37.7 213.87 37.9 213.99 ;
      RECT 40.58 213.87 40.78 213.99 ;
      RECT 37.34 213.24 37.54 213.36 ;
      RECT 38.06 213.24 38.26 213.36 ;
      RECT 40.22 213.24 40.42 213.36 ;
      RECT 40.94 213.24 41.14 213.36 ;
      RECT 37.7 215.13 37.9 215.25 ;
      RECT 40.58 215.13 40.78 215.25 ;
      RECT 37.34 214.5 37.54 214.62 ;
      RECT 38.06 214.5 38.26 214.62 ;
      RECT 40.22 214.5 40.42 214.62 ;
      RECT 40.94 214.5 41.14 214.62 ;
      RECT 37.34 217.02 37.54 217.14 ;
      RECT 38.06 217.02 38.26 217.14 ;
      RECT 40.22 217.02 40.42 217.14 ;
      RECT 40.94 217.02 41.14 217.14 ;
      RECT 40.58 216.39 40.78 216.51 ;
      RECT 37.7 216.39 37.9 216.51 ;
      RECT 37.34 215.76 37.54 215.88 ;
      RECT 38.06 215.76 38.26 215.88 ;
      RECT 40.22 215.76 40.42 215.88 ;
      RECT 40.94 215.76 41.14 215.88 ;
      RECT 37.34 218.28 37.54 218.4 ;
      RECT 38.06 218.28 38.26 218.4 ;
      RECT 40.22 218.28 40.42 218.4 ;
      RECT 40.94 218.28 41.14 218.4 ;
      RECT 37.7 217.65 37.9 217.77 ;
      RECT 40.58 217.65 40.78 217.77 ;
      RECT 40.94 219.54 41.14 219.66 ;
      RECT 40.22 219.54 40.42 219.66 ;
      RECT 37.34 141.18 37.54 141.3 ;
      RECT 40.22 141.18 40.42 141.3 ;
      RECT 36.98 142.2 37.18 142.32 ;
      RECT 40.22 143.7 40.42 143.82 ;
      RECT 38.06 143.7 38.26 143.82 ;
      RECT 37.34 143.46 37.54 143.58 ;
      RECT 40.94 143.46 41.14 143.58 ;
      RECT 37.34 145.98 37.54 146.1 ;
      RECT 38.06 145.98 38.26 146.1 ;
      RECT 40.22 145.98 40.42 146.1 ;
      RECT 40.94 145.98 41.14 146.1 ;
      RECT 36.98 144.96 37.18 145.08 ;
      RECT 37.34 148.74 37.54 148.86 ;
      RECT 40.22 148.74 40.42 148.86 ;
      RECT 40.94 148.74 41.14 148.86 ;
      RECT 38.06 148.5 38.26 148.62 ;
      RECT 36.98 149.76 37.18 149.88 ;
      RECT 40.94 151.26 41.14 151.38 ;
      RECT 40.22 151.26 40.42 151.38 ;
      RECT 38.06 151.26 38.26 151.38 ;
      RECT 37.34 151.02 37.54 151.14 ;
      RECT 36.98 152.52 37.18 152.64 ;
      RECT 40.22 153.78 40.42 153.9 ;
      RECT 38.06 153.78 38.26 153.9 ;
      RECT 40.94 153.54 41.14 153.66 ;
      RECT 37.34 153.54 37.54 153.66 ;
      RECT 36.98 155.04 37.18 155.16 ;
      RECT 40.58 156.842 40.78 156.962 ;
      RECT 37.7 156.602 37.9 156.722 ;
      RECT 38.06 156.3 38.26 156.42 ;
      RECT 40.94 156.3 41.14 156.42 ;
      RECT 40.22 156.06 40.42 156.18 ;
      RECT 37.34 156.06 37.54 156.18 ;
      RECT 40.58 158.278 40.78 158.398 ;
      RECT 37.7 158.038 37.9 158.158 ;
      RECT 36.98 157.56 37.18 157.68 ;
      RECT 40.94 158.82 41.14 158.94 ;
      RECT 37.34 158.82 37.54 158.94 ;
      RECT 38.06 158.58 38.26 158.7 ;
      RECT 40.22 158.58 40.42 158.7 ;
      RECT 36.98 159.84 37.18 159.96 ;
      RECT 37.34 161.1 37.54 161.22 ;
      RECT 38.06 161.1 38.26 161.22 ;
      RECT 40.22 161.1 40.42 161.22 ;
      RECT 40.94 161.1 41.14 161.22 ;
      RECT 37.34 163.62 37.54 163.74 ;
      RECT 36.98 162.6 37.18 162.72 ;
      RECT 36.98 165.12 37.18 165.24 ;
      RECT 40.94 163.86 41.14 163.98 ;
      RECT 40.22 163.86 40.42 163.98 ;
      RECT 38.06 163.86 38.26 163.98 ;
      RECT 37.34 166.38 37.54 166.5 ;
      RECT 40.94 166.14 41.14 166.26 ;
      RECT 40.22 166.14 40.42 166.26 ;
      RECT 38.06 166.14 38.26 166.26 ;
      RECT 36.98 167.4 37.18 167.52 ;
      RECT 40.94 168.9 41.14 169.02 ;
      RECT 40.22 168.9 40.42 169.02 ;
      RECT 37.34 168.9 37.54 169.02 ;
      RECT 38.06 168.66 38.26 168.78 ;
      RECT 36.98 170.16 37.18 170.28 ;
      RECT 40.22 171.42 40.42 171.54 ;
      RECT 38.06 171.42 38.26 171.54 ;
      RECT 37.34 171.42 37.54 171.54 ;
      RECT 40.94 171.18 41.14 171.3 ;
      RECT 36.98 172.68 37.18 172.8 ;
      RECT 40.94 173.94 41.14 174.06 ;
      RECT 38.06 173.94 38.26 174.06 ;
      RECT 40.22 173.7 40.42 173.82 ;
      RECT 37.34 173.7 37.54 173.82 ;
      RECT 36.98 174.96 37.18 175.08 ;
      RECT 40.94 176.46 41.14 176.58 ;
      RECT 40.22 176.46 40.42 176.58 ;
      RECT 38.06 176.22 38.26 176.34 ;
      RECT 37.34 176.22 37.54 176.34 ;
      RECT 40.94 178.74 41.14 178.86 ;
      RECT 36.98 177.48 37.18 177.6 ;
      RECT 36.98 180 37.18 180.12 ;
      RECT 37.34 178.98 37.54 179.1 ;
      RECT 40.22 178.98 40.42 179.1 ;
      RECT 38.06 178.98 38.26 179.1 ;
      RECT 38.06 181.5 38.26 181.62 ;
      RECT 40.22 181.5 40.42 181.62 ;
      RECT 40.94 181.26 41.14 181.38 ;
      RECT 37.34 181.26 37.54 181.38 ;
      RECT 36.98 182.52 37.18 182.64 ;
      RECT 40.22 184.02 40.42 184.14 ;
      RECT 37.34 184.02 37.54 184.14 ;
      RECT 40.94 183.78 41.14 183.9 ;
      RECT 38.06 183.78 38.26 183.9 ;
      RECT 36.98 185.28 37.18 185.4 ;
      RECT 37.34 186.54 37.54 186.66 ;
      RECT 40.22 186.54 40.42 186.66 ;
      RECT 38.06 186.3 38.26 186.42 ;
      RECT 40.94 186.3 41.14 186.42 ;
      RECT 36.98 187.8 37.18 187.92 ;
      RECT 38.06 189.06 38.26 189.18 ;
      RECT 40.94 189.06 41.14 189.18 ;
      RECT 40.22 188.82 40.42 188.94 ;
      RECT 37.34 188.82 37.54 188.94 ;
      RECT 37.7 190.862 37.9 190.982 ;
      RECT 40.58 190.622 40.78 190.742 ;
      RECT 34.46 278.76 34.66 278.88 ;
      RECT 35.18 278.76 35.38 278.88 ;
      RECT 35.9 278.76 36.1 278.88 ;
      RECT 36.62 278.76 36.82 278.88 ;
      RECT 34.46 283.087 34.66 283.207 ;
      RECT 35.18 283.087 35.38 283.207 ;
      RECT 35.9 283.087 36.1 283.207 ;
      RECT 36.62 283.087 36.82 283.207 ;
      RECT 35.54 305.498 35.74 305.618 ;
      RECT 36.62 305.967 36.82 306.087 ;
      RECT 35.9 305.967 36.1 306.087 ;
      RECT 35.18 305.967 35.38 306.087 ;
      RECT 34.46 305.967 34.66 306.087 ;
      RECT 35.54 323.3835 35.74 323.5035 ;
      RECT 36.62 325.9425 36.82 326.0625 ;
      RECT 35.9 325.9425 36.1 326.0625 ;
      RECT 35.18 325.9425 35.38 326.0625 ;
      RECT 34.46 325.9425 34.66 326.0625 ;
      RECT 35.54 348.339 35.74 348.459 ;
      RECT 37.34 118.26 37.54 118.38 ;
      RECT 38.06 118.26 38.26 118.38 ;
      RECT 40.94 118.26 41.14 118.38 ;
      RECT 40.22 118.5 40.42 118.62 ;
      RECT 40.94 118.978 41.14 119.098 ;
      RECT 40.22 118.978 40.42 119.098 ;
      RECT 38.06 118.978 38.26 119.098 ;
      RECT 37.34 118.978 37.54 119.098 ;
      RECT 36.98 119.52 37.18 119.64 ;
      RECT 40.22 120.78 40.42 120.9 ;
      RECT 38.06 120.78 38.26 120.9 ;
      RECT 40.94 121.02 41.14 121.14 ;
      RECT 37.34 121.02 37.54 121.14 ;
      RECT 40.94 121.498 41.14 121.618 ;
      RECT 40.22 121.498 40.42 121.618 ;
      RECT 38.06 121.498 38.26 121.618 ;
      RECT 37.34 121.498 37.54 121.618 ;
      RECT 36.98 122.28 37.18 122.4 ;
      RECT 40.94 123.3 41.14 123.42 ;
      RECT 38.06 123.3 38.26 123.42 ;
      RECT 37.34 123.54 37.54 123.66 ;
      RECT 40.22 123.54 40.42 123.66 ;
      RECT 40.94 124.018 41.14 124.138 ;
      RECT 40.22 124.018 40.42 124.138 ;
      RECT 38.06 124.018 38.26 124.138 ;
      RECT 37.34 124.018 37.54 124.138 ;
      RECT 36.98 124.8 37.18 124.92 ;
      RECT 40.94 125.82 41.14 125.94 ;
      RECT 40.22 126.06 40.42 126.18 ;
      RECT 38.06 126.06 38.26 126.18 ;
      RECT 37.34 126.06 37.54 126.18 ;
      RECT 40.94 126.538 41.14 126.658 ;
      RECT 40.22 126.538 40.42 126.658 ;
      RECT 38.06 126.538 38.26 126.658 ;
      RECT 37.34 126.538 37.54 126.658 ;
      RECT 36.98 127.08 37.18 127.2 ;
      RECT 38.06 128.34 38.26 128.46 ;
      RECT 40.22 128.34 40.42 128.46 ;
      RECT 37.34 128.58 37.54 128.7 ;
      RECT 40.94 128.58 41.14 128.7 ;
      RECT 40.94 129.058 41.14 129.178 ;
      RECT 40.22 129.058 40.42 129.178 ;
      RECT 38.06 129.058 38.26 129.178 ;
      RECT 37.34 129.058 37.54 129.178 ;
      RECT 36.98 129.6 37.18 129.72 ;
      RECT 40.22 130.86 40.42 130.98 ;
      RECT 37.34 131.1 37.54 131.22 ;
      RECT 38.06 131.1 38.26 131.22 ;
      RECT 40.94 131.1 41.14 131.22 ;
      RECT 40.94 131.578 41.14 131.698 ;
      RECT 40.22 131.578 40.42 131.698 ;
      RECT 38.06 131.578 38.26 131.698 ;
      RECT 37.34 131.578 37.54 131.698 ;
      RECT 36.98 132.12 37.18 132.24 ;
      RECT 38.06 133.38 38.26 133.5 ;
      RECT 40.22 133.38 40.42 133.5 ;
      RECT 40.94 133.62 41.14 133.74 ;
      RECT 37.34 133.62 37.54 133.74 ;
      RECT 40.94 134.098 41.14 134.218 ;
      RECT 40.22 134.098 40.42 134.218 ;
      RECT 38.06 134.098 38.26 134.218 ;
      RECT 37.34 134.098 37.54 134.218 ;
      RECT 36.98 134.88 37.18 135 ;
      RECT 38.06 135.9 38.26 136.02 ;
      RECT 40.22 135.9 40.42 136.02 ;
      RECT 40.94 136.14 41.14 136.26 ;
      RECT 37.34 136.14 37.54 136.26 ;
      RECT 40.94 136.618 41.14 136.738 ;
      RECT 40.22 136.618 40.42 136.738 ;
      RECT 38.06 136.618 38.26 136.738 ;
      RECT 37.34 136.618 37.54 136.738 ;
      RECT 36.98 137.16 37.18 137.28 ;
      RECT 38.06 138.42 38.26 138.54 ;
      RECT 40.94 138.42 41.14 138.54 ;
      RECT 37.34 138.66 37.54 138.78 ;
      RECT 40.22 138.66 40.42 138.78 ;
      RECT 40.94 139.138 41.14 139.258 ;
      RECT 40.22 139.138 40.42 139.258 ;
      RECT 38.06 139.138 38.26 139.258 ;
      RECT 37.34 139.138 37.54 139.258 ;
      RECT 36.98 139.92 37.18 140.04 ;
      RECT 40.94 140.94 41.14 141.06 ;
      RECT 38.06 140.94 38.26 141.06 ;
      RECT 34.46 257.34 34.66 257.46 ;
      RECT 35.18 257.34 35.38 257.46 ;
      RECT 35.9 257.34 36.1 257.46 ;
      RECT 36.62 257.34 36.82 257.46 ;
      RECT 34.82 257.97 35.02 258.09 ;
      RECT 36.26 257.97 36.46 258.09 ;
      RECT 34.46 258.6 34.66 258.72 ;
      RECT 35.18 258.6 35.38 258.72 ;
      RECT 35.9 258.6 36.1 258.72 ;
      RECT 36.62 258.6 36.82 258.72 ;
      RECT 34.82 259.23 35.02 259.35 ;
      RECT 36.26 259.23 36.46 259.35 ;
      RECT 36.26 260.49 36.46 260.61 ;
      RECT 34.82 260.49 35.02 260.61 ;
      RECT 36.62 259.86 36.82 259.98 ;
      RECT 35.9 259.86 36.1 259.98 ;
      RECT 35.18 259.86 35.38 259.98 ;
      RECT 34.46 259.86 34.66 259.98 ;
      RECT 36.26 261.75 36.46 261.87 ;
      RECT 34.82 261.75 35.02 261.87 ;
      RECT 36.62 261.12 36.82 261.24 ;
      RECT 35.9 261.12 36.1 261.24 ;
      RECT 35.18 261.12 35.38 261.24 ;
      RECT 34.46 261.12 34.66 261.24 ;
      RECT 36.26 263.01 36.46 263.13 ;
      RECT 34.82 263.01 35.02 263.13 ;
      RECT 36.62 262.38 36.82 262.5 ;
      RECT 35.9 262.38 36.1 262.5 ;
      RECT 35.18 262.38 35.38 262.5 ;
      RECT 34.46 262.38 34.66 262.5 ;
      RECT 36.26 264.27 36.46 264.39 ;
      RECT 34.82 264.27 35.02 264.39 ;
      RECT 36.62 263.64 36.82 263.76 ;
      RECT 35.9 263.64 36.1 263.76 ;
      RECT 35.18 263.64 35.38 263.76 ;
      RECT 34.46 263.64 34.66 263.76 ;
      RECT 36.62 266.16 36.82 266.28 ;
      RECT 35.9 266.16 36.1 266.28 ;
      RECT 35.18 266.16 35.38 266.28 ;
      RECT 34.46 266.16 34.66 266.28 ;
      RECT 36.26 265.53 36.46 265.65 ;
      RECT 34.82 265.53 35.02 265.65 ;
      RECT 36.62 264.9 36.82 265.02 ;
      RECT 35.9 264.9 36.1 265.02 ;
      RECT 35.18 264.9 35.38 265.02 ;
      RECT 34.46 264.9 34.66 265.02 ;
      RECT 36.62 267.42 36.82 267.54 ;
      RECT 35.9 267.42 36.1 267.54 ;
      RECT 35.18 267.42 35.38 267.54 ;
      RECT 34.46 267.42 34.66 267.54 ;
      RECT 36.26 266.79 36.46 266.91 ;
      RECT 34.82 266.79 35.02 266.91 ;
      RECT 36.62 268.68 36.82 268.8 ;
      RECT 35.9 268.68 36.1 268.8 ;
      RECT 35.18 268.68 35.38 268.8 ;
      RECT 34.46 268.68 34.66 268.8 ;
      RECT 36.26 268.05 36.46 268.17 ;
      RECT 34.82 268.05 35.02 268.17 ;
      RECT 36.62 269.94 36.82 270.06 ;
      RECT 35.9 269.94 36.1 270.06 ;
      RECT 35.18 269.94 35.38 270.06 ;
      RECT 34.46 269.94 34.66 270.06 ;
      RECT 36.26 269.31 36.46 269.43 ;
      RECT 34.82 269.31 35.02 269.43 ;
      RECT 36.62 271.2 36.82 271.32 ;
      RECT 35.9 271.2 36.1 271.32 ;
      RECT 35.18 271.2 35.38 271.32 ;
      RECT 34.46 271.2 34.66 271.32 ;
      RECT 36.26 270.57 36.46 270.69 ;
      RECT 34.82 270.57 35.02 270.69 ;
      RECT 36.26 271.83 36.46 271.95 ;
      RECT 34.82 271.83 35.02 271.95 ;
      RECT 35.9 272.46 36.1 272.58 ;
      RECT 36.62 272.46 36.82 272.58 ;
      RECT 34.46 272.46 34.66 272.58 ;
      RECT 35.18 272.46 35.38 272.58 ;
      RECT 34.82 273.09 35.02 273.21 ;
      RECT 36.26 273.09 36.46 273.21 ;
      RECT 34.46 273.72 34.66 273.84 ;
      RECT 35.18 273.72 35.38 273.84 ;
      RECT 35.9 273.72 36.1 273.84 ;
      RECT 36.62 273.72 36.82 273.84 ;
      RECT 34.82 274.35 35.02 274.47 ;
      RECT 36.26 274.35 36.46 274.47 ;
      RECT 34.46 274.98 34.66 275.1 ;
      RECT 35.18 274.98 35.38 275.1 ;
      RECT 35.9 274.98 36.1 275.1 ;
      RECT 36.62 274.98 36.82 275.1 ;
      RECT 34.82 275.61 35.02 275.73 ;
      RECT 36.26 275.61 36.46 275.73 ;
      RECT 34.46 276.24 34.66 276.36 ;
      RECT 35.18 276.24 35.38 276.36 ;
      RECT 35.9 276.24 36.1 276.36 ;
      RECT 36.62 276.24 36.82 276.36 ;
      RECT 34.82 276.87 35.02 276.99 ;
      RECT 36.26 276.87 36.46 276.99 ;
      RECT 35.18 277.5 35.38 277.62 ;
      RECT 34.46 277.5 34.66 277.62 ;
      RECT 35.9 277.5 36.1 277.62 ;
      RECT 36.62 277.5 36.82 277.62 ;
      RECT 34.82 278.13 35.02 278.25 ;
      RECT 36.26 278.13 36.46 278.25 ;
      RECT 35.18 235.92 35.38 236.04 ;
      RECT 34.46 235.92 34.66 236.04 ;
      RECT 36.26 235.29 36.46 235.41 ;
      RECT 34.82 235.29 35.02 235.41 ;
      RECT 34.46 237.18 34.66 237.3 ;
      RECT 35.18 237.18 35.38 237.3 ;
      RECT 35.9 237.18 36.1 237.3 ;
      RECT 36.62 237.18 36.82 237.3 ;
      RECT 36.26 236.55 36.46 236.67 ;
      RECT 34.82 236.55 35.02 236.67 ;
      RECT 36.62 238.44 36.82 238.56 ;
      RECT 35.9 238.44 36.1 238.56 ;
      RECT 35.18 238.44 35.38 238.56 ;
      RECT 34.46 238.44 34.66 238.56 ;
      RECT 34.82 237.81 35.02 237.93 ;
      RECT 36.26 237.81 36.46 237.93 ;
      RECT 36.62 239.7 36.82 239.82 ;
      RECT 35.9 239.7 36.1 239.82 ;
      RECT 35.18 239.7 35.38 239.82 ;
      RECT 34.46 239.7 34.66 239.82 ;
      RECT 36.26 239.07 36.46 239.19 ;
      RECT 34.82 239.07 35.02 239.19 ;
      RECT 34.82 241.59 35.02 241.71 ;
      RECT 36.26 241.59 36.46 241.71 ;
      RECT 34.46 240.96 34.66 241.08 ;
      RECT 35.18 240.96 35.38 241.08 ;
      RECT 35.9 240.96 36.1 241.08 ;
      RECT 36.62 240.96 36.82 241.08 ;
      RECT 36.26 240.33 36.46 240.45 ;
      RECT 34.82 240.33 35.02 240.45 ;
      RECT 36.26 242.85 36.46 242.97 ;
      RECT 34.82 242.85 35.02 242.97 ;
      RECT 36.62 242.22 36.82 242.34 ;
      RECT 35.9 242.22 36.1 242.34 ;
      RECT 35.18 242.22 35.38 242.34 ;
      RECT 34.46 242.22 34.66 242.34 ;
      RECT 36.26 244.11 36.46 244.23 ;
      RECT 34.82 244.11 35.02 244.23 ;
      RECT 36.62 243.48 36.82 243.6 ;
      RECT 35.9 243.48 36.1 243.6 ;
      RECT 35.18 243.48 35.38 243.6 ;
      RECT 34.46 243.48 34.66 243.6 ;
      RECT 34.82 245.37 35.02 245.49 ;
      RECT 36.26 245.37 36.46 245.49 ;
      RECT 34.46 244.74 34.66 244.86 ;
      RECT 35.18 244.74 35.38 244.86 ;
      RECT 35.9 244.74 36.1 244.86 ;
      RECT 36.62 244.74 36.82 244.86 ;
      RECT 34.46 246 34.66 246.12 ;
      RECT 35.18 246 35.38 246.12 ;
      RECT 35.9 246 36.1 246.12 ;
      RECT 36.62 246 36.82 246.12 ;
      RECT 34.82 246.63 35.02 246.75 ;
      RECT 36.26 246.63 36.46 246.75 ;
      RECT 34.46 247.26 34.66 247.38 ;
      RECT 35.18 247.26 35.38 247.38 ;
      RECT 35.9 247.26 36.1 247.38 ;
      RECT 36.62 247.26 36.82 247.38 ;
      RECT 34.82 247.89 35.02 248.01 ;
      RECT 36.26 247.89 36.46 248.01 ;
      RECT 34.46 248.52 34.66 248.64 ;
      RECT 35.18 248.52 35.38 248.64 ;
      RECT 35.9 248.52 36.1 248.64 ;
      RECT 36.62 248.52 36.82 248.64 ;
      RECT 34.82 249.15 35.02 249.27 ;
      RECT 36.26 249.15 36.46 249.27 ;
      RECT 34.46 249.78 34.66 249.9 ;
      RECT 35.18 249.78 35.38 249.9 ;
      RECT 35.9 249.78 36.1 249.9 ;
      RECT 36.62 249.78 36.82 249.9 ;
      RECT 34.82 250.41 35.02 250.53 ;
      RECT 36.26 250.41 36.46 250.53 ;
      RECT 34.46 251.04 34.66 251.16 ;
      RECT 35.18 251.04 35.38 251.16 ;
      RECT 35.9 251.04 36.1 251.16 ;
      RECT 36.62 251.04 36.82 251.16 ;
      RECT 34.82 251.67 35.02 251.79 ;
      RECT 36.26 251.67 36.46 251.79 ;
      RECT 34.46 252.3 34.66 252.42 ;
      RECT 35.18 252.3 35.38 252.42 ;
      RECT 35.9 252.3 36.1 252.42 ;
      RECT 36.62 252.3 36.82 252.42 ;
      RECT 34.82 252.93 35.02 253.05 ;
      RECT 36.26 252.93 36.46 253.05 ;
      RECT 34.46 253.56 34.66 253.68 ;
      RECT 35.18 253.56 35.38 253.68 ;
      RECT 35.9 253.56 36.1 253.68 ;
      RECT 36.62 253.56 36.82 253.68 ;
      RECT 34.82 254.19 35.02 254.31 ;
      RECT 36.26 254.19 36.46 254.31 ;
      RECT 34.46 254.82 34.66 254.94 ;
      RECT 35.18 254.82 35.38 254.94 ;
      RECT 35.9 254.82 36.1 254.94 ;
      RECT 36.62 254.82 36.82 254.94 ;
      RECT 34.82 255.45 35.02 255.57 ;
      RECT 36.26 255.45 36.46 255.57 ;
      RECT 34.46 256.08 34.66 256.2 ;
      RECT 35.18 256.08 35.38 256.2 ;
      RECT 35.9 256.08 36.1 256.2 ;
      RECT 36.62 256.08 36.82 256.2 ;
      RECT 36.26 256.71 36.46 256.83 ;
      RECT 34.82 256.71 35.02 256.83 ;
      RECT 34.82 215.13 35.02 215.25 ;
      RECT 36.26 215.13 36.46 215.25 ;
      RECT 36.62 214.5 36.82 214.62 ;
      RECT 35.9 214.5 36.1 214.62 ;
      RECT 35.18 214.5 35.38 214.62 ;
      RECT 34.46 214.5 34.66 214.62 ;
      RECT 34.46 217.02 34.66 217.14 ;
      RECT 35.18 217.02 35.38 217.14 ;
      RECT 35.9 217.02 36.1 217.14 ;
      RECT 36.62 217.02 36.82 217.14 ;
      RECT 36.26 216.39 36.46 216.51 ;
      RECT 34.82 216.39 35.02 216.51 ;
      RECT 34.46 215.76 34.66 215.88 ;
      RECT 35.18 215.76 35.38 215.88 ;
      RECT 35.9 215.76 36.1 215.88 ;
      RECT 36.62 215.76 36.82 215.88 ;
      RECT 34.46 218.28 34.66 218.4 ;
      RECT 35.18 218.28 35.38 218.4 ;
      RECT 35.9 218.28 36.1 218.4 ;
      RECT 36.62 218.28 36.82 218.4 ;
      RECT 34.82 217.65 35.02 217.77 ;
      RECT 36.26 217.65 36.46 217.77 ;
      RECT 36.62 219.54 36.82 219.66 ;
      RECT 35.9 219.54 36.1 219.66 ;
      RECT 35.18 219.54 35.38 219.66 ;
      RECT 34.46 219.54 34.66 219.66 ;
      RECT 34.82 218.91 35.02 219.03 ;
      RECT 36.26 218.91 36.46 219.03 ;
      RECT 36.26 220.17 36.46 220.29 ;
      RECT 34.82 220.17 35.02 220.29 ;
      RECT 34.46 220.8 34.66 220.92 ;
      RECT 35.18 220.8 35.38 220.92 ;
      RECT 35.9 220.8 36.1 220.92 ;
      RECT 36.62 220.8 36.82 220.92 ;
      RECT 34.46 222.06 34.66 222.18 ;
      RECT 35.18 222.06 35.38 222.18 ;
      RECT 35.9 222.06 36.1 222.18 ;
      RECT 36.62 222.06 36.82 222.18 ;
      RECT 36.26 221.43 36.46 221.55 ;
      RECT 34.82 221.43 35.02 221.55 ;
      RECT 34.46 223.32 34.66 223.44 ;
      RECT 35.18 223.32 35.38 223.44 ;
      RECT 35.9 223.32 36.1 223.44 ;
      RECT 36.62 223.32 36.82 223.44 ;
      RECT 34.82 222.69 35.02 222.81 ;
      RECT 36.26 222.69 36.46 222.81 ;
      RECT 34.82 225.21 35.02 225.33 ;
      RECT 36.26 225.21 36.46 225.33 ;
      RECT 34.46 224.58 34.66 224.7 ;
      RECT 35.18 224.58 35.38 224.7 ;
      RECT 35.9 224.58 36.1 224.7 ;
      RECT 36.62 224.58 36.82 224.7 ;
      RECT 34.82 223.95 35.02 224.07 ;
      RECT 36.26 223.95 36.46 224.07 ;
      RECT 34.82 226.47 35.02 226.59 ;
      RECT 36.26 226.47 36.46 226.59 ;
      RECT 34.46 225.84 34.66 225.96 ;
      RECT 35.18 225.84 35.38 225.96 ;
      RECT 35.9 225.84 36.1 225.96 ;
      RECT 36.62 225.84 36.82 225.96 ;
      RECT 34.82 227.73 35.02 227.85 ;
      RECT 36.26 227.73 36.46 227.85 ;
      RECT 34.46 227.1 34.66 227.22 ;
      RECT 35.18 227.1 35.38 227.22 ;
      RECT 35.9 227.1 36.1 227.22 ;
      RECT 36.62 227.1 36.82 227.22 ;
      RECT 34.82 228.99 35.02 229.11 ;
      RECT 36.26 228.99 36.46 229.11 ;
      RECT 34.46 228.36 34.66 228.48 ;
      RECT 35.18 228.36 35.38 228.48 ;
      RECT 35.9 228.36 36.1 228.48 ;
      RECT 36.62 228.36 36.82 228.48 ;
      RECT 36.26 230.25 36.46 230.37 ;
      RECT 34.82 230.25 35.02 230.37 ;
      RECT 34.46 229.62 34.66 229.74 ;
      RECT 35.18 229.62 35.38 229.74 ;
      RECT 35.9 229.62 36.1 229.74 ;
      RECT 36.62 229.62 36.82 229.74 ;
      RECT 36.26 231.51 36.46 231.63 ;
      RECT 34.82 231.51 35.02 231.63 ;
      RECT 36.62 230.88 36.82 231 ;
      RECT 35.9 230.88 36.1 231 ;
      RECT 35.18 230.88 35.38 231 ;
      RECT 34.46 230.88 34.66 231 ;
      RECT 34.46 233.4 34.66 233.52 ;
      RECT 35.18 233.4 35.38 233.52 ;
      RECT 35.9 233.4 36.1 233.52 ;
      RECT 36.62 233.4 36.82 233.52 ;
      RECT 36.26 232.77 36.46 232.89 ;
      RECT 34.82 232.77 35.02 232.89 ;
      RECT 36.62 232.14 36.82 232.26 ;
      RECT 35.9 232.14 36.1 232.26 ;
      RECT 35.18 232.14 35.38 232.26 ;
      RECT 34.46 232.14 34.66 232.26 ;
      RECT 36.62 234.66 36.82 234.78 ;
      RECT 35.9 234.66 36.1 234.78 ;
      RECT 35.18 234.66 35.38 234.78 ;
      RECT 34.46 234.66 34.66 234.78 ;
      RECT 34.82 234.03 35.02 234.15 ;
      RECT 36.26 234.03 36.46 234.15 ;
      RECT 36.62 235.92 36.82 236.04 ;
      RECT 35.9 235.92 36.1 236.04 ;
  END
END ringpll

END LIBRARY
