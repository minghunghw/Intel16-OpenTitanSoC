## ##############################################################################
## ## Intel Top Secret                                                         ##
## ##############################################################################
## ## Copyright © Intel Corporation.                                           ##
## ##                                                                          ##
## ## This is the property of Intel Corporation and may only be utilized       ##
## ## pursuant to a written Restricted Use Nondisclosure Agreement             ##
## ## with Intel Corporation.  It may not be used, reproduced, or              ##
## ## disclosed to others except in accordance with the terms and              ##
## ## conditions of such agreement.                                            ##
## ##                                                                          ##
## ## All products, processes, computer systems, dates, and figures            ##
## ## specified are preliminary based on current expectations, and are         ##
## ## subject to change without notice.                                        ##
## ##############################################################################
## ## Text_Tag % __Placeholder neutral1


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO b15qbfbf1bn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qbfbf1bn1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
      ANTENNAMAXAREACAR 6.0805555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
      ANTENNAMAXAREACAR 6.0805555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.222 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER m2 ;
        RECT 0.472 0.338 0.916 0.382 ;
      LAYER v1 ;
        RECT 0.726 0.338 0.786 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNADIFFAREA 0.04896 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 1.006 0.202 ;
        RECT 0.398 0.158 0.466 0.562 ;
        RECT 0.506 0.428 1.006 0.472 ;
      LAYER m2 ;
        RECT 0.488 0.158 0.916 0.202 ;
        RECT 0.272 0.428 0.916 0.472 ;
      LAYER v1 ;
        RECT 0.402 0.428 0.462 0.472 ;
        RECT 0.618 0.428 0.678 0.472 ;
        RECT 0.618 0.158 0.678 0.202 ;
        RECT 0.834 0.428 0.894 0.472 ;
        RECT 0.834 0.158 0.894 0.202 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
    END
  END o
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
        RECT 0.29 0.338 0.358 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.338 0.392 0.382 ;
      LAYER v1 ;
        RECT 0.186 0.338 0.246 0.382 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.363 0.142 0.407 ;
        RECT 0.182 0.498 0.25 0.542 ;
        RECT 0.182 0.363 0.25 0.407 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.363 0.358 0.407 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  OBS
    LAYER m2 ;
      RECT 1.352 0.428 1.564 0.472 ;
      RECT 1.352 0.158 1.564 0.202 ;
    LAYER m1 ;
      RECT 0.506 0.428 1.006 0.472 ;
      RECT 0.614 0.338 1.154 0.382 ;
      RECT 0.614 0.248 1.046 0.292 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.586 0.068 1.654 0.292 ;
    LAYER v1 ;
      RECT 1.482 0.158 1.542 0.202 ;
      RECT 1.482 0.428 1.542 0.472 ;
    LAYER v0 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.223 1.654 0.267 ;
      RECT 1.586 0.358 1.654 0.402 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.478 0.088 1.546 0.132 ;
      RECT 1.478 0.223 1.546 0.267 ;
      RECT 1.478 0.358 1.546 0.402 ;
      RECT 1.478 0.498 1.546 0.542 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.223 1.438 0.267 ;
      RECT 1.37 0.358 1.438 0.402 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.722 0.248 0.79 0.292 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.158 1.006 0.202 ;
      RECT 1.154 0.158 1.222 0.382 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.046 0.518 1.262 0.562 ;
      RECT 1.114 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.562 ;
  END
END b15qbfbf1bn1n16x5

MACRO b15qbfbf1bn1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qbfbf1bn1n32x5 0 0 ;
  SIZE 2.376 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
      ANTENNAMAXAREACAR 1.52222225 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.391111 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
      ANTENNAMAXAREACAR 1.52222225 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.391111 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER m2 ;
        RECT 0.364 0.338 1.024 0.382 ;
      LAYER v1 ;
        RECT 0.51 0.338 0.57 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05814 LAYER m1 ;
    ANTENNADIFFAREA 0.11628 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.978 0.202 ;
        RECT 0.938 0.158 1.006 0.562 ;
        RECT 1.046 0.428 1.978 0.472 ;
      LAYER m2 ;
        RECT 1.136 0.158 1.904 0.202 ;
        RECT 0.92 0.428 1.904 0.472 ;
      LAYER v1 ;
        RECT 0.942 0.428 1.002 0.472 ;
        RECT 1.158 0.428 1.218 0.472 ;
        RECT 1.158 0.158 1.218 0.202 ;
        RECT 1.374 0.428 1.434 0.472 ;
        RECT 1.374 0.158 1.434 0.202 ;
        RECT 1.59 0.428 1.65 0.472 ;
        RECT 1.59 0.158 1.65 0.202 ;
        RECT 1.806 0.428 1.866 0.472 ;
        RECT 1.806 0.158 1.866 0.202 ;
      LAYER v0 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
    END
  END o
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.41 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
        RECT 0.29 0.338 0.358 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.338 0.284 0.382 ;
      LAYER v1 ;
        RECT 0.186 0.338 0.246 0.382 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.363 0.142 0.407 ;
        RECT 0.182 0.498 0.25 0.542 ;
        RECT 0.182 0.363 0.25 0.407 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.363 0.358 0.407 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.41 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 1.046 0.538 1.114 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
    END
  END vcc
  OBS
    LAYER m2 ;
      RECT 1.984 0.428 2.212 0.472 ;
      RECT 1.984 0.158 2.212 0.202 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.046 0.428 1.978 0.472 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 2.234 0.068 2.302 0.292 ;
    LAYER v1 ;
      RECT 2.13 0.158 2.19 0.202 ;
      RECT 2.13 0.428 2.19 0.472 ;
    LAYER v0 ;
      RECT 2.234 0.088 2.302 0.132 ;
      RECT 2.234 0.223 2.302 0.267 ;
      RECT 2.234 0.358 2.302 0.402 ;
      RECT 2.234 0.498 2.302 0.542 ;
      RECT 2.126 0.088 2.194 0.132 ;
      RECT 2.126 0.223 2.194 0.267 ;
      RECT 2.126 0.358 2.194 0.402 ;
      RECT 2.126 0.498 2.194 0.542 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 2.018 0.223 2.086 0.267 ;
      RECT 2.018 0.358 2.086 0.402 ;
      RECT 2.018 0.498 2.086 0.542 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.616 0.4385 0.68 0.4825 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 1.006 0.158 1.978 0.202 ;
  END
END b15qbfbf1bn1n32x5

MACRO b15qbfff4gn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qbfff4gn1n08x5 0 0 ;
  SIZE 7.452 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0054 LAYER m2 ;
      ANTENNAMAXAREACAR 3.515 LAYER m1 ;
      ANTENNAMAXAREACAR 8.6024075 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0054 LAYER m2 ;
      ANTENNAMAXAREACAR 3.515 LAYER m1 ;
      ANTENNAMAXAREACAR 8.6024075 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.158 1.546 0.562 ;
      LAYER m2 ;
        RECT 1.028 0.428 1.58 0.472 ;
      LAYER v1 ;
        RECT 1.482 0.428 1.542 0.472 ;
      LAYER v0 ;
        RECT 1.478 0.498 1.546 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.472 ;
      LAYER m2 ;
        RECT 1.012 0.158 1.456 0.202 ;
      LAYER v1 ;
        RECT 1.158 0.158 1.218 0.202 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    ANTENNADIFFAREA 0.02448 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 6.554 0.158 6.946 0.202 ;
        RECT 6.554 0.158 6.622 0.562 ;
        RECT 6.77 0.338 6.838 0.562 ;
      LAYER m2 ;
        RECT 6.536 0.158 6.98 0.202 ;
        RECT 6.536 0.518 6.98 0.562 ;
      LAYER v1 ;
        RECT 6.558 0.518 6.618 0.562 ;
        RECT 6.774 0.518 6.834 0.562 ;
        RECT 6.774 0.158 6.834 0.202 ;
      LAYER v0 ;
        RECT 6.77 0.448 6.838 0.492 ;
        RECT 6.77 0.158 6.838 0.202 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 24.5444445 LAYER m2 ;
      ANTENNAMAXCUTCAR 2.29777775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 24.5444445 LAYER m2 ;
      ANTENNAMAXCUTCAR 2.29777775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.042 0.068 5.11 0.562 ;
        RECT 2.666 0.518 2.95 0.562 ;
      LAYER m2 ;
        RECT 4.808 0.068 5.252 0.112 ;
        RECT 2.756 0.518 5.128 0.562 ;
      LAYER v1 ;
        RECT 2.778 0.518 2.838 0.562 ;
        RECT 5.046 0.518 5.106 0.562 ;
        RECT 5.046 0.068 5.106 0.112 ;
      LAYER v0 ;
        RECT 2.774 0.518 2.842 0.562 ;
        RECT 5.042 0.248 5.11 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.068 4.678 0.382 ;
        RECT 3.942 0.338 4.246 0.382 ;
      LAYER m2 ;
        RECT 4.16 0.338 4.696 0.382 ;
      LAYER v1 ;
        RECT 4.182 0.338 4.242 0.382 ;
        RECT 4.614 0.338 4.674 0.382 ;
      LAYER v0 ;
        RECT 4.07 0.338 4.138 0.382 ;
        RECT 4.61 0.088 4.678 0.132 ;
    END
  END rb
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 7.486 0.022 ;
        RECT 6.878 -0.022 6.946 0.112 ;
        RECT 6.662 -0.022 6.73 0.112 ;
        RECT 6.446 -0.022 6.514 0.202 ;
        RECT 5.15 -0.022 5.218 0.202 ;
        RECT 4.718 -0.022 4.786 0.292 ;
        RECT 2.558 0.158 3.726 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.262 -0.022 1.33 0.292 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.29 0.338 0.358 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.596 0.158 0.932 0.202 ;
        RECT 0.164 0.428 0.376 0.472 ;
      LAYER v1 ;
        RECT 0.186 0.428 0.246 0.472 ;
        RECT 0.726 0.158 0.786 0.202 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.363 0.142 0.407 ;
        RECT 0.182 0.498 0.25 0.542 ;
        RECT 0.182 0.363 0.25 0.407 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.363 0.358 0.407 ;
        RECT 0.614 0.223 0.682 0.267 ;
        RECT 0.614 0.088 0.682 0.132 ;
        RECT 0.722 0.223 0.79 0.267 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 0.83 0.223 0.898 0.267 ;
        RECT 0.83 0.088 0.898 0.132 ;
        RECT 1.262 0.203 1.33 0.247 ;
        RECT 1.91 0.048 1.978 0.092 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.206 0.158 3.274 0.202 ;
        RECT 3.422 0.158 3.49 0.202 ;
        RECT 3.638 0.158 3.706 0.202 ;
        RECT 4.718 0.203 4.786 0.247 ;
        RECT 5.15 0.138 5.218 0.182 ;
        RECT 6.446 0.138 6.514 0.182 ;
        RECT 6.664 0.048 6.728 0.092 ;
        RECT 6.88 0.048 6.944 0.092 ;
    END
  END vssx
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 7.486 0.652 ;
        RECT 6.878 0.428 6.946 0.652 ;
        RECT 6.662 0.518 6.73 0.652 ;
        RECT 6.446 0.338 6.514 0.652 ;
        RECT 5.15 0.428 5.218 0.652 ;
        RECT 4.934 0.428 5.002 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.206 0.338 3.274 0.652 ;
        RECT 2.99 0.338 3.058 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.262 0.338 1.33 0.652 ;
      LAYER v0 ;
        RECT 1.262 0.408 1.33 0.452 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.99 0.3835 3.058 0.4275 ;
        RECT 3.208 0.428 3.272 0.472 ;
        RECT 3.962 0.538 4.03 0.582 ;
        RECT 4.61 0.448 4.678 0.492 ;
        RECT 4.934 0.448 5.002 0.492 ;
        RECT 5.15 0.448 5.218 0.492 ;
        RECT 6.446 0.428 6.514 0.472 ;
        RECT 6.664 0.538 6.728 0.582 ;
        RECT 6.878 0.448 6.946 0.492 ;
    END
  END vcc
  OBS
    LAYER m2 ;
      RECT 1.028 0.338 2.12 0.382 ;
      RECT 1.352 0.518 2.32 0.562 ;
      RECT 2.2 0.338 3.616 0.382 ;
      RECT 1.66 0.428 4.28 0.472 ;
      RECT 5.332 0.068 5.684 0.112 ;
      RECT 5.78 0.338 6.1 0.382 ;
      RECT 4.36 0.428 6.748 0.472 ;
      RECT 7.06 0.518 7.288 0.562 ;
      RECT 7.06 0.158 7.288 0.202 ;
    LAYER m1 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.91 0.248 1.978 0.382 ;
      RECT 2.234 0.158 2.302 0.472 ;
      RECT 2.342 0.248 2.41 0.472 ;
      RECT 2.234 0.518 2.43 0.562 ;
      RECT 2.558 0.248 2.626 0.472 ;
      RECT 2.666 0.518 2.95 0.562 ;
      RECT 3.422 0.338 3.834 0.382 ;
      RECT 3.942 0.338 4.246 0.382 ;
      RECT 4.07 0.428 4.286 0.472 ;
      RECT 4.178 0.158 4.394 0.202 ;
      RECT 2.774 0.068 4.502 0.112 ;
      RECT 4.826 0.248 4.894 0.562 ;
      RECT 4.61 0.068 4.678 0.382 ;
      RECT 4.718 0.428 4.786 0.562 ;
      RECT 6.554 0.158 6.622 0.562 ;
      RECT 5.042 0.068 5.11 0.562 ;
      RECT 5.366 0.068 5.434 0.292 ;
      RECT 5.474 0.068 5.542 0.292 ;
      RECT 5.582 0.068 5.65 0.292 ;
      RECT 5.906 0.338 5.974 0.562 ;
      RECT 6.014 0.338 6.082 0.562 ;
      RECT 6.122 0.338 6.19 0.562 ;
      RECT 6.338 0.068 6.406 0.562 ;
      RECT 6.662 0.248 6.73 0.472 ;
      RECT 6.77 0.338 6.838 0.562 ;
      RECT 7.094 0.338 7.162 0.562 ;
      RECT 7.094 0.068 7.162 0.292 ;
      RECT 7.202 0.338 7.27 0.562 ;
      RECT 7.202 0.068 7.27 0.292 ;
      RECT 7.31 0.338 7.378 0.562 ;
      RECT 7.31 0.068 7.378 0.292 ;
    LAYER v1 ;
      RECT 7.206 0.158 7.266 0.202 ;
      RECT 7.206 0.518 7.266 0.562 ;
      RECT 6.666 0.428 6.726 0.472 ;
      RECT 6.018 0.338 6.078 0.382 ;
      RECT 5.478 0.068 5.538 0.112 ;
      RECT 4.722 0.428 4.782 0.472 ;
      RECT 4.398 0.428 4.458 0.472 ;
      RECT 4.182 0.428 4.242 0.472 ;
      RECT 3.534 0.338 3.594 0.382 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 2.238 0.518 2.298 0.562 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 1.05 0.338 1.11 0.382 ;
    LAYER v0 ;
      RECT 7.31 0.088 7.378 0.132 ;
      RECT 7.31 0.223 7.378 0.267 ;
      RECT 7.31 0.358 7.378 0.402 ;
      RECT 7.31 0.498 7.378 0.542 ;
      RECT 7.202 0.088 7.27 0.132 ;
      RECT 7.202 0.223 7.27 0.267 ;
      RECT 7.202 0.358 7.27 0.402 ;
      RECT 7.202 0.498 7.27 0.542 ;
      RECT 7.094 0.088 7.162 0.132 ;
      RECT 7.094 0.223 7.162 0.267 ;
      RECT 7.094 0.358 7.162 0.402 ;
      RECT 7.094 0.498 7.162 0.542 ;
      RECT 6.662 0.338 6.73 0.382 ;
      RECT 6.338 0.138 6.406 0.182 ;
      RECT 6.338 0.428 6.406 0.472 ;
      RECT 6.122 0.363 6.19 0.407 ;
      RECT 6.122 0.498 6.19 0.542 ;
      RECT 6.014 0.363 6.082 0.407 ;
      RECT 6.014 0.498 6.082 0.542 ;
      RECT 5.906 0.363 5.974 0.407 ;
      RECT 5.906 0.498 5.974 0.542 ;
      RECT 5.582 0.088 5.65 0.132 ;
      RECT 5.582 0.223 5.65 0.267 ;
      RECT 5.474 0.088 5.542 0.132 ;
      RECT 5.474 0.223 5.542 0.267 ;
      RECT 5.366 0.088 5.434 0.132 ;
      RECT 5.366 0.223 5.434 0.267 ;
      RECT 4.934 0.138 5.002 0.182 ;
      RECT 4.826 0.448 4.894 0.492 ;
      RECT 4.718 0.448 4.786 0.492 ;
      RECT 4.502 0.338 4.57 0.382 ;
      RECT 4.394 0.068 4.462 0.112 ;
      RECT 4.394 0.428 4.462 0.472 ;
      RECT 4.286 0.158 4.354 0.202 ;
      RECT 4.286 0.338 4.354 0.382 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 3.854 0.248 3.922 0.292 ;
      RECT 3.854 0.428 3.922 0.472 ;
      RECT 3.746 0.338 3.814 0.382 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.558 0.293 2.626 0.337 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.342 0.518 2.41 0.562 ;
      RECT 2.234 0.3835 2.302 0.4275 ;
      RECT 2.128 0.088 2.192 0.132 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.37 0.408 1.438 0.452 ;
      RECT 1.046 0.203 1.114 0.247 ;
      RECT 1.046 0.4055 1.114 0.4495 ;
    LAYER m1 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.438 0.068 1.694 0.112 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.762 0.158 2.126 0.202 ;
      RECT 2.126 0.068 2.194 0.202 ;
      RECT 2.302 0.158 2.518 0.202 ;
      RECT 2.626 0.428 2.882 0.472 ;
      RECT 2.882 0.248 2.95 0.472 ;
      RECT 2.95 0.248 3.314 0.292 ;
      RECT 3.314 0.248 3.382 0.472 ;
      RECT 3.382 0.428 4.03 0.472 ;
      RECT 3.382 0.248 4.246 0.292 ;
      RECT 4.286 0.248 4.354 0.472 ;
      RECT 4.394 0.158 4.462 0.562 ;
      RECT 4.502 0.068 4.57 0.472 ;
      RECT 4.894 0.248 4.934 0.292 ;
      RECT 4.934 0.068 5.002 0.292 ;
      RECT 6.622 0.158 6.946 0.202 ;
  END
END b15qbfff4gn1n08x5

MACRO b15qbfin1bn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qbfin1bn1n16x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAGATEAREA 0.0288 LAYER m2 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
      ANTENNAMAXAREACAR 1.122639 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.1955555 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAGATEAREA 0.0288 LAYER m2 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
      ANTENNAMAXAREACAR 1.122639 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.1955555 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER m2 ;
        RECT 0.472 0.428 0.916 0.472 ;
      LAYER v1 ;
        RECT 0.51 0.428 0.57 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNADIFFAREA 0.04896 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 1.006 0.202 ;
        RECT 0.398 0.158 0.466 0.562 ;
        RECT 0.83 0.338 0.898 0.562 ;
        RECT 0.614 0.338 0.898 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.158 0.916 0.202 ;
        RECT 0.38 0.518 0.916 0.562 ;
      LAYER v1 ;
        RECT 0.402 0.518 0.462 0.562 ;
        RECT 0.618 0.518 0.678 0.562 ;
        RECT 0.618 0.158 0.678 0.202 ;
        RECT 0.834 0.518 0.894 0.562 ;
        RECT 0.834 0.158 0.894 0.202 ;
      LAYER v0 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 0.83 0.158 0.898 0.202 ;
    END
  END o1
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
        RECT 0.29 0.338 0.358 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.428 0.392 0.472 ;
      LAYER v1 ;
        RECT 0.186 0.428 0.246 0.472 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.363 0.142 0.407 ;
        RECT 0.182 0.498 0.25 0.542 ;
        RECT 0.182 0.363 0.25 0.407 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.363 0.358 0.407 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
    END
  END vssx
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.938 0.538 1.006 0.582 ;
    END
  END vcc
  OBS
    LAYER m2 ;
      RECT 1.244 0.518 1.472 0.562 ;
      RECT 1.244 0.158 1.472 0.202 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.262 0.068 1.33 0.292 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.292 ;
    LAYER v1 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.266 0.518 1.326 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.223 1.438 0.267 ;
      RECT 1.37 0.358 1.438 0.402 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.262 0.088 1.33 0.132 ;
      RECT 1.262 0.223 1.33 0.267 ;
      RECT 1.262 0.358 1.33 0.402 ;
      RECT 1.262 0.498 1.33 0.542 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.223 1.222 0.267 ;
      RECT 1.154 0.358 1.222 0.402 ;
      RECT 1.154 0.498 1.222 0.542 ;
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.466 0.158 1.006 0.202 ;
  END
END b15qbfin1bn1n16x5

MACRO b15qbfin1bn1n40x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qbfin1bn1n40x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.072 LAYER m1 ;
      ANTENNAGATEAREA 0.072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.5795 LAYER m1 ;
      ANTENNAMAXAREACAR 0.96327775 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.23466675 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.072 LAYER m1 ;
      ANTENNAGATEAREA 0.072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.5795 LAYER m1 ;
      ANTENNAMAXAREACAR 0.96327775 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.23466675 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.674 0.292 ;
      LAYER m2 ;
        RECT 0.92 0.248 1.672 0.292 ;
      LAYER v1 ;
        RECT 1.158 0.248 1.218 0.292 ;
        RECT 1.374 0.248 1.434 0.292 ;
        RECT 1.59 0.248 1.65 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.586 0.248 1.654 0.292 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    ANTENNADIFFAREA 0.1224 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 1.654 0.202 ;
        RECT 0.938 0.158 1.006 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
        RECT 0.506 0.428 1.654 0.472 ;
        RECT 1.586 0.338 1.654 0.472 ;
        RECT 1.37 0.338 1.438 0.472 ;
        RECT 1.154 0.338 1.222 0.472 ;
      LAYER m2 ;
        RECT 0.488 0.338 1.796 0.382 ;
        RECT 0.596 0.158 1.58 0.202 ;
      LAYER v1 ;
        RECT 0.51 0.338 0.57 0.382 ;
        RECT 0.618 0.158 0.678 0.202 ;
        RECT 0.726 0.338 0.786 0.382 ;
        RECT 0.834 0.158 0.894 0.202 ;
        RECT 0.942 0.338 1.002 0.382 ;
        RECT 1.05 0.158 1.11 0.202 ;
        RECT 1.158 0.338 1.218 0.382 ;
        RECT 1.266 0.158 1.326 0.202 ;
        RECT 1.374 0.338 1.434 0.382 ;
        RECT 1.482 0.158 1.542 0.202 ;
        RECT 1.59 0.338 1.65 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END o1
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
        RECT 0.29 0.338 0.358 0.562 ;
        RECT 0.182 0.248 0.25 0.562 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.248 0.268 0.292 ;
      LAYER v1 ;
        RECT 0.186 0.248 0.246 0.292 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.363 0.142 0.407 ;
        RECT 0.182 0.498 0.25 0.542 ;
        RECT 0.182 0.363 0.25 0.407 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.363 0.358 0.407 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
    END
  END vssx
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  OBS
    LAYER m2 ;
      RECT 1.66 0.158 1.996 0.202 ;
      RECT 1.876 0.338 2.12 0.382 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 1.046 0.248 1.674 0.292 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.91 0.068 1.978 0.292 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.018 0.068 2.086 0.292 ;
    LAYER v1 ;
      RECT 1.914 0.158 1.974 0.202 ;
      RECT 1.914 0.338 1.974 0.382 ;
    LAYER v0 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 2.018 0.223 2.086 0.267 ;
      RECT 2.018 0.358 2.086 0.402 ;
      RECT 2.018 0.498 2.086 0.542 ;
      RECT 1.91 0.088 1.978 0.132 ;
      RECT 1.91 0.223 1.978 0.267 ;
      RECT 1.91 0.358 1.978 0.402 ;
      RECT 1.91 0.498 1.978 0.542 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.223 1.87 0.267 ;
      RECT 1.802 0.358 1.87 0.402 ;
      RECT 1.802 0.498 1.87 0.542 ;
    LAYER m1 ;
      RECT 0.506 0.428 1.154 0.472 ;
      RECT 1.154 0.338 1.222 0.472 ;
      RECT 1.222 0.428 1.37 0.472 ;
      RECT 1.37 0.338 1.438 0.472 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.338 1.654 0.472 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 0.79 0.158 0.938 0.202 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.006 0.158 1.654 0.202 ;
  END
END b15qbfin1bn1n40x5

MACRO b15qbflf4gn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qbflf4gn1n08x5 0 0 ;
  SIZE 4.536 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 3.15 LAYER m1 ;
      ANTENNAMAXAREACAR 7.0555555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 6.3 LAYER m1 ;
      ANTENNAMAXAREACAR 14.111111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.338 1.762 0.562 ;
        RECT 0.938 0.248 1.438 0.292 ;
        RECT 0.938 0.248 1.006 0.382 ;
      LAYER m2 ;
        RECT 0.812 0.338 1.78 0.382 ;
      LAYER v1 ;
        RECT 0.942 0.338 1.002 0.382 ;
        RECT 1.698 0.338 1.758 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.694 0.473 1.762 0.517 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 5.2725 LAYER m1 ;
      ANTENNAMAXAREACAR 7.803611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 5.2725 LAYER m1 ;
      ANTENNAMAXAREACAR 7.803611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.202 ;
      LAYER m2 ;
        RECT 0.904 0.158 1.364 0.202 ;
      LAYER v1 ;
        RECT 0.942 0.158 1.002 0.202 ;
      LAYER v0 ;
        RECT 0.938 0.088 1.006 0.132 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    ANTENNADIFFAREA 0.02448 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.248 2.734 0.292 ;
        RECT 2.666 0.068 2.734 0.292 ;
        RECT 2.45 0.248 2.518 0.562 ;
        RECT 2.666 0.428 2.734 0.562 ;
      LAYER m2 ;
        RECT 2.524 0.158 3.076 0.202 ;
        RECT 2.432 0.518 3.076 0.562 ;
      LAYER v1 ;
        RECT 2.454 0.518 2.514 0.562 ;
        RECT 2.67 0.518 2.73 0.562 ;
        RECT 2.67 0.158 2.73 0.202 ;
      LAYER v0 ;
        RECT 2.666 0.473 2.734 0.517 ;
        RECT 2.666 0.138 2.734 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAGATEAREA 0.0045 LAYER m2 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
      ANTENNAMAXAREACAR 4.711111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.2515555 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0054 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 3.925926 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.248 2.194 0.292 ;
        RECT 1.91 0.158 1.978 0.292 ;
      LAYER m2 ;
        RECT 2 0.248 2.536 0.292 ;
      LAYER v1 ;
        RECT 2.022 0.248 2.082 0.292 ;
      LAYER v0 ;
        RECT 2.018 0.248 2.086 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0054 LAYER m2 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
      ANTENNAMAXAREACAR 3.20074075 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
      ANTENNAMAXAREACAR 2.4005555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.338 2.302 0.382 ;
      LAYER m2 ;
        RECT 2.108 0.338 2.752 0.382 ;
      LAYER v1 ;
        RECT 2.13 0.338 2.19 0.382 ;
      LAYER v0 ;
        RECT 2.126 0.338 2.194 0.382 ;
    END
  END rb
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.57 0.022 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.29 0.338 0.358 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.596 0.158 0.824 0.202 ;
        RECT 0.04 0.338 0.376 0.382 ;
      LAYER v1 ;
        RECT 0.078 0.338 0.138 0.382 ;
        RECT 0.294 0.338 0.354 0.382 ;
        RECT 0.618 0.158 0.678 0.202 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.363 0.142 0.407 ;
        RECT 0.182 0.498 0.25 0.542 ;
        RECT 0.182 0.363 0.25 0.407 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.363 0.358 0.407 ;
        RECT 0.614 0.223 0.682 0.267 ;
        RECT 0.614 0.088 0.682 0.132 ;
        RECT 0.722 0.223 0.79 0.267 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 0.83 0.223 0.898 0.267 ;
        RECT 0.83 0.088 0.898 0.132 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 2.018 0.1135 2.086 0.1575 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
    END
  END vssx
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.57 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
      LAYER v0 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.802 0.473 1.87 0.517 ;
        RECT 2.018 0.473 2.086 0.517 ;
        RECT 2.234 0.473 2.302 0.517 ;
        RECT 2.558 0.473 2.626 0.517 ;
        RECT 2.882 0.428 2.95 0.472 ;
    END
  END vcc
  OBS
    LAYER m2 ;
      RECT 1.568 0.428 2.444 0.472 ;
      RECT 1.784 0.158 2.444 0.202 ;
      RECT 3.188 0.338 3.508 0.382 ;
      RECT 3.712 0.248 4.048 0.292 ;
      RECT 4.036 0.518 4.496 0.562 ;
      RECT 4.036 0.158 4.496 0.202 ;
    LAYER m1 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.262 0.068 1.478 0.112 ;
      RECT 1.802 0.068 1.87 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.91 0.158 1.978 0.292 ;
      RECT 2.126 0.428 2.194 0.562 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.018 0.338 2.302 0.382 ;
      RECT 2.45 0.248 2.518 0.562 ;
      RECT 2.342 0.068 2.41 0.202 ;
      RECT 2.666 0.428 2.734 0.562 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.206 0.338 3.274 0.562 ;
      RECT 3.314 0.338 3.382 0.562 ;
      RECT 3.422 0.338 3.49 0.562 ;
      RECT 3.746 0.068 3.814 0.292 ;
      RECT 3.854 0.068 3.922 0.292 ;
      RECT 3.962 0.068 4.03 0.292 ;
      RECT 4.178 0.338 4.246 0.562 ;
      RECT 4.178 0.068 4.246 0.292 ;
      RECT 4.286 0.338 4.354 0.562 ;
      RECT 4.286 0.068 4.354 0.292 ;
      RECT 4.394 0.338 4.462 0.562 ;
      RECT 4.394 0.068 4.462 0.292 ;
    LAYER v1 ;
      RECT 4.398 0.158 4.458 0.202 ;
      RECT 4.398 0.518 4.458 0.562 ;
      RECT 4.182 0.158 4.242 0.202 ;
      RECT 4.182 0.518 4.242 0.562 ;
      RECT 3.966 0.248 4.026 0.292 ;
      RECT 3.75 0.248 3.81 0.292 ;
      RECT 3.426 0.338 3.486 0.382 ;
      RECT 3.21 0.338 3.27 0.382 ;
      RECT 2.346 0.158 2.406 0.202 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 1.59 0.428 1.65 0.472 ;
    LAYER v0 ;
      RECT 4.394 0.088 4.462 0.132 ;
      RECT 4.394 0.223 4.462 0.267 ;
      RECT 4.394 0.358 4.462 0.402 ;
      RECT 4.394 0.498 4.462 0.542 ;
      RECT 4.286 0.088 4.354 0.132 ;
      RECT 4.286 0.223 4.354 0.267 ;
      RECT 4.286 0.358 4.354 0.402 ;
      RECT 4.286 0.498 4.354 0.542 ;
      RECT 4.178 0.088 4.246 0.132 ;
      RECT 4.178 0.223 4.246 0.267 ;
      RECT 4.178 0.358 4.246 0.402 ;
      RECT 4.178 0.498 4.246 0.542 ;
      RECT 3.962 0.088 4.03 0.132 ;
      RECT 3.962 0.223 4.03 0.267 ;
      RECT 3.854 0.088 3.922 0.132 ;
      RECT 3.854 0.223 3.922 0.267 ;
      RECT 3.746 0.088 3.814 0.132 ;
      RECT 3.746 0.223 3.814 0.267 ;
      RECT 3.422 0.363 3.49 0.407 ;
      RECT 3.422 0.498 3.49 0.542 ;
      RECT 3.314 0.363 3.382 0.407 ;
      RECT 3.314 0.498 3.382 0.542 ;
      RECT 3.206 0.363 3.274 0.407 ;
      RECT 3.206 0.498 3.274 0.542 ;
      RECT 2.99 0.138 3.058 0.182 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.342 0.3445 2.41 0.3885 ;
      RECT 2.234 0.138 2.302 0.182 ;
      RECT 2.126 0.473 2.194 0.517 ;
      RECT 1.91 0.473 1.978 0.517 ;
      RECT 1.802 0.138 1.87 0.182 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.473 1.654 0.517 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.478 0.473 1.546 0.517 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.448 1.114 0.492 ;
    LAYER m1 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.338 1.438 0.382 ;
      RECT 1.006 0.248 1.438 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.87 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.978 0.248 2.194 0.292 ;
      RECT 2.302 0.248 2.342 0.292 ;
      RECT 2.342 0.248 2.41 0.472 ;
      RECT 2.518 0.248 2.666 0.292 ;
      RECT 2.666 0.068 2.734 0.292 ;
  END
END b15qbflf4gn1n08x5

MACRO b15qbfna2bn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qbfna2bn1n16x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAGATEAREA 0.0216 LAYER m2 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
      ANTENNAMAXAREACAR 1.39481475 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.26074075 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAGATEAREA 0.0288 LAYER m2 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
      ANTENNAMAXAREACAR 1.046111 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.1955555 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER m2 ;
        RECT 0.812 0.338 1.24 0.382 ;
      LAYER v1 ;
        RECT 1.158 0.338 1.218 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.2705 1.222 0.3145 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAGATEAREA 0.0216 LAYER m2 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59685175 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.39925925 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAGATEAREA 0.0288 LAYER m2 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
      ANTENNAMAXAREACAR 1.947639 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.2994445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.338 2.194 0.382 ;
        RECT 1.586 0.158 1.654 0.382 ;
      LAYER m2 ;
        RECT 1.46 0.248 1.888 0.292 ;
      LAYER v1 ;
        RECT 1.59 0.248 1.65 0.292 ;
      LAYER v0 ;
        RECT 1.802 0.338 1.87 0.382 ;
        RECT 2.018 0.338 2.086 0.382 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNADIFFAREA 0.07956 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0054 LAYER m2 ;
      ANTENNAMAXAREACAR 2.78666675 LAYER m1 ;
      ANTENNAMAXAREACAR 24.6014815 LAYER m2 ;
      ANTENNAMAXCUTCAR 3.4874075 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.428 2.214 0.472 ;
        RECT 1.046 0.158 1.114 0.472 ;
        RECT 1.262 0.338 1.546 0.382 ;
        RECT 1.478 0.158 1.546 0.382 ;
        RECT 1.262 0.158 1.33 0.382 ;
      LAYER m2 ;
        RECT 1.136 0.428 2.228 0.472 ;
        RECT 1.028 0.158 1.564 0.202 ;
      LAYER v1 ;
        RECT 1.05 0.158 1.11 0.202 ;
        RECT 1.158 0.428 1.218 0.472 ;
        RECT 1.266 0.158 1.326 0.202 ;
        RECT 1.374 0.428 1.434 0.472 ;
        RECT 1.482 0.158 1.542 0.202 ;
        RECT 1.59 0.428 1.65 0.472 ;
        RECT 1.914 0.428 1.974 0.472 ;
        RECT 2.13 0.428 2.19 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.262 0.178 1.33 0.222 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.478 0.178 1.546 0.222 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.126 0.428 2.194 0.472 ;
    END
  END o1
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.29 0.338 0.358 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.704 0.248 0.916 0.292 ;
        RECT 0.164 0.338 0.484 0.382 ;
      LAYER v1 ;
        RECT 0.186 0.338 0.246 0.382 ;
        RECT 0.726 0.248 0.786 0.292 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.363 0.142 0.407 ;
        RECT 0.182 0.498 0.25 0.542 ;
        RECT 0.182 0.363 0.25 0.407 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.363 0.358 0.407 ;
        RECT 0.614 0.223 0.682 0.267 ;
        RECT 0.614 0.088 0.682 0.132 ;
        RECT 0.722 0.223 0.79 0.267 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 0.83 0.223 0.898 0.267 ;
        RECT 0.83 0.088 0.898 0.132 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
    END
  END vssx
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
      LAYER v0 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.018 0.538 2.086 0.582 ;
    END
  END vcc
  OBS
    LAYER m2 ;
      RECT 2.308 0.428 2.536 0.472 ;
      RECT 2.324 0.158 2.536 0.202 ;
    LAYER m1 ;
      RECT 1.154 0.158 1.222 0.382 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 1.046 0.068 1.694 0.112 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.342 0.068 2.41 0.292 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 2.558 0.068 2.626 0.292 ;
    LAYER v1 ;
      RECT 2.454 0.158 2.514 0.202 ;
      RECT 2.454 0.428 2.514 0.472 ;
    LAYER v0 ;
      RECT 2.558 0.088 2.626 0.132 ;
      RECT 2.558 0.223 2.626 0.267 ;
      RECT 2.558 0.358 2.626 0.402 ;
      RECT 2.558 0.498 2.626 0.542 ;
      RECT 2.45 0.088 2.518 0.132 ;
      RECT 2.45 0.223 2.518 0.267 ;
      RECT 2.45 0.358 2.518 0.402 ;
      RECT 2.45 0.498 2.518 0.542 ;
      RECT 2.342 0.088 2.41 0.132 ;
      RECT 2.342 0.223 2.41 0.267 ;
      RECT 2.342 0.358 2.41 0.402 ;
      RECT 2.342 0.498 2.41 0.542 ;
      RECT 2.126 0.136 2.194 0.18 ;
      RECT 1.91 0.136 1.978 0.18 ;
      RECT 1.696 0.138 1.76 0.182 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.154 0.068 1.222 0.112 ;
    LAYER m1 ;
      RECT 1.262 0.158 1.33 0.382 ;
      RECT 1.33 0.338 1.478 0.382 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.654 0.338 2.194 0.382 ;
      RECT 1.694 0.068 1.762 0.292 ;
      RECT 1.762 0.248 1.91 0.292 ;
      RECT 1.91 0.068 1.978 0.292 ;
      RECT 1.978 0.248 2.126 0.292 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 1.114 0.428 2.214 0.472 ;
  END
END b15qbfna2bn1n16x5

MACRO b15qbfno2bn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qbfno2bn1n16x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAGATEAREA 0.0441 LAYER m2 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
      ANTENNAMAXAREACAR 1.04952375 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.18757375 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAGATEAREA 0.0297 LAYER m2 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
      ANTENNAMAXAREACAR 1.55838375 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.2785185 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.248 2.086 0.292 ;
        RECT 1.91 0.248 1.978 0.382 ;
        RECT 1.694 0.248 1.762 0.382 ;
      LAYER m2 ;
        RECT 1.46 0.338 1.996 0.382 ;
      LAYER v1 ;
        RECT 1.698 0.338 1.758 0.382 ;
        RECT 1.914 0.338 1.974 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.248 1.87 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAGATEAREA 0.0441 LAYER m2 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
      ANTENNAMAXAREACAR 0.84190475 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.1955555 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAGATEAREA 0.0297 LAYER m2 ;
      ANTENNAMAXAREACAR 0.63973075 LAYER m1 ;
      ANTENNAMAXAREACAR 1.250101 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.29037025 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.242 0.248 1.654 0.292 ;
      LAYER m2 ;
        RECT 1.012 0.248 1.472 0.292 ;
      LAYER v1 ;
        RECT 1.266 0.248 1.326 0.292 ;
      LAYER v0 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.478 0.248 1.546 0.292 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    ANTENNADIFFAREA 0.09792 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 2.302 0.202 ;
        RECT 1.046 0.158 1.114 0.562 ;
        RECT 1.694 0.518 2.302 0.562 ;
        RECT 2.234 0.338 2.302 0.562 ;
      LAYER m2 ;
        RECT 1.244 0.158 2.336 0.202 ;
        RECT 1.028 0.518 2.336 0.562 ;
      LAYER v1 ;
        RECT 1.05 0.518 1.11 0.562 ;
        RECT 1.266 0.158 1.326 0.202 ;
        RECT 1.482 0.158 1.542 0.202 ;
        RECT 1.698 0.158 1.758 0.202 ;
        RECT 1.806 0.518 1.866 0.562 ;
        RECT 1.914 0.158 1.974 0.202 ;
        RECT 2.022 0.518 2.082 0.562 ;
        RECT 2.13 0.158 2.19 0.202 ;
        RECT 2.238 0.518 2.298 0.562 ;
      LAYER v0 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.802 0.518 1.87 0.562 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.018 0.518 2.086 0.562 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.234 0.428 2.302 0.472 ;
    END
  END o1
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.29 0.338 0.358 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.596 0.248 0.932 0.292 ;
        RECT 0.164 0.338 0.376 0.382 ;
      LAYER v1 ;
        RECT 0.186 0.338 0.246 0.382 ;
        RECT 0.726 0.248 0.786 0.292 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.363 0.142 0.407 ;
        RECT 0.182 0.498 0.25 0.542 ;
        RECT 0.182 0.363 0.25 0.407 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.363 0.358 0.407 ;
        RECT 0.614 0.223 0.682 0.267 ;
        RECT 0.614 0.088 0.682 0.132 ;
        RECT 0.722 0.223 0.79 0.267 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 0.83 0.223 0.898 0.267 ;
        RECT 0.83 0.088 0.898 0.132 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
    END
  END vssx
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
      LAYER v0 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  OBS
    LAYER m2 ;
      RECT 2.416 0.518 2.644 0.562 ;
      RECT 2.416 0.158 2.644 0.202 ;
    LAYER m1 ;
      RECT 1.242 0.248 1.654 0.292 ;
      RECT 1.154 0.428 2.126 0.472 ;
      RECT 1.694 0.518 2.234 0.562 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 2.558 0.068 2.626 0.292 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.666 0.068 2.734 0.292 ;
    LAYER v1 ;
      RECT 2.562 0.158 2.622 0.202 ;
      RECT 2.562 0.518 2.622 0.562 ;
    LAYER v0 ;
      RECT 2.666 0.088 2.734 0.132 ;
      RECT 2.666 0.223 2.734 0.267 ;
      RECT 2.666 0.358 2.734 0.402 ;
      RECT 2.666 0.498 2.734 0.542 ;
      RECT 2.558 0.088 2.626 0.132 ;
      RECT 2.558 0.223 2.626 0.267 ;
      RECT 2.558 0.358 2.626 0.402 ;
      RECT 2.558 0.498 2.626 0.542 ;
      RECT 2.45 0.088 2.518 0.132 ;
      RECT 2.45 0.223 2.518 0.267 ;
      RECT 2.45 0.358 2.518 0.402 ;
      RECT 2.45 0.498 2.518 0.542 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.428 1.33 0.472 ;
    LAYER m1 ;
      RECT 1.694 0.248 1.762 0.382 ;
      RECT 1.762 0.248 1.91 0.292 ;
      RECT 1.91 0.248 1.978 0.382 ;
      RECT 1.978 0.248 2.086 0.292 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 1.114 0.158 2.302 0.202 ;
  END
END b15qbfno2bn1n16x5

MACRO b15qbnbf1bn1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qbnbf1bn1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.428 0.5 0.472 ;
      RECT 0.04 0.338 0.932 0.382 ;
      RECT 0.58 0.428 1.564 0.472 ;
      RECT 0.488 0.158 1.564 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.506 0.428 1.006 0.472 ;
      RECT 0.614 0.338 1.154 0.382 ;
      RECT 0.614 0.248 1.046 0.292 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.586 0.068 1.654 0.292 ;
    LAYER v1 ;
      RECT 1.482 0.158 1.542 0.202 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 0.834 0.158 0.894 0.202 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.618 0.158 0.678 0.202 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.402 0.428 0.462 0.472 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.223 1.654 0.267 ;
      RECT 1.586 0.358 1.654 0.402 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.478 0.088 1.546 0.132 ;
      RECT 1.478 0.223 1.546 0.267 ;
      RECT 1.478 0.358 1.546 0.402 ;
      RECT 1.478 0.498 1.546 0.542 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.223 1.438 0.267 ;
      RECT 1.37 0.358 1.438 0.402 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.29 0.363 0.358 0.407 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.363 0.25 0.407 ;
      RECT 0.182 0.498 0.25 0.542 ;
      RECT 0.074 0.363 0.142 0.407 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.158 1.006 0.202 ;
      RECT 1.154 0.158 1.222 0.382 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.046 0.518 1.262 0.562 ;
      RECT 1.114 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.562 ;
  END
END b15qbnbf1bn1n16x5

MACRO b15qbnbf1bn1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qbnbf1bn1n32x5 0 0 ;
  SIZE 2.376 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.41 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 1.046 0.538 1.114 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.41 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 0.592 0.382 ;
      RECT 0.812 0.428 1.04 0.472 ;
      RECT 1.12 0.428 2.212 0.472 ;
      RECT 1.136 0.158 2.212 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.046 0.428 1.978 0.472 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 2.234 0.068 2.302 0.292 ;
    LAYER v1 ;
      RECT 2.13 0.158 2.19 0.202 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.59 0.158 1.65 0.202 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.374 0.158 1.434 0.202 ;
      RECT 1.374 0.428 1.434 0.472 ;
      RECT 1.158 0.158 1.218 0.202 ;
      RECT 1.158 0.428 1.218 0.472 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 2.234 0.088 2.302 0.132 ;
      RECT 2.234 0.223 2.302 0.267 ;
      RECT 2.234 0.358 2.302 0.402 ;
      RECT 2.234 0.498 2.302 0.542 ;
      RECT 2.126 0.088 2.194 0.132 ;
      RECT 2.126 0.223 2.194 0.267 ;
      RECT 2.126 0.358 2.194 0.402 ;
      RECT 2.126 0.498 2.194 0.542 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 2.018 0.223 2.086 0.267 ;
      RECT 2.018 0.358 2.086 0.402 ;
      RECT 2.018 0.498 2.086 0.542 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.616 0.4385 0.68 0.4825 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.363 0.358 0.407 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.363 0.25 0.407 ;
      RECT 0.182 0.498 0.25 0.542 ;
      RECT 0.074 0.363 0.142 0.407 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 1.006 0.158 1.978 0.202 ;
  END
END b15qbnbf1bn1n32x5

MACRO b15qbnff4gn1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qbnff4gn1n08x5 0 0 ;
  SIZE 7.452 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 7.486 0.652 ;
        RECT 6.878 0.428 6.946 0.652 ;
        RECT 6.662 0.518 6.73 0.652 ;
        RECT 6.446 0.338 6.514 0.652 ;
        RECT 5.15 0.428 5.218 0.652 ;
        RECT 4.934 0.428 5.002 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.206 0.338 3.274 0.652 ;
        RECT 2.99 0.338 3.058 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.262 0.338 1.33 0.652 ;
      LAYER v0 ;
        RECT 1.262 0.408 1.33 0.452 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.99 0.3835 3.058 0.4275 ;
        RECT 3.208 0.428 3.272 0.472 ;
        RECT 3.962 0.538 4.03 0.582 ;
        RECT 4.61 0.448 4.678 0.492 ;
        RECT 4.934 0.448 5.002 0.492 ;
        RECT 5.15 0.448 5.218 0.492 ;
        RECT 6.446 0.428 6.514 0.472 ;
        RECT 6.664 0.538 6.728 0.582 ;
        RECT 6.878 0.448 6.946 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 7.486 0.022 ;
        RECT 6.878 -0.022 6.946 0.112 ;
        RECT 6.662 -0.022 6.73 0.112 ;
        RECT 6.446 -0.022 6.514 0.202 ;
        RECT 5.15 -0.022 5.218 0.202 ;
        RECT 4.718 -0.022 4.786 0.292 ;
        RECT 2.558 0.158 3.726 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.262 -0.022 1.33 0.292 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.262 0.203 1.33 0.247 ;
        RECT 1.91 0.048 1.978 0.092 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.206 0.158 3.274 0.202 ;
        RECT 3.422 0.158 3.49 0.202 ;
        RECT 3.638 0.158 3.706 0.202 ;
        RECT 4.718 0.203 4.786 0.247 ;
        RECT 5.15 0.138 5.218 0.182 ;
        RECT 6.446 0.138 6.514 0.182 ;
        RECT 6.664 0.048 6.728 0.092 ;
        RECT 6.88 0.048 6.944 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.596 0.158 1.456 0.202 ;
      RECT 0.164 0.428 1.58 0.472 ;
      RECT 1.028 0.338 2.12 0.382 ;
      RECT 1.352 0.518 2.32 0.562 ;
      RECT 2.2 0.338 3.616 0.382 ;
      RECT 1.66 0.428 4.28 0.472 ;
      RECT 2.756 0.518 5.128 0.562 ;
      RECT 4.808 0.068 5.668 0.112 ;
      RECT 4.16 0.338 6.1 0.382 ;
      RECT 6.428 0.518 6.656 0.562 ;
      RECT 4.36 0.428 6.748 0.472 ;
      RECT 6.736 0.518 7.288 0.562 ;
      RECT 6.536 0.158 7.288 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.91 0.248 1.978 0.382 ;
      RECT 2.234 0.158 2.302 0.472 ;
      RECT 2.342 0.248 2.41 0.472 ;
      RECT 2.234 0.518 2.43 0.562 ;
      RECT 2.558 0.248 2.626 0.472 ;
      RECT 2.666 0.518 2.95 0.562 ;
      RECT 3.422 0.338 3.834 0.382 ;
      RECT 3.942 0.338 4.246 0.382 ;
      RECT 4.07 0.428 4.286 0.472 ;
      RECT 4.178 0.158 4.394 0.202 ;
      RECT 2.774 0.068 4.502 0.112 ;
      RECT 4.826 0.248 4.894 0.562 ;
      RECT 4.61 0.068 4.678 0.382 ;
      RECT 4.718 0.428 4.786 0.562 ;
      RECT 6.554 0.158 6.622 0.562 ;
      RECT 5.042 0.068 5.11 0.562 ;
      RECT 5.366 0.068 5.434 0.292 ;
      RECT 5.474 0.068 5.542 0.292 ;
      RECT 5.582 0.068 5.65 0.292 ;
      RECT 5.906 0.338 5.974 0.562 ;
      RECT 6.014 0.338 6.082 0.562 ;
      RECT 6.122 0.338 6.19 0.562 ;
      RECT 6.338 0.068 6.406 0.562 ;
      RECT 6.662 0.248 6.73 0.472 ;
      RECT 6.77 0.338 6.838 0.562 ;
      RECT 7.094 0.338 7.162 0.562 ;
      RECT 7.094 0.068 7.162 0.292 ;
      RECT 7.202 0.338 7.27 0.562 ;
      RECT 7.202 0.068 7.27 0.292 ;
      RECT 7.31 0.338 7.378 0.562 ;
      RECT 7.31 0.068 7.378 0.292 ;
    LAYER v1 ;
      RECT 7.206 0.158 7.266 0.202 ;
      RECT 7.206 0.518 7.266 0.562 ;
      RECT 6.774 0.158 6.834 0.202 ;
      RECT 6.774 0.518 6.834 0.562 ;
      RECT 6.666 0.428 6.726 0.472 ;
      RECT 6.558 0.518 6.618 0.562 ;
      RECT 6.018 0.338 6.078 0.382 ;
      RECT 5.478 0.068 5.538 0.112 ;
      RECT 5.046 0.068 5.106 0.112 ;
      RECT 5.046 0.518 5.106 0.562 ;
      RECT 4.722 0.428 4.782 0.472 ;
      RECT 4.614 0.338 4.674 0.382 ;
      RECT 4.398 0.428 4.458 0.472 ;
      RECT 4.182 0.338 4.242 0.382 ;
      RECT 4.182 0.428 4.242 0.472 ;
      RECT 3.534 0.338 3.594 0.382 ;
      RECT 2.778 0.518 2.838 0.562 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 2.238 0.518 2.298 0.562 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 1.158 0.158 1.218 0.202 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.726 0.158 0.786 0.202 ;
      RECT 0.186 0.428 0.246 0.472 ;
    LAYER v0 ;
      RECT 7.31 0.088 7.378 0.132 ;
      RECT 7.31 0.223 7.378 0.267 ;
      RECT 7.31 0.358 7.378 0.402 ;
      RECT 7.31 0.498 7.378 0.542 ;
      RECT 7.202 0.088 7.27 0.132 ;
      RECT 7.202 0.223 7.27 0.267 ;
      RECT 7.202 0.358 7.27 0.402 ;
      RECT 7.202 0.498 7.27 0.542 ;
      RECT 7.094 0.088 7.162 0.132 ;
      RECT 7.094 0.223 7.162 0.267 ;
      RECT 7.094 0.358 7.162 0.402 ;
      RECT 7.094 0.498 7.162 0.542 ;
      RECT 6.77 0.158 6.838 0.202 ;
      RECT 6.77 0.448 6.838 0.492 ;
      RECT 6.662 0.338 6.73 0.382 ;
      RECT 6.338 0.138 6.406 0.182 ;
      RECT 6.338 0.428 6.406 0.472 ;
      RECT 6.122 0.363 6.19 0.407 ;
      RECT 6.122 0.498 6.19 0.542 ;
      RECT 6.014 0.363 6.082 0.407 ;
      RECT 6.014 0.498 6.082 0.542 ;
      RECT 5.906 0.363 5.974 0.407 ;
      RECT 5.906 0.498 5.974 0.542 ;
      RECT 5.582 0.088 5.65 0.132 ;
      RECT 5.582 0.223 5.65 0.267 ;
      RECT 5.474 0.088 5.542 0.132 ;
      RECT 5.474 0.223 5.542 0.267 ;
      RECT 5.366 0.088 5.434 0.132 ;
      RECT 5.366 0.223 5.434 0.267 ;
      RECT 5.042 0.248 5.11 0.292 ;
      RECT 4.934 0.138 5.002 0.182 ;
      RECT 4.826 0.448 4.894 0.492 ;
      RECT 4.718 0.448 4.786 0.492 ;
      RECT 4.61 0.088 4.678 0.132 ;
      RECT 4.502 0.338 4.57 0.382 ;
      RECT 4.394 0.068 4.462 0.112 ;
      RECT 4.394 0.428 4.462 0.472 ;
      RECT 4.286 0.158 4.354 0.202 ;
      RECT 4.286 0.338 4.354 0.382 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 4.07 0.338 4.138 0.382 ;
      RECT 3.854 0.248 3.922 0.292 ;
      RECT 3.854 0.428 3.922 0.472 ;
      RECT 3.746 0.338 3.814 0.382 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.774 0.518 2.842 0.562 ;
      RECT 2.558 0.293 2.626 0.337 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.342 0.518 2.41 0.562 ;
      RECT 2.234 0.3835 2.302 0.4275 ;
      RECT 2.128 0.088 2.192 0.132 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.478 0.498 1.546 0.542 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.37 0.408 1.438 0.452 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.203 1.114 0.247 ;
      RECT 1.046 0.4055 1.114 0.4495 ;
      RECT 0.83 0.088 0.898 0.132 ;
      RECT 0.83 0.223 0.898 0.267 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.223 0.79 0.267 ;
      RECT 0.614 0.088 0.682 0.132 ;
      RECT 0.614 0.223 0.682 0.267 ;
      RECT 0.29 0.363 0.358 0.407 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.363 0.25 0.407 ;
      RECT 0.182 0.498 0.25 0.542 ;
      RECT 0.074 0.363 0.142 0.407 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.438 0.068 1.694 0.112 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.762 0.158 2.126 0.202 ;
      RECT 2.126 0.068 2.194 0.202 ;
      RECT 2.302 0.158 2.518 0.202 ;
      RECT 2.626 0.428 2.882 0.472 ;
      RECT 2.882 0.248 2.95 0.472 ;
      RECT 2.95 0.248 3.314 0.292 ;
      RECT 3.314 0.248 3.382 0.472 ;
      RECT 3.382 0.428 4.03 0.472 ;
      RECT 3.382 0.248 4.246 0.292 ;
      RECT 4.286 0.248 4.354 0.472 ;
      RECT 4.394 0.158 4.462 0.562 ;
      RECT 4.502 0.068 4.57 0.472 ;
      RECT 4.894 0.248 4.934 0.292 ;
      RECT 4.934 0.068 5.002 0.292 ;
      RECT 6.622 0.158 6.946 0.202 ;
  END
END b15qbnff4gn1n08x5

MACRO b15qbnin1bn1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qbnin1bn1n16x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.938 0.538 1.006 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.518 0.5 0.562 ;
      RECT 0.04 0.428 0.916 0.472 ;
      RECT 0.58 0.518 1.472 0.562 ;
      RECT 0.488 0.158 1.472 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.262 0.068 1.33 0.292 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.292 ;
    LAYER v1 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.266 0.518 1.326 0.562 ;
      RECT 0.834 0.158 0.894 0.202 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.618 0.158 0.678 0.202 ;
      RECT 0.618 0.518 0.678 0.562 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.402 0.518 0.462 0.562 ;
      RECT 0.186 0.428 0.246 0.472 ;
    LAYER v0 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.223 1.438 0.267 ;
      RECT 1.37 0.358 1.438 0.402 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.262 0.088 1.33 0.132 ;
      RECT 1.262 0.223 1.33 0.267 ;
      RECT 1.262 0.358 1.33 0.402 ;
      RECT 1.262 0.498 1.33 0.542 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.223 1.222 0.267 ;
      RECT 1.154 0.358 1.222 0.402 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.363 0.358 0.407 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.363 0.25 0.407 ;
      RECT 0.182 0.498 0.25 0.542 ;
      RECT 0.074 0.363 0.142 0.407 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.466 0.158 1.006 0.202 ;
  END
END b15qbnin1bn1n16x5

MACRO b15qbnin1bn1n40x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qbnin1bn1n40x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 1.04 0.382 ;
      RECT 0.04 0.248 1.672 0.292 ;
      RECT 0.596 0.158 1.996 0.202 ;
      RECT 1.12 0.338 2.12 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.182 0.248 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 1.046 0.248 1.674 0.292 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.91 0.068 1.978 0.292 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.018 0.068 2.086 0.292 ;
    LAYER v1 ;
      RECT 1.914 0.158 1.974 0.202 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.59 0.248 1.65 0.292 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.482 0.158 1.542 0.202 ;
      RECT 1.374 0.248 1.434 0.292 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.158 0.248 1.218 0.292 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 1.05 0.158 1.11 0.202 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.158 0.894 0.202 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.618 0.158 0.678 0.202 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.248 0.246 0.292 ;
    LAYER v0 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 2.018 0.223 2.086 0.267 ;
      RECT 2.018 0.358 2.086 0.402 ;
      RECT 2.018 0.498 2.086 0.542 ;
      RECT 1.91 0.088 1.978 0.132 ;
      RECT 1.91 0.223 1.978 0.267 ;
      RECT 1.91 0.358 1.978 0.402 ;
      RECT 1.91 0.498 1.978 0.542 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.223 1.87 0.267 ;
      RECT 1.802 0.358 1.87 0.402 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.29 0.363 0.358 0.407 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.363 0.25 0.407 ;
      RECT 0.182 0.498 0.25 0.542 ;
      RECT 0.074 0.363 0.142 0.407 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 0.506 0.428 1.154 0.472 ;
      RECT 1.154 0.338 1.222 0.472 ;
      RECT 1.222 0.428 1.37 0.472 ;
      RECT 1.37 0.338 1.438 0.472 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.338 1.654 0.472 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 0.79 0.158 0.938 0.202 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.006 0.158 1.654 0.202 ;
  END
END b15qbnin1bn1n40x5

MACRO b15qbnlf4gn1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qbnlf4gn1n08x5 0 0 ;
  SIZE 4.536 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.57 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
      LAYER v0 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.802 0.473 1.87 0.517 ;
        RECT 2.018 0.473 2.086 0.517 ;
        RECT 2.234 0.473 2.302 0.517 ;
        RECT 2.558 0.473 2.626 0.517 ;
        RECT 2.882 0.428 2.95 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.57 0.022 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 2.018 0.1135 2.086 0.1575 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.596 0.158 1.348 0.202 ;
      RECT 0.04 0.338 1.78 0.382 ;
      RECT 1.568 0.428 2.428 0.472 ;
      RECT 1.784 0.158 2.444 0.202 ;
      RECT 2.324 0.518 2.552 0.562 ;
      RECT 2.108 0.338 3.508 0.382 ;
      RECT 2 0.248 4.048 0.292 ;
      RECT 2.632 0.518 4.496 0.562 ;
      RECT 2.524 0.158 4.496 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.262 0.068 1.478 0.112 ;
      RECT 1.802 0.068 1.87 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.91 0.158 1.978 0.292 ;
      RECT 2.126 0.428 2.194 0.562 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.018 0.338 2.302 0.382 ;
      RECT 2.45 0.248 2.518 0.562 ;
      RECT 2.342 0.068 2.41 0.202 ;
      RECT 2.666 0.428 2.734 0.562 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.206 0.338 3.274 0.562 ;
      RECT 3.314 0.338 3.382 0.562 ;
      RECT 3.422 0.338 3.49 0.562 ;
      RECT 3.746 0.068 3.814 0.292 ;
      RECT 3.854 0.068 3.922 0.292 ;
      RECT 3.962 0.068 4.03 0.292 ;
      RECT 4.178 0.338 4.246 0.562 ;
      RECT 4.178 0.068 4.246 0.292 ;
      RECT 4.286 0.338 4.354 0.562 ;
      RECT 4.286 0.068 4.354 0.292 ;
      RECT 4.394 0.338 4.462 0.562 ;
      RECT 4.394 0.068 4.462 0.292 ;
    LAYER v1 ;
      RECT 4.398 0.158 4.458 0.202 ;
      RECT 4.398 0.518 4.458 0.562 ;
      RECT 4.182 0.158 4.242 0.202 ;
      RECT 4.182 0.518 4.242 0.562 ;
      RECT 3.966 0.248 4.026 0.292 ;
      RECT 3.75 0.248 3.81 0.292 ;
      RECT 3.426 0.338 3.486 0.382 ;
      RECT 3.21 0.338 3.27 0.382 ;
      RECT 2.67 0.158 2.73 0.202 ;
      RECT 2.67 0.518 2.73 0.562 ;
      RECT 2.454 0.518 2.514 0.562 ;
      RECT 2.346 0.158 2.406 0.202 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.13 0.338 2.19 0.382 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 2.022 0.248 2.082 0.292 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 0.942 0.158 1.002 0.202 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.618 0.158 0.678 0.202 ;
      RECT 0.294 0.338 0.354 0.382 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 4.394 0.088 4.462 0.132 ;
      RECT 4.394 0.223 4.462 0.267 ;
      RECT 4.394 0.358 4.462 0.402 ;
      RECT 4.394 0.498 4.462 0.542 ;
      RECT 4.286 0.088 4.354 0.132 ;
      RECT 4.286 0.223 4.354 0.267 ;
      RECT 4.286 0.358 4.354 0.402 ;
      RECT 4.286 0.498 4.354 0.542 ;
      RECT 4.178 0.088 4.246 0.132 ;
      RECT 4.178 0.223 4.246 0.267 ;
      RECT 4.178 0.358 4.246 0.402 ;
      RECT 4.178 0.498 4.246 0.542 ;
      RECT 3.962 0.088 4.03 0.132 ;
      RECT 3.962 0.223 4.03 0.267 ;
      RECT 3.854 0.088 3.922 0.132 ;
      RECT 3.854 0.223 3.922 0.267 ;
      RECT 3.746 0.088 3.814 0.132 ;
      RECT 3.746 0.223 3.814 0.267 ;
      RECT 3.422 0.363 3.49 0.407 ;
      RECT 3.422 0.498 3.49 0.542 ;
      RECT 3.314 0.363 3.382 0.407 ;
      RECT 3.314 0.498 3.382 0.542 ;
      RECT 3.206 0.363 3.274 0.407 ;
      RECT 3.206 0.498 3.274 0.542 ;
      RECT 2.99 0.138 3.058 0.182 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.666 0.138 2.734 0.182 ;
      RECT 2.666 0.473 2.734 0.517 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.342 0.3445 2.41 0.3885 ;
      RECT 2.234 0.138 2.302 0.182 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.126 0.473 2.194 0.517 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.91 0.473 1.978 0.517 ;
      RECT 1.802 0.138 1.87 0.182 ;
      RECT 1.694 0.473 1.762 0.517 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.473 1.654 0.517 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.478 0.473 1.546 0.517 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.83 0.088 0.898 0.132 ;
      RECT 0.83 0.223 0.898 0.267 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.223 0.79 0.267 ;
      RECT 0.614 0.088 0.682 0.132 ;
      RECT 0.614 0.223 0.682 0.267 ;
      RECT 0.29 0.363 0.358 0.407 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.363 0.25 0.407 ;
      RECT 0.182 0.498 0.25 0.542 ;
      RECT 0.074 0.363 0.142 0.407 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.338 1.438 0.382 ;
      RECT 1.006 0.248 1.438 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.87 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.978 0.248 2.194 0.292 ;
      RECT 2.302 0.248 2.342 0.292 ;
      RECT 2.342 0.248 2.41 0.472 ;
      RECT 2.518 0.248 2.666 0.292 ;
      RECT 2.666 0.068 2.734 0.292 ;
  END
END b15qbnlf4gn1n08x5

MACRO b15qbnna2bn1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qbnna2bn1n16x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
      LAYER v0 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.018 0.538 2.086 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.158 1.148 0.202 ;
      RECT 0.164 0.338 1.24 0.382 ;
      RECT 0.704 0.248 1.888 0.292 ;
      RECT 1.136 0.428 2.536 0.472 ;
      RECT 1.228 0.158 2.536 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 1.154 0.158 1.222 0.382 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 1.046 0.068 1.694 0.112 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.342 0.068 2.41 0.292 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 2.558 0.068 2.626 0.292 ;
    LAYER v1 ;
      RECT 2.454 0.158 2.514 0.202 ;
      RECT 2.454 0.428 2.514 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.59 0.248 1.65 0.292 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.482 0.158 1.542 0.202 ;
      RECT 1.374 0.428 1.434 0.472 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 1.158 0.428 1.218 0.472 ;
      RECT 1.05 0.158 1.11 0.202 ;
      RECT 0.726 0.248 0.786 0.292 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 2.558 0.088 2.626 0.132 ;
      RECT 2.558 0.223 2.626 0.267 ;
      RECT 2.558 0.358 2.626 0.402 ;
      RECT 2.558 0.498 2.626 0.542 ;
      RECT 2.45 0.088 2.518 0.132 ;
      RECT 2.45 0.223 2.518 0.267 ;
      RECT 2.45 0.358 2.518 0.402 ;
      RECT 2.45 0.498 2.518 0.542 ;
      RECT 2.342 0.088 2.41 0.132 ;
      RECT 2.342 0.223 2.41 0.267 ;
      RECT 2.342 0.358 2.41 0.402 ;
      RECT 2.342 0.498 2.41 0.542 ;
      RECT 2.126 0.136 2.194 0.18 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.136 1.978 0.18 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.696 0.138 1.76 0.182 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.2705 1.222 0.3145 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.83 0.088 0.898 0.132 ;
      RECT 0.83 0.223 0.898 0.267 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.223 0.79 0.267 ;
      RECT 0.614 0.088 0.682 0.132 ;
      RECT 0.614 0.223 0.682 0.267 ;
      RECT 0.29 0.363 0.358 0.407 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.363 0.25 0.407 ;
      RECT 0.182 0.498 0.25 0.542 ;
      RECT 0.074 0.363 0.142 0.407 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 1.262 0.158 1.33 0.382 ;
      RECT 1.33 0.338 1.478 0.382 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.654 0.338 2.194 0.382 ;
      RECT 1.694 0.068 1.762 0.292 ;
      RECT 1.762 0.248 1.91 0.292 ;
      RECT 1.91 0.068 1.978 0.292 ;
      RECT 1.978 0.248 2.126 0.292 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 1.114 0.428 2.214 0.472 ;
  END
END b15qbnna2bn1n16x5

MACRO b15qbnno2bn1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qbnno2bn1n16x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
      LAYER v0 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.028 0.518 1.256 0.562 ;
      RECT 0.596 0.248 1.456 0.292 ;
      RECT 0.164 0.338 1.996 0.382 ;
      RECT 1.336 0.518 2.644 0.562 ;
      RECT 1.244 0.158 2.644 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 1.242 0.248 1.654 0.292 ;
      RECT 1.154 0.428 2.126 0.472 ;
      RECT 1.694 0.518 2.234 0.562 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 2.558 0.068 2.626 0.292 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.666 0.068 2.734 0.292 ;
    LAYER v1 ;
      RECT 2.562 0.158 2.622 0.202 ;
      RECT 2.562 0.518 2.622 0.562 ;
      RECT 2.238 0.518 2.298 0.562 ;
      RECT 2.13 0.158 2.19 0.202 ;
      RECT 2.022 0.518 2.082 0.562 ;
      RECT 1.914 0.158 1.974 0.202 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.698 0.158 1.758 0.202 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.482 0.158 1.542 0.202 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.266 0.248 1.326 0.292 ;
      RECT 1.05 0.518 1.11 0.562 ;
      RECT 0.726 0.248 0.786 0.292 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 2.666 0.088 2.734 0.132 ;
      RECT 2.666 0.223 2.734 0.267 ;
      RECT 2.666 0.358 2.734 0.402 ;
      RECT 2.666 0.498 2.734 0.542 ;
      RECT 2.558 0.088 2.626 0.132 ;
      RECT 2.558 0.223 2.626 0.267 ;
      RECT 2.558 0.358 2.626 0.402 ;
      RECT 2.558 0.498 2.626 0.542 ;
      RECT 2.45 0.088 2.518 0.132 ;
      RECT 2.45 0.223 2.518 0.267 ;
      RECT 2.45 0.358 2.518 0.402 ;
      RECT 2.45 0.498 2.518 0.542 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 0.83 0.088 0.898 0.132 ;
      RECT 0.83 0.223 0.898 0.267 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.223 0.79 0.267 ;
      RECT 0.614 0.088 0.682 0.132 ;
      RECT 0.614 0.223 0.682 0.267 ;
      RECT 0.29 0.363 0.358 0.407 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.363 0.25 0.407 ;
      RECT 0.182 0.498 0.25 0.542 ;
      RECT 0.074 0.363 0.142 0.407 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 1.694 0.248 1.762 0.382 ;
      RECT 1.762 0.248 1.91 0.292 ;
      RECT 1.91 0.248 1.978 0.382 ;
      RECT 1.978 0.248 2.086 0.292 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 1.114 0.158 2.302 0.202 ;
  END
END b15qbnno2bn1n16x5

MACRO b15qfd1x2an1nnpx5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qfd1x2an1nnpx5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.182 0.338 0.898 0.382 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.506 0.338 0.574 0.562 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.182 0.338 0.25 0.562 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.518 0.142 0.562 ;
        RECT 0.184 0.4125 0.248 0.4565 ;
        RECT 0.29 0.518 0.358 0.562 ;
        RECT 0.508 0.4125 0.572 0.4565 ;
        RECT 0.614 0.518 0.682 0.562 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.182 0.248 0.898 0.292 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.506 0.068 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.182 0.068 0.25 0.292 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.184 0.1755 0.248 0.2195 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.508 0.1755 0.572 0.2195 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.046 0.068 1.114 0.112 ;
        RECT 1.262 0.068 1.33 0.112 ;
        RECT 1.478 0.068 1.546 0.112 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.154 0.068 1.222 0.202 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.202 ;
  END
END b15qfd1x2an1nnpx5

MACRO b15qfdglban1v00x5
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN b15qfdglban1v00x5 0 0 ;
  SIZE 9.504 BY 10.08 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 9.538 0.652 ;
        RECT 7.958 0.608 8.026 0.742 ;
        RECT 1.478 0.608 1.546 0.742 ;
        RECT -0.034 1.868 9.538 1.912 ;
        RECT 7.526 1.778 7.594 1.912 ;
        RECT 7.094 1.868 7.162 2.002 ;
        RECT 2.342 1.868 2.41 2.002 ;
        RECT 1.91 1.778 1.978 1.912 ;
        RECT -0.034 3.128 9.538 3.172 ;
        RECT 6.662 3.038 6.73 3.172 ;
        RECT 6.23 3.128 6.298 3.262 ;
        RECT 3.206 3.128 3.274 3.262 ;
        RECT 2.774 3.038 2.842 3.172 ;
        RECT -0.034 4.388 9.538 4.432 ;
        RECT 5.798 4.298 5.866 4.432 ;
        RECT 5.366 4.388 5.434 4.612 ;
        RECT 5.15 4.388 5.218 4.612 ;
        RECT 4.934 4.388 5.002 4.612 ;
        RECT 4.07 4.658 4.786 4.702 ;
        RECT 4.718 4.388 4.786 4.702 ;
        RECT 4.502 4.388 4.57 4.612 ;
        RECT 4.394 4.478 4.462 4.702 ;
        RECT 4.178 4.388 4.246 4.612 ;
        RECT 4.07 4.478 4.138 4.702 ;
        RECT 3.962 4.388 4.03 4.612 ;
        RECT 3.638 4.298 3.706 4.432 ;
        RECT -0.034 5.648 9.538 5.692 ;
        RECT 5.798 5.648 5.866 5.782 ;
        RECT 5.366 5.468 5.434 5.692 ;
        RECT 5.15 5.468 5.218 5.692 ;
        RECT 4.934 5.468 5.002 5.692 ;
        RECT 4.718 5.378 4.786 5.692 ;
        RECT 4.07 5.378 4.786 5.422 ;
        RECT 4.502 5.468 4.57 5.692 ;
        RECT 4.394 5.378 4.462 5.602 ;
        RECT 4.178 5.468 4.246 5.692 ;
        RECT 4.07 5.378 4.138 5.602 ;
        RECT 3.962 5.468 4.03 5.692 ;
        RECT 3.638 5.648 3.706 5.782 ;
        RECT -0.034 6.908 9.538 6.952 ;
        RECT 6.662 6.908 6.73 7.042 ;
        RECT 6.23 6.818 6.298 6.952 ;
        RECT 3.206 6.818 3.274 6.952 ;
        RECT 2.774 6.908 2.842 7.042 ;
        RECT -0.034 8.168 9.538 8.212 ;
        RECT 7.526 8.168 7.594 8.302 ;
        RECT 7.094 8.078 7.162 8.212 ;
        RECT 2.342 8.078 2.41 8.212 ;
        RECT 1.91 8.168 1.978 8.302 ;
        RECT -0.034 9.428 9.538 9.472 ;
        RECT 7.958 9.338 8.026 9.472 ;
        RECT 1.478 9.338 1.546 9.472 ;
      LAYER v0 ;
        RECT 1.48 9.358 1.544 9.402 ;
        RECT 1.48 0.678 1.544 0.722 ;
        RECT 1.912 8.238 1.976 8.282 ;
        RECT 1.912 1.798 1.976 1.842 ;
        RECT 2.344 8.098 2.408 8.142 ;
        RECT 2.344 1.938 2.408 1.982 ;
        RECT 2.776 6.978 2.84 7.022 ;
        RECT 2.776 3.058 2.84 3.102 ;
        RECT 3.208 6.838 3.272 6.882 ;
        RECT 3.208 3.198 3.272 3.242 ;
        RECT 3.64 5.718 3.704 5.762 ;
        RECT 3.64 4.318 3.704 4.362 ;
        RECT 3.962 5.558 4.03 5.602 ;
        RECT 3.962 4.478 4.03 4.522 ;
        RECT 4.072 5.4525 4.136 5.4965 ;
        RECT 4.072 4.5835 4.136 4.6275 ;
        RECT 4.178 5.558 4.246 5.602 ;
        RECT 4.178 4.478 4.246 4.522 ;
        RECT 4.396 5.4525 4.46 5.4965 ;
        RECT 4.396 4.5835 4.46 4.6275 ;
        RECT 4.502 5.558 4.57 5.602 ;
        RECT 4.502 4.478 4.57 4.522 ;
        RECT 4.936 5.578 5 5.622 ;
        RECT 4.936 4.458 5 4.502 ;
        RECT 5.152 5.578 5.216 5.622 ;
        RECT 5.152 4.458 5.216 4.502 ;
        RECT 5.368 5.578 5.432 5.622 ;
        RECT 5.368 4.458 5.432 4.502 ;
        RECT 5.8 5.718 5.864 5.762 ;
        RECT 5.8 4.318 5.864 4.362 ;
        RECT 6.232 6.838 6.296 6.882 ;
        RECT 6.232 3.198 6.296 3.242 ;
        RECT 6.664 6.978 6.728 7.022 ;
        RECT 6.664 3.058 6.728 3.102 ;
        RECT 7.096 8.098 7.16 8.142 ;
        RECT 7.096 1.938 7.16 1.982 ;
        RECT 7.528 8.238 7.592 8.282 ;
        RECT 7.528 1.798 7.592 1.842 ;
        RECT 7.96 9.358 8.024 9.402 ;
        RECT 7.96 0.678 8.024 0.722 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 9.538 0.022 ;
        RECT -0.034 1.238 9.538 1.282 ;
        RECT 7.958 1.148 8.026 1.282 ;
        RECT 7.526 1.238 7.594 1.372 ;
        RECT 1.91 1.238 1.978 1.372 ;
        RECT 1.478 1.148 1.546 1.282 ;
        RECT -0.034 2.498 9.538 2.542 ;
        RECT 7.094 2.408 7.162 2.542 ;
        RECT 6.662 2.498 6.73 2.632 ;
        RECT 2.774 2.498 2.842 2.632 ;
        RECT 2.342 2.408 2.41 2.542 ;
        RECT -0.034 3.758 9.538 3.802 ;
        RECT 6.23 3.668 6.298 3.802 ;
        RECT 5.798 3.758 5.866 3.892 ;
        RECT 3.638 3.758 3.706 3.892 ;
        RECT 3.206 3.668 3.274 3.802 ;
        RECT -0.034 5.018 9.538 5.062 ;
        RECT 5.366 4.838 5.434 5.242 ;
        RECT 5.15 4.838 5.218 5.242 ;
        RECT 4.934 4.838 5.002 5.242 ;
        RECT 4.07 5.288 4.786 5.332 ;
        RECT 4.718 4.748 4.786 5.332 ;
        RECT 4.07 4.748 4.786 4.792 ;
        RECT 4.502 4.838 4.57 5.242 ;
        RECT 4.394 5.108 4.462 5.332 ;
        RECT 4.394 4.748 4.462 4.972 ;
        RECT 4.178 4.838 4.246 5.242 ;
        RECT 4.07 5.108 4.138 5.332 ;
        RECT 4.07 4.748 4.138 4.972 ;
        RECT 3.962 4.838 4.03 5.242 ;
        RECT -0.034 6.278 9.538 6.322 ;
        RECT 6.23 6.278 6.298 6.412 ;
        RECT 5.798 6.188 5.866 6.322 ;
        RECT 3.638 6.188 3.706 6.322 ;
        RECT 3.206 6.278 3.274 6.412 ;
        RECT -0.034 7.538 9.538 7.582 ;
        RECT 7.094 7.538 7.162 7.672 ;
        RECT 6.662 7.448 6.73 7.582 ;
        RECT 2.774 7.448 2.842 7.582 ;
        RECT 2.342 7.538 2.41 7.672 ;
        RECT -0.034 8.798 9.538 8.842 ;
        RECT 7.958 8.798 8.026 8.932 ;
        RECT 7.526 8.708 7.594 8.842 ;
        RECT 1.91 8.708 1.978 8.842 ;
        RECT 1.478 8.798 1.546 8.932 ;
        RECT -0.034 10.058 9.538 10.102 ;
      LAYER v0 ;
        RECT 1.48 8.868 1.544 8.912 ;
        RECT 1.48 1.168 1.544 1.212 ;
        RECT 1.912 8.728 1.976 8.772 ;
        RECT 1.912 1.308 1.976 1.352 ;
        RECT 2.344 7.608 2.408 7.652 ;
        RECT 2.344 2.428 2.408 2.472 ;
        RECT 2.776 7.468 2.84 7.512 ;
        RECT 2.776 2.568 2.84 2.612 ;
        RECT 3.208 6.348 3.272 6.392 ;
        RECT 3.208 3.688 3.272 3.732 ;
        RECT 3.64 6.208 3.704 6.252 ;
        RECT 3.64 3.828 3.704 3.872 ;
        RECT 3.962 5.108 4.03 5.152 ;
        RECT 3.962 4.928 4.03 4.972 ;
        RECT 4.072 5.2155 4.136 5.2595 ;
        RECT 4.072 4.8205 4.136 4.8645 ;
        RECT 4.178 5.108 4.246 5.152 ;
        RECT 4.178 4.928 4.246 4.972 ;
        RECT 4.396 5.2155 4.46 5.2595 ;
        RECT 4.396 4.8205 4.46 4.8645 ;
        RECT 4.502 5.108 4.57 5.152 ;
        RECT 4.502 4.928 4.57 4.972 ;
        RECT 4.934 5.108 5.002 5.152 ;
        RECT 4.934 4.928 5.002 4.972 ;
        RECT 5.15 5.108 5.218 5.152 ;
        RECT 5.15 4.928 5.218 4.972 ;
        RECT 5.366 5.108 5.434 5.152 ;
        RECT 5.366 4.928 5.434 4.972 ;
        RECT 5.8 6.208 5.864 6.252 ;
        RECT 5.8 3.828 5.864 3.872 ;
        RECT 6.232 6.348 6.296 6.392 ;
        RECT 6.232 3.688 6.296 3.732 ;
        RECT 6.664 7.468 6.728 7.512 ;
        RECT 6.664 2.568 6.728 2.612 ;
        RECT 7.096 7.608 7.16 7.652 ;
        RECT 7.096 2.428 7.16 2.472 ;
        RECT 7.528 8.728 7.592 8.772 ;
        RECT 7.528 1.308 7.592 1.352 ;
        RECT 7.96 8.868 8.024 8.912 ;
        RECT 7.96 1.168 8.024 1.212 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 9.608 0.142 9.922 ;
      RECT 0.074 8.978 0.142 9.292 ;
      RECT 0.074 8.348 0.142 8.662 ;
      RECT 0.074 7.718 0.142 8.032 ;
      RECT 0.074 7.088 0.142 7.402 ;
      RECT 0.074 6.458 0.142 6.772 ;
      RECT 0.074 5.828 0.142 6.142 ;
      RECT 0.074 5.198 0.142 5.512 ;
      RECT 0.074 4.568 0.142 4.882 ;
      RECT 0.074 3.938 0.142 4.252 ;
      RECT 0.074 3.308 0.142 3.622 ;
      RECT 0.074 2.678 0.142 2.992 ;
      RECT 0.074 2.048 0.142 2.362 ;
      RECT 0.074 1.418 0.142 1.732 ;
      RECT 0.074 0.788 0.142 1.102 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.182 9.608 0.25 9.922 ;
      RECT 0.182 8.978 0.25 9.292 ;
      RECT 0.182 8.348 0.25 8.662 ;
      RECT 0.182 7.718 0.25 8.032 ;
      RECT 0.182 7.088 0.25 7.402 ;
      RECT 0.182 6.458 0.25 6.772 ;
      RECT 0.182 5.828 0.25 6.142 ;
      RECT 0.182 5.198 0.25 5.512 ;
      RECT 0.182 4.568 0.25 4.882 ;
      RECT 0.182 3.938 0.25 4.252 ;
      RECT 0.182 3.308 0.25 3.622 ;
      RECT 0.182 2.678 0.25 2.992 ;
      RECT 0.182 2.048 0.25 2.362 ;
      RECT 0.182 1.418 0.25 1.732 ;
      RECT 0.182 0.788 0.25 1.102 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.29 9.608 0.358 9.922 ;
      RECT 0.29 8.978 0.358 9.292 ;
      RECT 0.29 8.348 0.358 8.662 ;
      RECT 0.29 7.718 0.358 8.032 ;
      RECT 0.29 7.088 0.358 7.402 ;
      RECT 0.29 6.458 0.358 6.772 ;
      RECT 0.29 5.828 0.358 6.142 ;
      RECT 0.29 5.198 0.358 5.512 ;
      RECT 0.29 4.568 0.358 4.882 ;
      RECT 0.29 3.938 0.358 4.252 ;
      RECT 0.29 3.308 0.358 3.622 ;
      RECT 0.29 2.678 0.358 2.992 ;
      RECT 0.29 2.048 0.358 2.362 ;
      RECT 0.29 1.418 0.358 1.732 ;
      RECT 0.29 0.788 0.358 1.102 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.054 9.968 0.378 10.012 ;
      RECT 0.054 9.518 0.378 9.562 ;
      RECT 0.054 9.338 0.378 9.382 ;
      RECT 0.054 8.888 0.378 8.932 ;
      RECT 0.054 8.708 0.378 8.752 ;
      RECT 0.054 8.258 0.378 8.302 ;
      RECT 0.054 8.078 0.378 8.122 ;
      RECT 0.054 7.628 0.378 7.672 ;
      RECT 0.054 7.448 0.378 7.492 ;
      RECT 0.054 6.998 0.378 7.042 ;
      RECT 0.054 6.818 0.378 6.862 ;
      RECT 0.054 6.368 0.378 6.412 ;
      RECT 0.054 6.188 0.378 6.232 ;
      RECT 0.054 5.738 0.378 5.782 ;
      RECT 0.054 5.558 0.378 5.602 ;
      RECT 0.054 5.108 0.378 5.152 ;
      RECT 0.054 4.928 0.378 4.972 ;
      RECT 0.054 4.478 0.378 4.522 ;
      RECT 0.054 4.298 0.378 4.342 ;
      RECT 0.054 3.848 0.378 3.892 ;
      RECT 0.054 3.668 0.378 3.712 ;
      RECT 0.054 3.218 0.378 3.262 ;
      RECT 0.054 3.038 0.378 3.082 ;
      RECT 0.054 2.588 0.378 2.632 ;
      RECT 0.054 2.408 0.378 2.452 ;
      RECT 0.054 1.958 0.378 2.002 ;
      RECT 0.054 1.778 0.378 1.822 ;
      RECT 0.054 1.328 0.378 1.372 ;
      RECT 0.054 1.148 0.378 1.192 ;
      RECT 0.054 0.698 0.378 0.742 ;
      RECT 0.054 0.518 0.378 0.562 ;
      RECT 0.054 0.068 0.378 0.112 ;
      RECT 0.506 9.608 0.574 9.922 ;
      RECT 0.506 8.978 0.574 9.292 ;
      RECT 0.506 8.348 0.574 8.662 ;
      RECT 0.506 7.718 0.574 8.032 ;
      RECT 0.506 7.088 0.574 7.402 ;
      RECT 0.506 6.458 0.574 6.772 ;
      RECT 0.506 5.828 0.574 6.142 ;
      RECT 0.506 5.198 0.574 5.512 ;
      RECT 0.506 4.568 0.574 4.882 ;
      RECT 0.506 3.938 0.574 4.252 ;
      RECT 0.506 3.308 0.574 3.622 ;
      RECT 0.506 2.678 0.574 2.992 ;
      RECT 0.506 2.048 0.574 2.362 ;
      RECT 0.506 1.418 0.574 1.732 ;
      RECT 0.506 0.788 0.574 1.102 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.614 9.608 0.682 9.922 ;
      RECT 0.614 8.978 0.682 9.292 ;
      RECT 0.614 8.348 0.682 8.662 ;
      RECT 0.614 7.718 0.682 8.032 ;
      RECT 0.614 7.088 0.682 7.402 ;
      RECT 0.614 6.458 0.682 6.772 ;
      RECT 0.614 5.828 0.682 6.142 ;
      RECT 0.614 5.198 0.682 5.512 ;
      RECT 0.614 4.568 0.682 4.882 ;
      RECT 0.614 3.938 0.682 4.252 ;
      RECT 0.614 3.308 0.682 3.622 ;
      RECT 0.614 2.678 0.682 2.992 ;
      RECT 0.614 2.048 0.682 2.362 ;
      RECT 0.614 1.418 0.682 1.732 ;
      RECT 0.614 0.788 0.682 1.102 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.722 9.608 0.79 9.922 ;
      RECT 0.722 8.978 0.79 9.292 ;
      RECT 0.722 8.348 0.79 8.662 ;
      RECT 0.722 7.718 0.79 8.032 ;
      RECT 0.722 7.088 0.79 7.402 ;
      RECT 0.722 6.458 0.79 6.772 ;
      RECT 0.722 5.828 0.79 6.142 ;
      RECT 0.722 5.198 0.79 5.512 ;
      RECT 0.722 4.568 0.79 4.882 ;
      RECT 0.722 3.938 0.79 4.252 ;
      RECT 0.722 3.308 0.79 3.622 ;
      RECT 0.722 2.678 0.79 2.992 ;
      RECT 0.722 2.048 0.79 2.362 ;
      RECT 0.722 1.418 0.79 1.732 ;
      RECT 0.722 0.788 0.79 1.102 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.486 9.968 0.81 10.012 ;
      RECT 0.486 9.518 0.81 9.562 ;
      RECT 0.486 9.338 0.81 9.382 ;
      RECT 0.486 8.888 0.81 8.932 ;
      RECT 0.486 8.708 0.81 8.752 ;
      RECT 0.486 8.258 0.81 8.302 ;
      RECT 0.486 8.078 0.81 8.122 ;
      RECT 0.486 7.628 0.81 7.672 ;
      RECT 0.486 7.448 0.81 7.492 ;
      RECT 0.486 6.998 0.81 7.042 ;
      RECT 0.486 6.818 0.81 6.862 ;
      RECT 0.486 6.368 0.81 6.412 ;
      RECT 0.486 6.188 0.81 6.232 ;
      RECT 0.486 5.738 0.81 5.782 ;
      RECT 0.486 5.558 0.81 5.602 ;
      RECT 0.486 5.108 0.81 5.152 ;
      RECT 0.486 4.928 0.81 4.972 ;
      RECT 0.486 4.478 0.81 4.522 ;
      RECT 0.486 4.298 0.81 4.342 ;
      RECT 0.486 3.848 0.81 3.892 ;
      RECT 0.486 3.668 0.81 3.712 ;
      RECT 0.486 3.218 0.81 3.262 ;
      RECT 0.486 3.038 0.81 3.082 ;
      RECT 0.486 2.588 0.81 2.632 ;
      RECT 0.486 2.408 0.81 2.452 ;
      RECT 0.486 1.958 0.81 2.002 ;
      RECT 0.486 1.778 0.81 1.822 ;
      RECT 0.486 1.328 0.81 1.372 ;
      RECT 0.486 1.148 0.81 1.192 ;
      RECT 0.486 0.698 0.81 0.742 ;
      RECT 0.486 0.518 0.81 0.562 ;
      RECT 0.486 0.068 0.81 0.112 ;
      RECT 0.938 9.608 1.006 9.922 ;
      RECT 0.938 8.978 1.006 9.292 ;
      RECT 0.938 8.348 1.006 8.662 ;
      RECT 0.938 7.718 1.006 8.032 ;
      RECT 0.938 7.088 1.006 7.402 ;
      RECT 0.938 6.458 1.006 6.772 ;
      RECT 0.938 5.828 1.006 6.142 ;
      RECT 0.938 5.198 1.006 5.512 ;
      RECT 0.938 4.568 1.006 4.882 ;
      RECT 0.938 3.938 1.006 4.252 ;
      RECT 0.938 3.308 1.006 3.622 ;
      RECT 0.938 2.678 1.006 2.992 ;
      RECT 0.938 2.048 1.006 2.362 ;
      RECT 0.938 1.418 1.006 1.732 ;
      RECT 0.938 0.788 1.006 1.102 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.046 9.608 1.114 9.922 ;
      RECT 1.046 9.158 1.114 9.292 ;
      RECT 1.046 8.978 1.114 9.112 ;
      RECT 1.046 8.348 1.114 8.662 ;
      RECT 1.046 7.718 1.114 8.032 ;
      RECT 1.046 7.088 1.114 7.402 ;
      RECT 1.046 6.458 1.114 6.772 ;
      RECT 1.046 5.828 1.114 6.142 ;
      RECT 1.046 5.198 1.114 5.512 ;
      RECT 1.046 4.568 1.114 4.882 ;
      RECT 1.046 3.938 1.114 4.252 ;
      RECT 1.046 3.308 1.114 3.622 ;
      RECT 1.046 2.678 1.114 2.992 ;
      RECT 1.046 2.048 1.114 2.362 ;
      RECT 1.046 1.418 1.114 1.732 ;
      RECT 1.046 0.968 1.114 1.102 ;
      RECT 1.046 0.788 1.114 0.922 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.154 9.608 1.222 9.922 ;
      RECT 1.154 8.978 1.222 9.292 ;
      RECT 1.154 8.348 1.222 8.662 ;
      RECT 1.154 7.718 1.222 8.032 ;
      RECT 1.154 7.088 1.222 7.402 ;
      RECT 1.154 6.458 1.222 6.772 ;
      RECT 1.154 5.828 1.222 6.142 ;
      RECT 1.154 5.198 1.222 5.512 ;
      RECT 1.154 4.568 1.222 4.882 ;
      RECT 1.154 3.938 1.222 4.252 ;
      RECT 1.154 3.308 1.222 3.622 ;
      RECT 1.154 2.678 1.222 2.992 ;
      RECT 1.154 2.048 1.222 2.362 ;
      RECT 1.154 1.418 1.222 1.732 ;
      RECT 1.154 0.788 1.222 1.102 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.918 9.968 1.242 10.012 ;
      RECT 0.918 9.518 1.242 9.562 ;
      RECT 0.918 8.708 1.242 8.752 ;
      RECT 0.918 8.258 1.242 8.302 ;
      RECT 0.918 8.078 1.242 8.122 ;
      RECT 0.918 7.628 1.242 7.672 ;
      RECT 0.918 7.448 1.242 7.492 ;
      RECT 0.918 6.998 1.242 7.042 ;
      RECT 0.918 6.818 1.242 6.862 ;
      RECT 0.918 6.368 1.242 6.412 ;
      RECT 0.918 6.188 1.242 6.232 ;
      RECT 0.918 5.738 1.242 5.782 ;
      RECT 0.918 5.558 1.242 5.602 ;
      RECT 0.918 5.108 1.242 5.152 ;
      RECT 0.918 4.928 1.242 4.972 ;
      RECT 0.918 4.478 1.242 4.522 ;
      RECT 0.918 4.298 1.242 4.342 ;
      RECT 0.918 3.848 1.242 3.892 ;
      RECT 0.918 3.668 1.242 3.712 ;
      RECT 0.918 3.218 1.242 3.262 ;
      RECT 0.918 3.038 1.242 3.082 ;
      RECT 0.918 2.588 1.242 2.632 ;
      RECT 0.918 2.408 1.242 2.452 ;
      RECT 0.918 1.958 1.242 2.002 ;
      RECT 0.918 1.778 1.242 1.822 ;
      RECT 0.918 1.328 1.242 1.372 ;
      RECT 0.918 0.518 1.242 0.562 ;
      RECT 0.918 0.068 1.242 0.112 ;
      RECT 1.262 8.978 1.33 9.292 ;
      RECT 1.262 0.788 1.33 1.102 ;
      RECT 1.37 9.608 1.438 9.922 ;
      RECT 1.37 9.158 1.438 9.292 ;
      RECT 1.37 8.978 1.438 9.112 ;
      RECT 1.37 8.348 1.438 8.662 ;
      RECT 1.37 7.718 1.438 8.032 ;
      RECT 1.37 7.088 1.438 7.402 ;
      RECT 1.37 6.458 1.438 6.772 ;
      RECT 1.37 5.828 1.438 6.142 ;
      RECT 1.37 5.198 1.438 5.512 ;
      RECT 1.37 4.568 1.438 4.882 ;
      RECT 1.37 3.938 1.438 4.252 ;
      RECT 1.37 3.308 1.438 3.622 ;
      RECT 1.37 2.678 1.438 2.992 ;
      RECT 1.37 2.048 1.438 2.362 ;
      RECT 1.37 1.418 1.438 1.732 ;
      RECT 1.37 0.968 1.438 1.102 ;
      RECT 1.37 0.788 1.438 0.922 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 1.478 9.608 1.546 9.922 ;
      RECT 1.478 8.528 1.546 8.662 ;
      RECT 1.478 8.348 1.546 8.482 ;
      RECT 1.478 7.718 1.546 8.032 ;
      RECT 1.478 7.088 1.546 7.402 ;
      RECT 1.478 6.458 1.546 6.772 ;
      RECT 1.478 5.828 1.546 6.142 ;
      RECT 1.478 5.198 1.546 5.512 ;
      RECT 1.478 4.568 1.546 4.882 ;
      RECT 1.478 3.938 1.546 4.252 ;
      RECT 1.478 3.308 1.546 3.622 ;
      RECT 1.478 2.678 1.546 2.992 ;
      RECT 1.478 2.048 1.546 2.362 ;
      RECT 1.478 1.598 1.546 1.732 ;
      RECT 1.478 1.418 1.546 1.552 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.586 9.608 1.654 9.922 ;
      RECT 1.586 9.158 1.654 9.292 ;
      RECT 1.586 8.978 1.654 9.112 ;
      RECT 1.586 8.348 1.654 8.662 ;
      RECT 1.586 7.718 1.654 8.032 ;
      RECT 1.586 7.088 1.654 7.402 ;
      RECT 1.586 6.458 1.654 6.772 ;
      RECT 1.586 5.828 1.654 6.142 ;
      RECT 1.586 5.198 1.654 5.512 ;
      RECT 1.586 4.568 1.654 4.882 ;
      RECT 1.586 3.938 1.654 4.252 ;
      RECT 1.586 3.308 1.654 3.622 ;
      RECT 1.586 2.678 1.654 2.992 ;
      RECT 1.586 2.048 1.654 2.362 ;
      RECT 1.586 1.418 1.654 1.732 ;
      RECT 1.586 0.968 1.654 1.102 ;
      RECT 1.586 0.788 1.654 0.922 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.35 9.968 1.674 10.012 ;
      RECT 1.35 9.518 1.674 9.562 ;
      RECT 1.35 8.078 1.674 8.122 ;
      RECT 1.35 7.628 1.674 7.672 ;
      RECT 1.35 7.448 1.674 7.492 ;
      RECT 1.35 6.998 1.674 7.042 ;
      RECT 1.35 6.818 1.674 6.862 ;
      RECT 1.35 6.368 1.674 6.412 ;
      RECT 1.35 6.188 1.674 6.232 ;
      RECT 1.35 5.738 1.674 5.782 ;
      RECT 1.35 5.558 1.674 5.602 ;
      RECT 1.35 5.108 1.674 5.152 ;
      RECT 1.35 4.928 1.674 4.972 ;
      RECT 1.35 4.478 1.674 4.522 ;
      RECT 1.35 4.298 1.674 4.342 ;
      RECT 1.35 3.848 1.674 3.892 ;
      RECT 1.35 3.668 1.674 3.712 ;
      RECT 1.35 3.218 1.674 3.262 ;
      RECT 1.35 3.038 1.674 3.082 ;
      RECT 1.35 2.588 1.674 2.632 ;
      RECT 1.35 2.408 1.674 2.452 ;
      RECT 1.35 1.958 1.674 2.002 ;
      RECT 1.35 0.518 1.674 0.562 ;
      RECT 1.35 0.068 1.674 0.112 ;
      RECT 1.694 8.978 1.762 9.292 ;
      RECT 1.694 8.348 1.762 8.662 ;
      RECT 1.694 1.418 1.762 1.732 ;
      RECT 1.694 0.788 1.762 1.102 ;
      RECT 1.802 9.608 1.87 9.922 ;
      RECT 1.802 8.978 1.87 9.292 ;
      RECT 1.802 8.528 1.87 8.662 ;
      RECT 1.802 8.348 1.87 8.482 ;
      RECT 1.802 7.718 1.87 8.032 ;
      RECT 1.802 7.088 1.87 7.402 ;
      RECT 1.802 6.458 1.87 6.772 ;
      RECT 1.802 5.828 1.87 6.142 ;
      RECT 1.802 5.198 1.87 5.512 ;
      RECT 1.802 4.568 1.87 4.882 ;
      RECT 1.802 3.938 1.87 4.252 ;
      RECT 1.802 3.308 1.87 3.622 ;
      RECT 1.802 2.678 1.87 2.992 ;
      RECT 1.802 2.048 1.87 2.362 ;
      RECT 1.802 1.598 1.87 1.732 ;
      RECT 1.802 1.418 1.87 1.552 ;
      RECT 1.802 0.788 1.87 1.102 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 1.91 9.608 1.978 9.922 ;
      RECT 1.91 9.158 1.978 9.292 ;
      RECT 1.91 8.978 1.978 9.112 ;
      RECT 1.91 7.898 1.978 8.032 ;
      RECT 1.91 7.718 1.978 7.852 ;
      RECT 1.91 7.088 1.978 7.402 ;
      RECT 1.91 6.458 1.978 6.772 ;
      RECT 1.91 5.828 1.978 6.142 ;
      RECT 1.91 5.198 1.978 5.512 ;
      RECT 1.91 4.568 1.978 4.882 ;
      RECT 1.91 3.938 1.978 4.252 ;
      RECT 1.91 3.308 1.978 3.622 ;
      RECT 1.91 2.678 1.978 2.992 ;
      RECT 1.91 2.228 1.978 2.362 ;
      RECT 1.91 2.048 1.978 2.182 ;
      RECT 1.91 0.968 1.978 1.102 ;
      RECT 1.91 0.788 1.978 0.922 ;
      RECT 1.91 0.158 1.978 0.472 ;
      RECT 2.018 9.608 2.086 9.922 ;
      RECT 2.018 8.978 2.086 9.292 ;
      RECT 2.018 8.528 2.086 8.662 ;
      RECT 2.018 8.348 2.086 8.482 ;
      RECT 2.018 7.718 2.086 8.032 ;
      RECT 2.018 7.088 2.086 7.402 ;
      RECT 2.018 6.458 2.086 6.772 ;
      RECT 2.018 5.828 2.086 6.142 ;
      RECT 2.018 5.198 2.086 5.512 ;
      RECT 2.018 4.568 2.086 4.882 ;
      RECT 2.018 3.938 2.086 4.252 ;
      RECT 2.018 3.308 2.086 3.622 ;
      RECT 2.018 2.678 2.086 2.992 ;
      RECT 2.018 2.048 2.086 2.362 ;
      RECT 2.018 1.598 2.086 1.732 ;
      RECT 2.018 1.418 2.086 1.552 ;
      RECT 2.018 0.788 2.086 1.102 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 1.782 9.968 2.106 10.012 ;
      RECT 1.782 9.518 2.106 9.562 ;
      RECT 1.782 7.448 2.106 7.492 ;
      RECT 1.782 6.998 2.106 7.042 ;
      RECT 1.782 6.818 2.106 6.862 ;
      RECT 1.782 6.368 2.106 6.412 ;
      RECT 1.782 6.188 2.106 6.232 ;
      RECT 1.782 5.738 2.106 5.782 ;
      RECT 1.782 5.558 2.106 5.602 ;
      RECT 1.782 5.108 2.106 5.152 ;
      RECT 1.782 4.928 2.106 4.972 ;
      RECT 1.782 4.478 2.106 4.522 ;
      RECT 1.782 4.298 2.106 4.342 ;
      RECT 1.782 3.848 2.106 3.892 ;
      RECT 1.782 3.668 2.106 3.712 ;
      RECT 1.782 3.218 2.106 3.262 ;
      RECT 1.782 3.038 2.106 3.082 ;
      RECT 1.782 2.588 2.106 2.632 ;
      RECT 1.782 0.518 2.106 0.562 ;
      RECT 1.782 0.068 2.106 0.112 ;
      RECT 2.126 8.348 2.194 8.662 ;
      RECT 2.126 7.718 2.194 8.032 ;
      RECT 2.126 2.048 2.194 2.362 ;
      RECT 2.126 1.418 2.194 1.732 ;
      RECT 2.234 9.608 2.302 9.922 ;
      RECT 2.234 8.978 2.302 9.292 ;
      RECT 2.234 8.348 2.302 8.662 ;
      RECT 2.234 7.898 2.302 8.032 ;
      RECT 2.234 7.718 2.302 7.852 ;
      RECT 2.234 7.088 2.302 7.402 ;
      RECT 2.234 6.458 2.302 6.772 ;
      RECT 2.234 5.828 2.302 6.142 ;
      RECT 2.234 5.198 2.302 5.512 ;
      RECT 2.234 4.568 2.302 4.882 ;
      RECT 2.234 3.938 2.302 4.252 ;
      RECT 2.234 3.308 2.302 3.622 ;
      RECT 2.234 2.678 2.302 2.992 ;
      RECT 2.234 2.228 2.302 2.362 ;
      RECT 2.234 2.048 2.302 2.182 ;
      RECT 2.234 1.418 2.302 1.732 ;
      RECT 2.234 0.788 2.302 1.102 ;
      RECT 2.234 0.158 2.302 0.472 ;
      RECT 2.342 9.608 2.41 9.922 ;
      RECT 2.342 8.978 2.41 9.292 ;
      RECT 2.342 8.528 2.41 8.662 ;
      RECT 2.342 8.348 2.41 8.482 ;
      RECT 2.342 7.268 2.41 7.402 ;
      RECT 2.342 7.088 2.41 7.222 ;
      RECT 2.342 6.458 2.41 6.772 ;
      RECT 2.342 5.828 2.41 6.142 ;
      RECT 2.342 5.198 2.41 5.512 ;
      RECT 2.342 4.568 2.41 4.882 ;
      RECT 2.342 3.938 2.41 4.252 ;
      RECT 2.342 3.308 2.41 3.622 ;
      RECT 2.342 2.858 2.41 2.992 ;
      RECT 2.342 2.678 2.41 2.812 ;
      RECT 2.342 1.598 2.41 1.732 ;
      RECT 2.342 1.418 2.41 1.552 ;
      RECT 2.342 0.788 2.41 1.102 ;
      RECT 2.342 0.158 2.41 0.472 ;
      RECT 2.45 9.608 2.518 9.922 ;
      RECT 2.45 8.978 2.518 9.292 ;
      RECT 2.45 8.348 2.518 8.662 ;
      RECT 2.45 7.898 2.518 8.032 ;
      RECT 2.45 7.718 2.518 7.852 ;
      RECT 2.45 7.088 2.518 7.402 ;
      RECT 2.45 6.458 2.518 6.772 ;
      RECT 2.45 5.828 2.518 6.142 ;
      RECT 2.45 5.198 2.518 5.512 ;
      RECT 2.45 4.568 2.518 4.882 ;
      RECT 2.45 3.938 2.518 4.252 ;
      RECT 2.45 3.308 2.518 3.622 ;
      RECT 2.45 2.678 2.518 2.992 ;
      RECT 2.45 2.228 2.518 2.362 ;
      RECT 2.45 2.048 2.518 2.182 ;
      RECT 2.45 1.418 2.518 1.732 ;
      RECT 2.45 0.788 2.518 1.102 ;
      RECT 2.45 0.158 2.518 0.472 ;
      RECT 2.214 9.968 2.538 10.012 ;
      RECT 2.214 9.518 2.538 9.562 ;
      RECT 2.214 9.338 2.538 9.382 ;
      RECT 2.214 8.888 2.538 8.932 ;
      RECT 2.214 6.818 2.538 6.862 ;
      RECT 2.214 6.368 2.538 6.412 ;
      RECT 2.214 6.188 2.538 6.232 ;
      RECT 2.214 5.738 2.538 5.782 ;
      RECT 2.214 5.558 2.538 5.602 ;
      RECT 2.214 5.108 2.538 5.152 ;
      RECT 2.214 4.928 2.538 4.972 ;
      RECT 2.214 4.478 2.538 4.522 ;
      RECT 2.214 4.298 2.538 4.342 ;
      RECT 2.214 3.848 2.538 3.892 ;
      RECT 2.214 3.668 2.538 3.712 ;
      RECT 2.214 3.218 2.538 3.262 ;
      RECT 2.214 1.148 2.538 1.192 ;
      RECT 2.214 0.698 2.538 0.742 ;
      RECT 2.214 0.518 2.538 0.562 ;
      RECT 2.214 0.068 2.538 0.112 ;
      RECT 2.558 7.718 2.626 8.032 ;
      RECT 2.558 7.088 2.626 7.402 ;
      RECT 2.558 2.678 2.626 2.992 ;
      RECT 2.558 2.048 2.626 2.362 ;
      RECT 2.666 9.608 2.734 9.922 ;
      RECT 2.666 8.978 2.734 9.292 ;
      RECT 2.666 8.348 2.734 8.662 ;
      RECT 2.666 7.718 2.734 8.032 ;
      RECT 2.666 7.268 2.734 7.402 ;
      RECT 2.666 7.088 2.734 7.222 ;
      RECT 2.666 6.458 2.734 6.772 ;
      RECT 2.666 5.828 2.734 6.142 ;
      RECT 2.666 5.198 2.734 5.512 ;
      RECT 2.666 4.568 2.734 4.882 ;
      RECT 2.666 3.938 2.734 4.252 ;
      RECT 2.666 3.308 2.734 3.622 ;
      RECT 2.666 2.858 2.734 2.992 ;
      RECT 2.666 2.678 2.734 2.812 ;
      RECT 2.666 2.048 2.734 2.362 ;
      RECT 2.666 1.418 2.734 1.732 ;
      RECT 2.666 0.788 2.734 1.102 ;
      RECT 2.666 0.158 2.734 0.472 ;
      RECT 2.774 9.608 2.842 9.922 ;
      RECT 2.774 8.978 2.842 9.292 ;
      RECT 2.774 8.348 2.842 8.662 ;
      RECT 2.774 7.898 2.842 8.032 ;
      RECT 2.774 7.718 2.842 7.852 ;
      RECT 2.774 6.638 2.842 6.772 ;
      RECT 2.774 6.458 2.842 6.592 ;
      RECT 2.774 5.828 2.842 6.142 ;
      RECT 2.774 5.198 2.842 5.512 ;
      RECT 2.774 4.568 2.842 4.882 ;
      RECT 2.774 3.938 2.842 4.252 ;
      RECT 2.774 3.488 2.842 3.622 ;
      RECT 2.774 3.308 2.842 3.442 ;
      RECT 2.774 2.228 2.842 2.362 ;
      RECT 2.774 2.048 2.842 2.182 ;
      RECT 2.774 1.418 2.842 1.732 ;
      RECT 2.774 0.788 2.842 1.102 ;
      RECT 2.774 0.158 2.842 0.472 ;
      RECT 2.882 9.608 2.95 9.922 ;
      RECT 2.882 8.978 2.95 9.292 ;
      RECT 2.882 8.348 2.95 8.662 ;
      RECT 2.882 7.718 2.95 8.032 ;
      RECT 2.882 7.268 2.95 7.402 ;
      RECT 2.882 7.088 2.95 7.222 ;
      RECT 2.882 6.458 2.95 6.772 ;
      RECT 2.882 5.828 2.95 6.142 ;
      RECT 2.882 5.198 2.95 5.512 ;
      RECT 2.882 4.568 2.95 4.882 ;
      RECT 2.882 3.938 2.95 4.252 ;
      RECT 2.882 3.308 2.95 3.622 ;
      RECT 2.882 2.858 2.95 2.992 ;
      RECT 2.882 2.678 2.95 2.812 ;
      RECT 2.882 2.048 2.95 2.362 ;
      RECT 2.882 1.418 2.95 1.732 ;
      RECT 2.882 0.788 2.95 1.102 ;
      RECT 2.882 0.158 2.95 0.472 ;
      RECT 2.646 9.968 2.97 10.012 ;
      RECT 2.646 9.518 2.97 9.562 ;
      RECT 2.646 9.338 2.97 9.382 ;
      RECT 2.646 8.888 2.97 8.932 ;
      RECT 2.646 8.708 2.97 8.752 ;
      RECT 2.646 8.258 2.97 8.302 ;
      RECT 2.646 6.188 2.97 6.232 ;
      RECT 2.646 5.738 2.97 5.782 ;
      RECT 2.646 5.558 2.97 5.602 ;
      RECT 2.646 5.108 2.97 5.152 ;
      RECT 2.646 4.928 2.97 4.972 ;
      RECT 2.646 4.478 2.97 4.522 ;
      RECT 2.646 4.298 2.97 4.342 ;
      RECT 2.646 3.848 2.97 3.892 ;
      RECT 2.646 1.778 2.97 1.822 ;
      RECT 2.646 1.328 2.97 1.372 ;
      RECT 2.646 1.148 2.97 1.192 ;
      RECT 2.646 0.698 2.97 0.742 ;
      RECT 2.646 0.518 2.97 0.562 ;
      RECT 2.646 0.068 2.97 0.112 ;
      RECT 2.99 7.088 3.058 7.402 ;
      RECT 2.99 6.458 3.058 6.772 ;
      RECT 2.99 3.308 3.058 3.622 ;
      RECT 2.99 2.678 3.058 2.992 ;
      RECT 3.098 9.608 3.166 9.922 ;
      RECT 3.098 8.978 3.166 9.292 ;
      RECT 3.098 8.348 3.166 8.662 ;
      RECT 3.098 7.718 3.166 8.032 ;
      RECT 3.098 7.088 3.166 7.402 ;
      RECT 3.098 6.638 3.166 6.772 ;
      RECT 3.098 6.458 3.166 6.592 ;
      RECT 3.098 5.828 3.166 6.142 ;
      RECT 3.098 5.198 3.166 5.512 ;
      RECT 3.098 4.568 3.166 4.882 ;
      RECT 3.098 3.938 3.166 4.252 ;
      RECT 3.098 3.488 3.166 3.622 ;
      RECT 3.098 3.308 3.166 3.442 ;
      RECT 3.098 2.678 3.166 2.992 ;
      RECT 3.098 2.048 3.166 2.362 ;
      RECT 3.098 1.418 3.166 1.732 ;
      RECT 3.098 0.788 3.166 1.102 ;
      RECT 3.098 0.158 3.166 0.472 ;
      RECT 3.206 9.608 3.274 9.922 ;
      RECT 3.206 8.978 3.274 9.292 ;
      RECT 3.206 8.348 3.274 8.662 ;
      RECT 3.206 7.718 3.274 8.032 ;
      RECT 3.206 7.268 3.274 7.402 ;
      RECT 3.206 7.088 3.274 7.222 ;
      RECT 3.206 6.008 3.274 6.142 ;
      RECT 3.206 5.828 3.274 5.962 ;
      RECT 3.206 5.198 3.274 5.512 ;
      RECT 3.206 4.568 3.274 4.882 ;
      RECT 3.206 4.118 3.274 4.252 ;
      RECT 3.206 3.938 3.274 4.072 ;
      RECT 3.206 2.858 3.274 2.992 ;
      RECT 3.206 2.678 3.274 2.812 ;
      RECT 3.206 2.048 3.274 2.362 ;
      RECT 3.206 1.418 3.274 1.732 ;
      RECT 3.206 0.788 3.274 1.102 ;
      RECT 3.206 0.158 3.274 0.472 ;
      RECT 3.314 9.608 3.382 9.922 ;
      RECT 3.314 8.978 3.382 9.292 ;
      RECT 3.314 8.348 3.382 8.662 ;
      RECT 3.314 7.718 3.382 8.032 ;
      RECT 3.314 7.088 3.382 7.402 ;
      RECT 3.314 6.638 3.382 6.772 ;
      RECT 3.314 6.458 3.382 6.592 ;
      RECT 3.314 5.828 3.382 6.142 ;
      RECT 3.314 5.198 3.382 5.512 ;
      RECT 3.314 4.568 3.382 4.882 ;
      RECT 3.314 3.938 3.382 4.252 ;
      RECT 3.314 3.488 3.382 3.622 ;
      RECT 3.314 3.308 3.382 3.442 ;
      RECT 3.314 2.678 3.382 2.992 ;
      RECT 3.314 2.048 3.382 2.362 ;
      RECT 3.314 1.418 3.382 1.732 ;
      RECT 3.314 0.788 3.382 1.102 ;
      RECT 3.314 0.158 3.382 0.472 ;
      RECT 3.078 9.968 3.402 10.012 ;
      RECT 3.078 9.518 3.402 9.562 ;
      RECT 3.078 9.338 3.402 9.382 ;
      RECT 3.078 8.888 3.402 8.932 ;
      RECT 3.078 8.708 3.402 8.752 ;
      RECT 3.078 8.258 3.402 8.302 ;
      RECT 3.078 8.078 3.402 8.122 ;
      RECT 3.078 7.628 3.402 7.672 ;
      RECT 3.078 5.558 3.402 5.602 ;
      RECT 3.078 5.108 3.402 5.152 ;
      RECT 3.078 4.928 3.402 4.972 ;
      RECT 3.078 4.478 3.402 4.522 ;
      RECT 3.078 2.408 3.402 2.452 ;
      RECT 3.078 1.958 3.402 2.002 ;
      RECT 3.078 1.778 3.402 1.822 ;
      RECT 3.078 1.328 3.402 1.372 ;
      RECT 3.078 1.148 3.402 1.192 ;
      RECT 3.078 0.698 3.402 0.742 ;
      RECT 3.078 0.518 3.402 0.562 ;
      RECT 3.078 0.068 3.402 0.112 ;
      RECT 3.422 6.458 3.49 6.772 ;
      RECT 3.422 5.828 3.49 6.142 ;
      RECT 3.422 3.938 3.49 4.252 ;
      RECT 3.422 3.308 3.49 3.622 ;
      RECT 3.53 9.608 3.598 9.922 ;
      RECT 3.53 8.978 3.598 9.292 ;
      RECT 3.53 8.348 3.598 8.662 ;
      RECT 3.53 7.718 3.598 8.032 ;
      RECT 3.53 7.088 3.598 7.402 ;
      RECT 3.53 6.458 3.598 6.772 ;
      RECT 3.53 6.008 3.598 6.142 ;
      RECT 3.53 5.828 3.598 5.962 ;
      RECT 3.53 5.198 3.598 5.512 ;
      RECT 3.53 4.568 3.598 4.882 ;
      RECT 3.53 4.118 3.598 4.252 ;
      RECT 3.53 3.938 3.598 4.072 ;
      RECT 3.53 3.308 3.598 3.622 ;
      RECT 3.53 2.678 3.598 2.992 ;
      RECT 3.53 2.048 3.598 2.362 ;
      RECT 3.53 1.418 3.598 1.732 ;
      RECT 3.53 0.788 3.598 1.102 ;
      RECT 3.53 0.158 3.598 0.472 ;
      RECT 3.638 9.608 3.706 9.922 ;
      RECT 3.638 8.978 3.706 9.292 ;
      RECT 3.638 8.348 3.706 8.662 ;
      RECT 3.638 7.718 3.706 8.032 ;
      RECT 3.638 7.088 3.706 7.402 ;
      RECT 3.638 6.638 3.706 6.772 ;
      RECT 3.638 6.458 3.706 6.592 ;
      RECT 3.638 5.198 3.706 5.512 ;
      RECT 3.638 4.568 3.706 4.882 ;
      RECT 3.638 3.488 3.706 3.622 ;
      RECT 3.638 3.308 3.706 3.442 ;
      RECT 3.638 2.678 3.706 2.992 ;
      RECT 3.638 2.048 3.706 2.362 ;
      RECT 3.638 1.418 3.706 1.732 ;
      RECT 3.638 0.788 3.706 1.102 ;
      RECT 3.638 0.158 3.706 0.472 ;
      RECT 3.746 9.608 3.814 9.922 ;
      RECT 3.746 8.978 3.814 9.292 ;
      RECT 3.746 8.348 3.814 8.662 ;
      RECT 3.746 7.718 3.814 8.032 ;
      RECT 3.746 7.088 3.814 7.402 ;
      RECT 3.746 6.458 3.814 6.772 ;
      RECT 3.746 6.008 3.814 6.142 ;
      RECT 3.746 5.828 3.814 5.962 ;
      RECT 3.746 5.198 3.814 5.512 ;
      RECT 3.746 4.568 3.814 4.882 ;
      RECT 3.746 4.118 3.814 4.252 ;
      RECT 3.746 3.938 3.814 4.072 ;
      RECT 3.746 3.308 3.814 3.622 ;
      RECT 3.746 2.678 3.814 2.992 ;
      RECT 3.746 2.048 3.814 2.362 ;
      RECT 3.746 1.418 3.814 1.732 ;
      RECT 3.746 0.788 3.814 1.102 ;
      RECT 3.746 0.158 3.814 0.472 ;
      RECT 3.51 9.968 3.834 10.012 ;
      RECT 3.51 9.518 3.834 9.562 ;
      RECT 3.51 9.338 3.834 9.382 ;
      RECT 3.51 8.888 3.834 8.932 ;
      RECT 3.51 8.708 3.834 8.752 ;
      RECT 3.51 8.258 3.834 8.302 ;
      RECT 3.51 8.078 3.834 8.122 ;
      RECT 3.51 7.628 3.834 7.672 ;
      RECT 3.51 7.448 3.834 7.492 ;
      RECT 3.51 6.998 3.834 7.042 ;
      RECT 3.51 5.558 3.834 5.602 ;
      RECT 3.51 5.108 3.834 5.152 ;
      RECT 3.51 4.928 3.834 4.972 ;
      RECT 3.51 4.478 3.834 4.522 ;
      RECT 3.51 3.038 3.834 3.082 ;
      RECT 3.51 2.588 3.834 2.632 ;
      RECT 3.51 2.408 3.834 2.452 ;
      RECT 3.51 1.958 3.834 2.002 ;
      RECT 3.51 1.778 3.834 1.822 ;
      RECT 3.51 1.328 3.834 1.372 ;
      RECT 3.51 1.148 3.834 1.192 ;
      RECT 3.51 0.698 3.834 0.742 ;
      RECT 3.51 0.518 3.834 0.562 ;
      RECT 3.51 0.068 3.834 0.112 ;
      RECT 3.854 5.828 3.922 6.142 ;
      RECT 3.854 3.938 3.922 4.252 ;
      RECT 3.962 9.608 4.03 9.922 ;
      RECT 3.962 8.978 4.03 9.292 ;
      RECT 3.962 8.348 4.03 8.662 ;
      RECT 3.962 7.718 4.03 8.032 ;
      RECT 3.962 7.088 4.03 7.402 ;
      RECT 3.962 6.458 4.03 6.772 ;
      RECT 3.962 5.828 4.03 6.142 ;
      RECT 3.962 3.938 4.03 4.252 ;
      RECT 3.962 3.308 4.03 3.622 ;
      RECT 3.962 2.678 4.03 2.992 ;
      RECT 3.962 2.048 4.03 2.362 ;
      RECT 3.962 1.418 4.03 1.732 ;
      RECT 3.962 0.788 4.03 1.102 ;
      RECT 3.962 0.158 4.03 0.472 ;
      RECT 4.07 9.608 4.138 9.922 ;
      RECT 4.07 8.978 4.138 9.292 ;
      RECT 4.07 8.348 4.138 8.662 ;
      RECT 4.07 7.718 4.138 8.032 ;
      RECT 4.07 7.088 4.138 7.402 ;
      RECT 4.07 6.458 4.138 6.772 ;
      RECT 4.07 6.008 4.138 6.142 ;
      RECT 4.07 5.828 4.138 5.962 ;
      RECT 4.07 4.118 4.138 4.252 ;
      RECT 4.07 3.938 4.138 4.072 ;
      RECT 4.07 3.308 4.138 3.622 ;
      RECT 4.07 2.678 4.138 2.992 ;
      RECT 4.07 2.048 4.138 2.362 ;
      RECT 4.07 1.418 4.138 1.732 ;
      RECT 4.07 0.788 4.138 1.102 ;
      RECT 4.07 0.158 4.138 0.472 ;
      RECT 4.178 9.608 4.246 9.922 ;
      RECT 4.178 8.978 4.246 9.292 ;
      RECT 4.178 8.348 4.246 8.662 ;
      RECT 4.178 7.718 4.246 8.032 ;
      RECT 4.178 7.088 4.246 7.402 ;
      RECT 4.178 6.458 4.246 6.772 ;
      RECT 4.178 5.828 4.246 6.142 ;
      RECT 4.178 3.938 4.246 4.252 ;
      RECT 4.178 3.308 4.246 3.622 ;
      RECT 4.178 2.678 4.246 2.992 ;
      RECT 4.178 2.048 4.246 2.362 ;
      RECT 4.178 1.418 4.246 1.732 ;
      RECT 4.178 0.788 4.246 1.102 ;
      RECT 4.178 0.158 4.246 0.472 ;
      RECT 3.942 9.968 4.266 10.012 ;
      RECT 3.942 9.518 4.266 9.562 ;
      RECT 3.942 9.338 4.266 9.382 ;
      RECT 3.942 8.888 4.266 8.932 ;
      RECT 3.942 8.708 4.266 8.752 ;
      RECT 3.942 8.258 4.266 8.302 ;
      RECT 3.942 8.078 4.266 8.122 ;
      RECT 3.942 7.628 4.266 7.672 ;
      RECT 3.942 7.448 4.266 7.492 ;
      RECT 3.942 6.998 4.266 7.042 ;
      RECT 3.942 6.818 4.266 6.862 ;
      RECT 3.942 6.368 4.266 6.412 ;
      RECT 3.942 3.668 4.266 3.712 ;
      RECT 3.942 3.218 4.266 3.262 ;
      RECT 3.942 3.038 4.266 3.082 ;
      RECT 3.942 2.588 4.266 2.632 ;
      RECT 3.942 2.408 4.266 2.452 ;
      RECT 3.942 1.958 4.266 2.002 ;
      RECT 3.942 1.778 4.266 1.822 ;
      RECT 3.942 1.328 4.266 1.372 ;
      RECT 3.942 1.148 4.266 1.192 ;
      RECT 3.942 0.698 4.266 0.742 ;
      RECT 3.942 0.518 4.266 0.562 ;
      RECT 3.942 0.068 4.266 0.112 ;
      RECT 4.394 9.608 4.462 9.922 ;
      RECT 4.394 8.978 4.462 9.292 ;
      RECT 4.394 8.348 4.462 8.662 ;
      RECT 4.394 7.718 4.462 8.032 ;
      RECT 4.394 7.088 4.462 7.402 ;
      RECT 4.394 6.458 4.462 6.772 ;
      RECT 4.394 5.828 4.462 6.142 ;
      RECT 4.394 3.938 4.462 4.252 ;
      RECT 4.394 3.308 4.462 3.622 ;
      RECT 4.394 2.678 4.462 2.992 ;
      RECT 4.394 2.048 4.462 2.362 ;
      RECT 4.394 1.418 4.462 1.732 ;
      RECT 4.394 0.788 4.462 1.102 ;
      RECT 4.394 0.158 4.462 0.472 ;
      RECT 4.502 9.608 4.57 9.922 ;
      RECT 4.502 8.978 4.57 9.292 ;
      RECT 4.502 8.348 4.57 8.662 ;
      RECT 4.502 7.718 4.57 8.032 ;
      RECT 4.502 7.088 4.57 7.402 ;
      RECT 4.502 6.458 4.57 6.772 ;
      RECT 4.502 5.828 4.57 6.142 ;
      RECT 4.502 3.938 4.57 4.252 ;
      RECT 4.502 3.308 4.57 3.622 ;
      RECT 4.502 2.678 4.57 2.992 ;
      RECT 4.502 2.048 4.57 2.362 ;
      RECT 4.502 1.418 4.57 1.732 ;
      RECT 4.502 0.788 4.57 1.102 ;
      RECT 4.502 0.158 4.57 0.472 ;
      RECT 4.61 9.608 4.678 9.922 ;
      RECT 4.61 8.978 4.678 9.292 ;
      RECT 4.61 8.348 4.678 8.662 ;
      RECT 4.61 7.718 4.678 8.032 ;
      RECT 4.61 7.088 4.678 7.402 ;
      RECT 4.61 6.458 4.678 6.772 ;
      RECT 4.61 5.828 4.678 6.142 ;
      RECT 4.61 3.938 4.678 4.252 ;
      RECT 4.61 3.308 4.678 3.622 ;
      RECT 4.61 2.678 4.678 2.992 ;
      RECT 4.61 2.048 4.678 2.362 ;
      RECT 4.61 1.418 4.678 1.732 ;
      RECT 4.61 0.788 4.678 1.102 ;
      RECT 4.61 0.158 4.678 0.472 ;
      RECT 4.374 9.968 4.698 10.012 ;
      RECT 4.374 9.518 4.698 9.562 ;
      RECT 4.374 9.338 4.698 9.382 ;
      RECT 4.374 8.888 4.698 8.932 ;
      RECT 4.374 8.708 4.698 8.752 ;
      RECT 4.374 8.258 4.698 8.302 ;
      RECT 4.374 8.078 4.698 8.122 ;
      RECT 4.374 7.628 4.698 7.672 ;
      RECT 4.374 7.448 4.698 7.492 ;
      RECT 4.374 6.998 4.698 7.042 ;
      RECT 4.374 6.818 4.698 6.862 ;
      RECT 4.374 6.368 4.698 6.412 ;
      RECT 4.374 6.188 4.698 6.232 ;
      RECT 4.374 5.738 4.698 5.782 ;
      RECT 4.374 4.298 4.698 4.342 ;
      RECT 4.374 3.848 4.698 3.892 ;
      RECT 4.374 3.668 4.698 3.712 ;
      RECT 4.374 3.218 4.698 3.262 ;
      RECT 4.374 3.038 4.698 3.082 ;
      RECT 4.374 2.588 4.698 2.632 ;
      RECT 4.374 2.408 4.698 2.452 ;
      RECT 4.374 1.958 4.698 2.002 ;
      RECT 4.374 1.778 4.698 1.822 ;
      RECT 4.374 1.328 4.698 1.372 ;
      RECT 4.374 1.148 4.698 1.192 ;
      RECT 4.374 0.698 4.698 0.742 ;
      RECT 4.374 0.518 4.698 0.562 ;
      RECT 4.374 0.068 4.698 0.112 ;
      RECT 4.826 9.608 4.894 9.922 ;
      RECT 4.826 8.978 4.894 9.292 ;
      RECT 4.826 8.348 4.894 8.662 ;
      RECT 4.826 7.718 4.894 8.032 ;
      RECT 4.826 7.088 4.894 7.402 ;
      RECT 4.826 6.458 4.894 6.772 ;
      RECT 4.826 5.828 4.894 6.142 ;
      RECT 4.826 3.938 4.894 4.252 ;
      RECT 4.826 3.308 4.894 3.622 ;
      RECT 4.826 2.678 4.894 2.992 ;
      RECT 4.826 2.048 4.894 2.362 ;
      RECT 4.826 1.418 4.894 1.732 ;
      RECT 4.826 0.788 4.894 1.102 ;
      RECT 4.826 0.158 4.894 0.472 ;
      RECT 4.934 9.608 5.002 9.922 ;
      RECT 4.934 8.978 5.002 9.292 ;
      RECT 4.934 8.348 5.002 8.662 ;
      RECT 4.934 7.718 5.002 8.032 ;
      RECT 4.934 7.088 5.002 7.402 ;
      RECT 4.934 6.458 5.002 6.772 ;
      RECT 4.934 5.828 5.002 6.142 ;
      RECT 4.934 3.938 5.002 4.252 ;
      RECT 4.934 3.308 5.002 3.622 ;
      RECT 4.934 2.678 5.002 2.992 ;
      RECT 4.934 2.048 5.002 2.362 ;
      RECT 4.934 1.418 5.002 1.732 ;
      RECT 4.934 0.788 5.002 1.102 ;
      RECT 4.934 0.158 5.002 0.472 ;
      RECT 5.042 9.608 5.11 9.922 ;
      RECT 5.042 8.978 5.11 9.292 ;
      RECT 5.042 8.348 5.11 8.662 ;
      RECT 5.042 7.718 5.11 8.032 ;
      RECT 5.042 7.088 5.11 7.402 ;
      RECT 5.042 6.458 5.11 6.772 ;
      RECT 5.042 5.828 5.11 6.142 ;
      RECT 5.042 5.468 5.11 5.602 ;
      RECT 5.042 5.108 5.11 5.242 ;
      RECT 5.042 4.838 5.11 4.972 ;
      RECT 5.042 4.478 5.11 4.612 ;
      RECT 5.042 3.938 5.11 4.252 ;
      RECT 5.042 3.308 5.11 3.622 ;
      RECT 5.042 2.678 5.11 2.992 ;
      RECT 5.042 2.048 5.11 2.362 ;
      RECT 5.042 1.418 5.11 1.732 ;
      RECT 5.042 0.788 5.11 1.102 ;
      RECT 5.042 0.158 5.11 0.472 ;
      RECT 4.806 9.968 5.13 10.012 ;
      RECT 4.806 9.518 5.13 9.562 ;
      RECT 4.806 9.338 5.13 9.382 ;
      RECT 4.806 8.888 5.13 8.932 ;
      RECT 4.806 8.708 5.13 8.752 ;
      RECT 4.806 8.258 5.13 8.302 ;
      RECT 4.806 8.078 5.13 8.122 ;
      RECT 4.806 7.628 5.13 7.672 ;
      RECT 4.806 7.448 5.13 7.492 ;
      RECT 4.806 6.998 5.13 7.042 ;
      RECT 4.806 6.818 5.13 6.862 ;
      RECT 4.806 6.368 5.13 6.412 ;
      RECT 4.806 6.188 5.13 6.232 ;
      RECT 4.806 5.738 5.13 5.782 ;
      RECT 4.806 4.298 5.13 4.342 ;
      RECT 4.806 3.848 5.13 3.892 ;
      RECT 4.806 3.668 5.13 3.712 ;
      RECT 4.806 3.218 5.13 3.262 ;
      RECT 4.806 3.038 5.13 3.082 ;
      RECT 4.806 2.588 5.13 2.632 ;
      RECT 4.806 2.408 5.13 2.452 ;
      RECT 4.806 1.958 5.13 2.002 ;
      RECT 4.806 1.778 5.13 1.822 ;
      RECT 4.806 1.328 5.13 1.372 ;
      RECT 4.806 1.148 5.13 1.192 ;
      RECT 4.806 0.698 5.13 0.742 ;
      RECT 4.806 0.518 5.13 0.562 ;
      RECT 4.806 0.068 5.13 0.112 ;
      RECT 5.258 9.608 5.326 9.922 ;
      RECT 5.258 8.978 5.326 9.292 ;
      RECT 5.258 8.348 5.326 8.662 ;
      RECT 5.258 7.718 5.326 8.032 ;
      RECT 5.258 7.088 5.326 7.402 ;
      RECT 5.258 6.458 5.326 6.772 ;
      RECT 5.258 5.828 5.326 6.142 ;
      RECT 5.258 5.468 5.326 5.602 ;
      RECT 5.258 5.108 5.326 5.242 ;
      RECT 5.258 4.838 5.326 4.972 ;
      RECT 5.258 4.478 5.326 4.612 ;
      RECT 5.258 3.938 5.326 4.252 ;
      RECT 5.258 3.308 5.326 3.622 ;
      RECT 5.258 2.678 5.326 2.992 ;
      RECT 5.258 2.048 5.326 2.362 ;
      RECT 5.258 1.418 5.326 1.732 ;
      RECT 5.258 0.788 5.326 1.102 ;
      RECT 5.258 0.158 5.326 0.472 ;
      RECT 5.366 9.608 5.434 9.922 ;
      RECT 5.366 8.978 5.434 9.292 ;
      RECT 5.366 8.348 5.434 8.662 ;
      RECT 5.366 7.718 5.434 8.032 ;
      RECT 5.366 7.088 5.434 7.402 ;
      RECT 5.366 6.458 5.434 6.772 ;
      RECT 5.366 6.008 5.434 6.142 ;
      RECT 5.366 5.828 5.434 5.962 ;
      RECT 5.366 4.118 5.434 4.252 ;
      RECT 5.366 3.938 5.434 4.072 ;
      RECT 5.366 3.308 5.434 3.622 ;
      RECT 5.366 2.678 5.434 2.992 ;
      RECT 5.366 2.048 5.434 2.362 ;
      RECT 5.366 1.418 5.434 1.732 ;
      RECT 5.366 0.788 5.434 1.102 ;
      RECT 5.366 0.158 5.434 0.472 ;
      RECT 5.474 9.608 5.542 9.922 ;
      RECT 5.474 8.978 5.542 9.292 ;
      RECT 5.474 8.348 5.542 8.662 ;
      RECT 5.474 7.718 5.542 8.032 ;
      RECT 5.474 7.088 5.542 7.402 ;
      RECT 5.474 6.458 5.542 6.772 ;
      RECT 5.474 5.828 5.542 6.142 ;
      RECT 5.474 3.938 5.542 4.252 ;
      RECT 5.474 3.308 5.542 3.622 ;
      RECT 5.474 2.678 5.542 2.992 ;
      RECT 5.474 2.048 5.542 2.362 ;
      RECT 5.474 1.418 5.542 1.732 ;
      RECT 5.474 0.788 5.542 1.102 ;
      RECT 5.474 0.158 5.542 0.472 ;
      RECT 5.238 9.968 5.562 10.012 ;
      RECT 5.238 9.518 5.562 9.562 ;
      RECT 5.238 9.338 5.562 9.382 ;
      RECT 5.238 8.888 5.562 8.932 ;
      RECT 5.238 8.708 5.562 8.752 ;
      RECT 5.238 8.258 5.562 8.302 ;
      RECT 5.238 8.078 5.562 8.122 ;
      RECT 5.238 7.628 5.562 7.672 ;
      RECT 5.238 7.448 5.562 7.492 ;
      RECT 5.238 6.998 5.562 7.042 ;
      RECT 5.238 6.818 5.562 6.862 ;
      RECT 5.238 6.368 5.562 6.412 ;
      RECT 5.238 3.668 5.562 3.712 ;
      RECT 5.238 3.218 5.562 3.262 ;
      RECT 5.238 3.038 5.562 3.082 ;
      RECT 5.238 2.588 5.562 2.632 ;
      RECT 5.238 2.408 5.562 2.452 ;
      RECT 5.238 1.958 5.562 2.002 ;
      RECT 5.238 1.778 5.562 1.822 ;
      RECT 5.238 1.328 5.562 1.372 ;
      RECT 5.238 1.148 5.562 1.192 ;
      RECT 5.238 0.698 5.562 0.742 ;
      RECT 5.238 0.518 5.562 0.562 ;
      RECT 5.238 0.068 5.562 0.112 ;
      RECT 5.582 5.828 5.65 6.142 ;
      RECT 5.582 3.938 5.65 4.252 ;
      RECT 5.69 9.608 5.758 9.922 ;
      RECT 5.69 8.978 5.758 9.292 ;
      RECT 5.69 8.348 5.758 8.662 ;
      RECT 5.69 7.718 5.758 8.032 ;
      RECT 5.69 7.088 5.758 7.402 ;
      RECT 5.69 6.458 5.758 6.772 ;
      RECT 5.69 6.008 5.758 6.142 ;
      RECT 5.69 5.828 5.758 5.962 ;
      RECT 5.69 5.198 5.758 5.512 ;
      RECT 5.69 4.568 5.758 4.882 ;
      RECT 5.69 4.118 5.758 4.252 ;
      RECT 5.69 3.938 5.758 4.072 ;
      RECT 5.69 3.308 5.758 3.622 ;
      RECT 5.69 2.678 5.758 2.992 ;
      RECT 5.69 2.048 5.758 2.362 ;
      RECT 5.69 1.418 5.758 1.732 ;
      RECT 5.69 0.788 5.758 1.102 ;
      RECT 5.69 0.158 5.758 0.472 ;
      RECT 5.798 9.608 5.866 9.922 ;
      RECT 5.798 8.978 5.866 9.292 ;
      RECT 5.798 8.348 5.866 8.662 ;
      RECT 5.798 7.718 5.866 8.032 ;
      RECT 5.798 7.088 5.866 7.402 ;
      RECT 5.798 6.638 5.866 6.772 ;
      RECT 5.798 6.458 5.866 6.592 ;
      RECT 5.798 5.198 5.866 5.512 ;
      RECT 5.798 4.568 5.866 4.882 ;
      RECT 5.798 3.488 5.866 3.622 ;
      RECT 5.798 3.308 5.866 3.442 ;
      RECT 5.798 2.678 5.866 2.992 ;
      RECT 5.798 2.048 5.866 2.362 ;
      RECT 5.798 1.418 5.866 1.732 ;
      RECT 5.798 0.788 5.866 1.102 ;
      RECT 5.798 0.158 5.866 0.472 ;
      RECT 5.906 9.608 5.974 9.922 ;
      RECT 5.906 8.978 5.974 9.292 ;
      RECT 5.906 8.348 5.974 8.662 ;
      RECT 5.906 7.718 5.974 8.032 ;
      RECT 5.906 7.088 5.974 7.402 ;
      RECT 5.906 6.458 5.974 6.772 ;
      RECT 5.906 6.008 5.974 6.142 ;
      RECT 5.906 5.828 5.974 5.962 ;
      RECT 5.906 5.198 5.974 5.512 ;
      RECT 5.906 4.568 5.974 4.882 ;
      RECT 5.906 4.118 5.974 4.252 ;
      RECT 5.906 3.938 5.974 4.072 ;
      RECT 5.906 3.308 5.974 3.622 ;
      RECT 5.906 2.678 5.974 2.992 ;
      RECT 5.906 2.048 5.974 2.362 ;
      RECT 5.906 1.418 5.974 1.732 ;
      RECT 5.906 0.788 5.974 1.102 ;
      RECT 5.906 0.158 5.974 0.472 ;
      RECT 5.67 9.968 5.994 10.012 ;
      RECT 5.67 9.518 5.994 9.562 ;
      RECT 5.67 9.338 5.994 9.382 ;
      RECT 5.67 8.888 5.994 8.932 ;
      RECT 5.67 8.708 5.994 8.752 ;
      RECT 5.67 8.258 5.994 8.302 ;
      RECT 5.67 8.078 5.994 8.122 ;
      RECT 5.67 7.628 5.994 7.672 ;
      RECT 5.67 7.448 5.994 7.492 ;
      RECT 5.67 6.998 5.994 7.042 ;
      RECT 5.67 5.558 5.994 5.602 ;
      RECT 5.67 5.108 5.994 5.152 ;
      RECT 5.67 4.928 5.994 4.972 ;
      RECT 5.67 4.478 5.994 4.522 ;
      RECT 5.67 3.038 5.994 3.082 ;
      RECT 5.67 2.588 5.994 2.632 ;
      RECT 5.67 2.408 5.994 2.452 ;
      RECT 5.67 1.958 5.994 2.002 ;
      RECT 5.67 1.778 5.994 1.822 ;
      RECT 5.67 1.328 5.994 1.372 ;
      RECT 5.67 1.148 5.994 1.192 ;
      RECT 5.67 0.698 5.994 0.742 ;
      RECT 5.67 0.518 5.994 0.562 ;
      RECT 5.67 0.068 5.994 0.112 ;
      RECT 6.014 6.458 6.082 6.772 ;
      RECT 6.014 5.828 6.082 6.142 ;
      RECT 6.014 3.938 6.082 4.252 ;
      RECT 6.014 3.308 6.082 3.622 ;
      RECT 6.122 9.608 6.19 9.922 ;
      RECT 6.122 8.978 6.19 9.292 ;
      RECT 6.122 8.348 6.19 8.662 ;
      RECT 6.122 7.718 6.19 8.032 ;
      RECT 6.122 7.088 6.19 7.402 ;
      RECT 6.122 6.638 6.19 6.772 ;
      RECT 6.122 6.458 6.19 6.592 ;
      RECT 6.122 5.828 6.19 6.142 ;
      RECT 6.122 5.198 6.19 5.512 ;
      RECT 6.122 4.568 6.19 4.882 ;
      RECT 6.122 3.938 6.19 4.252 ;
      RECT 6.122 3.488 6.19 3.622 ;
      RECT 6.122 3.308 6.19 3.442 ;
      RECT 6.122 2.678 6.19 2.992 ;
      RECT 6.122 2.048 6.19 2.362 ;
      RECT 6.122 1.418 6.19 1.732 ;
      RECT 6.122 0.788 6.19 1.102 ;
      RECT 6.122 0.158 6.19 0.472 ;
      RECT 6.23 9.608 6.298 9.922 ;
      RECT 6.23 8.978 6.298 9.292 ;
      RECT 6.23 8.348 6.298 8.662 ;
      RECT 6.23 7.718 6.298 8.032 ;
      RECT 6.23 7.268 6.298 7.402 ;
      RECT 6.23 7.088 6.298 7.222 ;
      RECT 6.23 6.008 6.298 6.142 ;
      RECT 6.23 5.828 6.298 5.962 ;
      RECT 6.23 5.198 6.298 5.512 ;
      RECT 6.23 4.568 6.298 4.882 ;
      RECT 6.23 4.118 6.298 4.252 ;
      RECT 6.23 3.938 6.298 4.072 ;
      RECT 6.23 2.858 6.298 2.992 ;
      RECT 6.23 2.678 6.298 2.812 ;
      RECT 6.23 2.048 6.298 2.362 ;
      RECT 6.23 1.418 6.298 1.732 ;
      RECT 6.23 0.788 6.298 1.102 ;
      RECT 6.23 0.158 6.298 0.472 ;
      RECT 6.338 9.608 6.406 9.922 ;
      RECT 6.338 8.978 6.406 9.292 ;
      RECT 6.338 8.348 6.406 8.662 ;
      RECT 6.338 7.718 6.406 8.032 ;
      RECT 6.338 7.088 6.406 7.402 ;
      RECT 6.338 6.638 6.406 6.772 ;
      RECT 6.338 6.458 6.406 6.592 ;
      RECT 6.338 5.828 6.406 6.142 ;
      RECT 6.338 5.198 6.406 5.512 ;
      RECT 6.338 4.568 6.406 4.882 ;
      RECT 6.338 3.938 6.406 4.252 ;
      RECT 6.338 3.488 6.406 3.622 ;
      RECT 6.338 3.308 6.406 3.442 ;
      RECT 6.338 2.678 6.406 2.992 ;
      RECT 6.338 2.048 6.406 2.362 ;
      RECT 6.338 1.418 6.406 1.732 ;
      RECT 6.338 0.788 6.406 1.102 ;
      RECT 6.338 0.158 6.406 0.472 ;
      RECT 6.102 9.968 6.426 10.012 ;
      RECT 6.102 9.518 6.426 9.562 ;
      RECT 6.102 9.338 6.426 9.382 ;
      RECT 6.102 8.888 6.426 8.932 ;
      RECT 6.102 8.708 6.426 8.752 ;
      RECT 6.102 8.258 6.426 8.302 ;
      RECT 6.102 8.078 6.426 8.122 ;
      RECT 6.102 7.628 6.426 7.672 ;
      RECT 6.102 5.558 6.426 5.602 ;
      RECT 6.102 5.108 6.426 5.152 ;
      RECT 6.102 4.928 6.426 4.972 ;
      RECT 6.102 4.478 6.426 4.522 ;
      RECT 6.102 2.408 6.426 2.452 ;
      RECT 6.102 1.958 6.426 2.002 ;
      RECT 6.102 1.778 6.426 1.822 ;
      RECT 6.102 1.328 6.426 1.372 ;
      RECT 6.102 1.148 6.426 1.192 ;
      RECT 6.102 0.698 6.426 0.742 ;
      RECT 6.102 0.518 6.426 0.562 ;
      RECT 6.102 0.068 6.426 0.112 ;
      RECT 6.446 7.088 6.514 7.402 ;
      RECT 6.446 6.458 6.514 6.772 ;
      RECT 6.446 3.308 6.514 3.622 ;
      RECT 6.446 2.678 6.514 2.992 ;
      RECT 6.554 9.608 6.622 9.922 ;
      RECT 6.554 8.978 6.622 9.292 ;
      RECT 6.554 8.348 6.622 8.662 ;
      RECT 6.554 7.718 6.622 8.032 ;
      RECT 6.554 7.268 6.622 7.402 ;
      RECT 6.554 7.088 6.622 7.222 ;
      RECT 6.554 6.458 6.622 6.772 ;
      RECT 6.554 5.828 6.622 6.142 ;
      RECT 6.554 5.198 6.622 5.512 ;
      RECT 6.554 4.568 6.622 4.882 ;
      RECT 6.554 3.938 6.622 4.252 ;
      RECT 6.554 3.308 6.622 3.622 ;
      RECT 6.554 2.858 6.622 2.992 ;
      RECT 6.554 2.678 6.622 2.812 ;
      RECT 6.554 2.048 6.622 2.362 ;
      RECT 6.554 1.418 6.622 1.732 ;
      RECT 6.554 0.788 6.622 1.102 ;
      RECT 6.554 0.158 6.622 0.472 ;
      RECT 6.662 9.608 6.73 9.922 ;
      RECT 6.662 8.978 6.73 9.292 ;
      RECT 6.662 8.348 6.73 8.662 ;
      RECT 6.662 7.898 6.73 8.032 ;
      RECT 6.662 7.718 6.73 7.852 ;
      RECT 6.662 6.638 6.73 6.772 ;
      RECT 6.662 6.458 6.73 6.592 ;
      RECT 6.662 5.828 6.73 6.142 ;
      RECT 6.662 5.198 6.73 5.512 ;
      RECT 6.662 4.568 6.73 4.882 ;
      RECT 6.662 3.938 6.73 4.252 ;
      RECT 6.662 3.488 6.73 3.622 ;
      RECT 6.662 3.308 6.73 3.442 ;
      RECT 6.662 2.228 6.73 2.362 ;
      RECT 6.662 2.048 6.73 2.182 ;
      RECT 6.662 1.418 6.73 1.732 ;
      RECT 6.662 0.788 6.73 1.102 ;
      RECT 6.662 0.158 6.73 0.472 ;
      RECT 6.77 9.608 6.838 9.922 ;
      RECT 6.77 8.978 6.838 9.292 ;
      RECT 6.77 8.348 6.838 8.662 ;
      RECT 6.77 7.718 6.838 8.032 ;
      RECT 6.77 7.268 6.838 7.402 ;
      RECT 6.77 7.088 6.838 7.222 ;
      RECT 6.77 6.458 6.838 6.772 ;
      RECT 6.77 5.828 6.838 6.142 ;
      RECT 6.77 5.198 6.838 5.512 ;
      RECT 6.77 4.568 6.838 4.882 ;
      RECT 6.77 3.938 6.838 4.252 ;
      RECT 6.77 3.308 6.838 3.622 ;
      RECT 6.77 2.858 6.838 2.992 ;
      RECT 6.77 2.678 6.838 2.812 ;
      RECT 6.77 2.048 6.838 2.362 ;
      RECT 6.77 1.418 6.838 1.732 ;
      RECT 6.77 0.788 6.838 1.102 ;
      RECT 6.77 0.158 6.838 0.472 ;
      RECT 6.534 9.968 6.858 10.012 ;
      RECT 6.534 9.518 6.858 9.562 ;
      RECT 6.534 9.338 6.858 9.382 ;
      RECT 6.534 8.888 6.858 8.932 ;
      RECT 6.534 8.708 6.858 8.752 ;
      RECT 6.534 8.258 6.858 8.302 ;
      RECT 6.534 6.188 6.858 6.232 ;
      RECT 6.534 5.738 6.858 5.782 ;
      RECT 6.534 5.558 6.858 5.602 ;
      RECT 6.534 5.108 6.858 5.152 ;
      RECT 6.534 4.928 6.858 4.972 ;
      RECT 6.534 4.478 6.858 4.522 ;
      RECT 6.534 4.298 6.858 4.342 ;
      RECT 6.534 3.848 6.858 3.892 ;
      RECT 6.534 1.778 6.858 1.822 ;
      RECT 6.534 1.328 6.858 1.372 ;
      RECT 6.534 1.148 6.858 1.192 ;
      RECT 6.534 0.698 6.858 0.742 ;
      RECT 6.534 0.518 6.858 0.562 ;
      RECT 6.534 0.068 6.858 0.112 ;
      RECT 6.878 7.718 6.946 8.032 ;
      RECT 6.878 7.088 6.946 7.402 ;
      RECT 6.878 2.678 6.946 2.992 ;
      RECT 6.878 2.048 6.946 2.362 ;
      RECT 6.986 9.608 7.054 9.922 ;
      RECT 6.986 8.978 7.054 9.292 ;
      RECT 6.986 8.348 7.054 8.662 ;
      RECT 6.986 7.898 7.054 8.032 ;
      RECT 6.986 7.718 7.054 7.852 ;
      RECT 6.986 7.088 7.054 7.402 ;
      RECT 6.986 6.458 7.054 6.772 ;
      RECT 6.986 5.828 7.054 6.142 ;
      RECT 6.986 5.198 7.054 5.512 ;
      RECT 6.986 4.568 7.054 4.882 ;
      RECT 6.986 3.938 7.054 4.252 ;
      RECT 6.986 3.308 7.054 3.622 ;
      RECT 6.986 2.678 7.054 2.992 ;
      RECT 6.986 2.228 7.054 2.362 ;
      RECT 6.986 2.048 7.054 2.182 ;
      RECT 6.986 1.418 7.054 1.732 ;
      RECT 6.986 0.788 7.054 1.102 ;
      RECT 6.986 0.158 7.054 0.472 ;
      RECT 7.094 9.608 7.162 9.922 ;
      RECT 7.094 8.978 7.162 9.292 ;
      RECT 7.094 8.528 7.162 8.662 ;
      RECT 7.094 8.348 7.162 8.482 ;
      RECT 7.094 7.268 7.162 7.402 ;
      RECT 7.094 7.088 7.162 7.222 ;
      RECT 7.094 6.458 7.162 6.772 ;
      RECT 7.094 5.828 7.162 6.142 ;
      RECT 7.094 5.198 7.162 5.512 ;
      RECT 7.094 4.568 7.162 4.882 ;
      RECT 7.094 3.938 7.162 4.252 ;
      RECT 7.094 3.308 7.162 3.622 ;
      RECT 7.094 2.858 7.162 2.992 ;
      RECT 7.094 2.678 7.162 2.812 ;
      RECT 7.094 1.598 7.162 1.732 ;
      RECT 7.094 1.418 7.162 1.552 ;
      RECT 7.094 0.788 7.162 1.102 ;
      RECT 7.094 0.158 7.162 0.472 ;
      RECT 7.202 9.608 7.27 9.922 ;
      RECT 7.202 8.978 7.27 9.292 ;
      RECT 7.202 8.348 7.27 8.662 ;
      RECT 7.202 7.898 7.27 8.032 ;
      RECT 7.202 7.718 7.27 7.852 ;
      RECT 7.202 7.088 7.27 7.402 ;
      RECT 7.202 6.458 7.27 6.772 ;
      RECT 7.202 5.828 7.27 6.142 ;
      RECT 7.202 5.198 7.27 5.512 ;
      RECT 7.202 4.568 7.27 4.882 ;
      RECT 7.202 3.938 7.27 4.252 ;
      RECT 7.202 3.308 7.27 3.622 ;
      RECT 7.202 2.678 7.27 2.992 ;
      RECT 7.202 2.228 7.27 2.362 ;
      RECT 7.202 2.048 7.27 2.182 ;
      RECT 7.202 1.418 7.27 1.732 ;
      RECT 7.202 0.788 7.27 1.102 ;
      RECT 7.202 0.158 7.27 0.472 ;
      RECT 6.966 9.968 7.29 10.012 ;
      RECT 6.966 9.518 7.29 9.562 ;
      RECT 6.966 9.338 7.29 9.382 ;
      RECT 6.966 8.888 7.29 8.932 ;
      RECT 6.966 6.818 7.29 6.862 ;
      RECT 6.966 6.368 7.29 6.412 ;
      RECT 6.966 6.188 7.29 6.232 ;
      RECT 6.966 5.738 7.29 5.782 ;
      RECT 6.966 5.558 7.29 5.602 ;
      RECT 6.966 5.108 7.29 5.152 ;
      RECT 6.966 4.928 7.29 4.972 ;
      RECT 6.966 4.478 7.29 4.522 ;
      RECT 6.966 4.298 7.29 4.342 ;
      RECT 6.966 3.848 7.29 3.892 ;
      RECT 6.966 3.668 7.29 3.712 ;
      RECT 6.966 3.218 7.29 3.262 ;
      RECT 6.966 1.148 7.29 1.192 ;
      RECT 6.966 0.698 7.29 0.742 ;
      RECT 6.966 0.518 7.29 0.562 ;
      RECT 6.966 0.068 7.29 0.112 ;
      RECT 7.31 8.348 7.378 8.662 ;
      RECT 7.31 7.718 7.378 8.032 ;
      RECT 7.31 2.048 7.378 2.362 ;
      RECT 7.31 1.418 7.378 1.732 ;
      RECT 7.418 9.608 7.486 9.922 ;
      RECT 7.418 8.978 7.486 9.292 ;
      RECT 7.418 8.528 7.486 8.662 ;
      RECT 7.418 8.348 7.486 8.482 ;
      RECT 7.418 7.718 7.486 8.032 ;
      RECT 7.418 7.088 7.486 7.402 ;
      RECT 7.418 6.458 7.486 6.772 ;
      RECT 7.418 5.828 7.486 6.142 ;
      RECT 7.418 5.198 7.486 5.512 ;
      RECT 7.418 4.568 7.486 4.882 ;
      RECT 7.418 3.938 7.486 4.252 ;
      RECT 7.418 3.308 7.486 3.622 ;
      RECT 7.418 2.678 7.486 2.992 ;
      RECT 7.418 2.048 7.486 2.362 ;
      RECT 7.418 1.598 7.486 1.732 ;
      RECT 7.418 1.418 7.486 1.552 ;
      RECT 7.418 0.788 7.486 1.102 ;
      RECT 7.418 0.158 7.486 0.472 ;
      RECT 7.526 9.608 7.594 9.922 ;
      RECT 7.526 9.158 7.594 9.292 ;
      RECT 7.526 8.978 7.594 9.112 ;
      RECT 7.526 7.898 7.594 8.032 ;
      RECT 7.526 7.718 7.594 7.852 ;
      RECT 7.526 7.088 7.594 7.402 ;
      RECT 7.526 6.458 7.594 6.772 ;
      RECT 7.526 5.828 7.594 6.142 ;
      RECT 7.526 5.198 7.594 5.512 ;
      RECT 7.526 4.568 7.594 4.882 ;
      RECT 7.526 3.938 7.594 4.252 ;
      RECT 7.526 3.308 7.594 3.622 ;
      RECT 7.526 2.678 7.594 2.992 ;
      RECT 7.526 2.228 7.594 2.362 ;
      RECT 7.526 2.048 7.594 2.182 ;
      RECT 7.526 0.968 7.594 1.102 ;
      RECT 7.526 0.788 7.594 0.922 ;
      RECT 7.526 0.158 7.594 0.472 ;
      RECT 7.634 9.608 7.702 9.922 ;
      RECT 7.634 8.978 7.702 9.292 ;
      RECT 7.634 8.528 7.702 8.662 ;
      RECT 7.634 8.348 7.702 8.482 ;
      RECT 7.634 7.718 7.702 8.032 ;
      RECT 7.634 7.088 7.702 7.402 ;
      RECT 7.634 6.458 7.702 6.772 ;
      RECT 7.634 5.828 7.702 6.142 ;
      RECT 7.634 5.198 7.702 5.512 ;
      RECT 7.634 4.568 7.702 4.882 ;
      RECT 7.634 3.938 7.702 4.252 ;
      RECT 7.634 3.308 7.702 3.622 ;
      RECT 7.634 2.678 7.702 2.992 ;
      RECT 7.634 2.048 7.702 2.362 ;
      RECT 7.634 1.598 7.702 1.732 ;
      RECT 7.634 1.418 7.702 1.552 ;
      RECT 7.634 0.788 7.702 1.102 ;
      RECT 7.634 0.158 7.702 0.472 ;
      RECT 7.398 9.968 7.722 10.012 ;
      RECT 7.398 9.518 7.722 9.562 ;
      RECT 7.398 7.448 7.722 7.492 ;
      RECT 7.398 6.998 7.722 7.042 ;
      RECT 7.398 6.818 7.722 6.862 ;
      RECT 7.398 6.368 7.722 6.412 ;
      RECT 7.398 6.188 7.722 6.232 ;
      RECT 7.398 5.738 7.722 5.782 ;
      RECT 7.398 5.558 7.722 5.602 ;
      RECT 7.398 5.108 7.722 5.152 ;
      RECT 7.398 4.928 7.722 4.972 ;
      RECT 7.398 4.478 7.722 4.522 ;
      RECT 7.398 4.298 7.722 4.342 ;
      RECT 7.398 3.848 7.722 3.892 ;
      RECT 7.398 3.668 7.722 3.712 ;
      RECT 7.398 3.218 7.722 3.262 ;
      RECT 7.398 3.038 7.722 3.082 ;
      RECT 7.398 2.588 7.722 2.632 ;
      RECT 7.398 0.518 7.722 0.562 ;
      RECT 7.398 0.068 7.722 0.112 ;
      RECT 7.742 8.978 7.81 9.292 ;
      RECT 7.742 8.348 7.81 8.662 ;
      RECT 7.742 1.418 7.81 1.732 ;
      RECT 7.742 0.788 7.81 1.102 ;
      RECT 7.85 9.608 7.918 9.922 ;
      RECT 7.85 9.158 7.918 9.292 ;
      RECT 7.85 8.978 7.918 9.112 ;
      RECT 7.85 8.348 7.918 8.662 ;
      RECT 7.85 7.718 7.918 8.032 ;
      RECT 7.85 7.088 7.918 7.402 ;
      RECT 7.85 6.458 7.918 6.772 ;
      RECT 7.85 5.828 7.918 6.142 ;
      RECT 7.85 5.198 7.918 5.512 ;
      RECT 7.85 4.568 7.918 4.882 ;
      RECT 7.85 3.938 7.918 4.252 ;
      RECT 7.85 3.308 7.918 3.622 ;
      RECT 7.85 2.678 7.918 2.992 ;
      RECT 7.85 2.048 7.918 2.362 ;
      RECT 7.85 1.418 7.918 1.732 ;
      RECT 7.85 0.968 7.918 1.102 ;
      RECT 7.85 0.788 7.918 0.922 ;
      RECT 7.85 0.158 7.918 0.472 ;
      RECT 7.958 9.608 8.026 9.922 ;
      RECT 7.958 8.528 8.026 8.662 ;
      RECT 7.958 8.348 8.026 8.482 ;
      RECT 7.958 7.718 8.026 8.032 ;
      RECT 7.958 7.088 8.026 7.402 ;
      RECT 7.958 6.458 8.026 6.772 ;
      RECT 7.958 5.828 8.026 6.142 ;
      RECT 7.958 5.198 8.026 5.512 ;
      RECT 7.958 4.568 8.026 4.882 ;
      RECT 7.958 3.938 8.026 4.252 ;
      RECT 7.958 3.308 8.026 3.622 ;
      RECT 7.958 2.678 8.026 2.992 ;
      RECT 7.958 2.048 8.026 2.362 ;
      RECT 7.958 1.598 8.026 1.732 ;
      RECT 7.958 1.418 8.026 1.552 ;
      RECT 7.958 0.158 8.026 0.472 ;
      RECT 8.066 9.608 8.134 9.922 ;
      RECT 8.066 9.158 8.134 9.292 ;
      RECT 8.066 8.978 8.134 9.112 ;
      RECT 8.066 8.348 8.134 8.662 ;
      RECT 8.066 7.718 8.134 8.032 ;
      RECT 8.066 7.088 8.134 7.402 ;
      RECT 8.066 6.458 8.134 6.772 ;
      RECT 8.066 5.828 8.134 6.142 ;
      RECT 8.066 5.198 8.134 5.512 ;
      RECT 8.066 4.568 8.134 4.882 ;
      RECT 8.066 3.938 8.134 4.252 ;
      RECT 8.066 3.308 8.134 3.622 ;
      RECT 8.066 2.678 8.134 2.992 ;
      RECT 8.066 2.048 8.134 2.362 ;
      RECT 8.066 1.418 8.134 1.732 ;
      RECT 8.066 0.968 8.134 1.102 ;
      RECT 8.066 0.788 8.134 0.922 ;
      RECT 8.066 0.158 8.134 0.472 ;
      RECT 7.83 9.968 8.154 10.012 ;
      RECT 7.83 9.518 8.154 9.562 ;
      RECT 7.83 8.078 8.154 8.122 ;
      RECT 7.83 7.628 8.154 7.672 ;
      RECT 7.83 7.448 8.154 7.492 ;
      RECT 7.83 6.998 8.154 7.042 ;
      RECT 7.83 6.818 8.154 6.862 ;
      RECT 7.83 6.368 8.154 6.412 ;
      RECT 7.83 6.188 8.154 6.232 ;
      RECT 7.83 5.738 8.154 5.782 ;
      RECT 7.83 5.558 8.154 5.602 ;
      RECT 7.83 5.108 8.154 5.152 ;
      RECT 7.83 4.928 8.154 4.972 ;
      RECT 7.83 4.478 8.154 4.522 ;
      RECT 7.83 4.298 8.154 4.342 ;
      RECT 7.83 3.848 8.154 3.892 ;
      RECT 7.83 3.668 8.154 3.712 ;
      RECT 7.83 3.218 8.154 3.262 ;
      RECT 7.83 3.038 8.154 3.082 ;
      RECT 7.83 2.588 8.154 2.632 ;
      RECT 7.83 2.408 8.154 2.452 ;
      RECT 7.83 1.958 8.154 2.002 ;
      RECT 7.83 0.518 8.154 0.562 ;
      RECT 7.83 0.068 8.154 0.112 ;
      RECT 8.174 8.978 8.242 9.292 ;
      RECT 8.174 0.788 8.242 1.102 ;
      RECT 8.282 9.608 8.35 9.922 ;
      RECT 8.282 8.978 8.35 9.292 ;
      RECT 8.282 8.348 8.35 8.662 ;
      RECT 8.282 7.718 8.35 8.032 ;
      RECT 8.282 7.088 8.35 7.402 ;
      RECT 8.282 6.458 8.35 6.772 ;
      RECT 8.282 5.828 8.35 6.142 ;
      RECT 8.282 5.198 8.35 5.512 ;
      RECT 8.282 4.568 8.35 4.882 ;
      RECT 8.282 3.938 8.35 4.252 ;
      RECT 8.282 3.308 8.35 3.622 ;
      RECT 8.282 2.678 8.35 2.992 ;
      RECT 8.282 2.048 8.35 2.362 ;
      RECT 8.282 1.418 8.35 1.732 ;
      RECT 8.282 0.788 8.35 1.102 ;
      RECT 8.282 0.158 8.35 0.472 ;
      RECT 8.39 9.608 8.458 9.922 ;
      RECT 8.39 9.158 8.458 9.292 ;
      RECT 8.39 8.978 8.458 9.112 ;
      RECT 8.39 8.348 8.458 8.662 ;
      RECT 8.39 7.718 8.458 8.032 ;
      RECT 8.39 7.088 8.458 7.402 ;
      RECT 8.39 6.458 8.458 6.772 ;
      RECT 8.39 5.828 8.458 6.142 ;
      RECT 8.39 5.198 8.458 5.512 ;
      RECT 8.39 4.568 8.458 4.882 ;
      RECT 8.39 3.938 8.458 4.252 ;
      RECT 8.39 3.308 8.458 3.622 ;
      RECT 8.39 2.678 8.458 2.992 ;
      RECT 8.39 2.048 8.458 2.362 ;
      RECT 8.39 1.418 8.458 1.732 ;
      RECT 8.39 0.968 8.458 1.102 ;
      RECT 8.39 0.788 8.458 0.922 ;
      RECT 8.39 0.158 8.458 0.472 ;
      RECT 8.498 9.608 8.566 9.922 ;
      RECT 8.498 8.978 8.566 9.292 ;
      RECT 8.498 8.348 8.566 8.662 ;
      RECT 8.498 7.718 8.566 8.032 ;
      RECT 8.498 7.088 8.566 7.402 ;
      RECT 8.498 6.458 8.566 6.772 ;
      RECT 8.498 5.828 8.566 6.142 ;
      RECT 8.498 5.198 8.566 5.512 ;
      RECT 8.498 4.568 8.566 4.882 ;
      RECT 8.498 3.938 8.566 4.252 ;
      RECT 8.498 3.308 8.566 3.622 ;
      RECT 8.498 2.678 8.566 2.992 ;
      RECT 8.498 2.048 8.566 2.362 ;
      RECT 8.498 1.418 8.566 1.732 ;
      RECT 8.498 0.788 8.566 1.102 ;
      RECT 8.498 0.158 8.566 0.472 ;
      RECT 8.262 9.968 8.586 10.012 ;
      RECT 8.262 9.518 8.586 9.562 ;
      RECT 8.262 8.708 8.586 8.752 ;
      RECT 8.262 8.258 8.586 8.302 ;
      RECT 8.262 8.078 8.586 8.122 ;
      RECT 8.262 7.628 8.586 7.672 ;
      RECT 8.262 7.448 8.586 7.492 ;
      RECT 8.262 6.998 8.586 7.042 ;
      RECT 8.262 6.818 8.586 6.862 ;
      RECT 8.262 6.368 8.586 6.412 ;
      RECT 8.262 6.188 8.586 6.232 ;
      RECT 8.262 5.738 8.586 5.782 ;
      RECT 8.262 5.558 8.586 5.602 ;
      RECT 8.262 5.108 8.586 5.152 ;
      RECT 8.262 4.928 8.586 4.972 ;
      RECT 8.262 4.478 8.586 4.522 ;
      RECT 8.262 4.298 8.586 4.342 ;
      RECT 8.262 3.848 8.586 3.892 ;
      RECT 8.262 3.668 8.586 3.712 ;
      RECT 8.262 3.218 8.586 3.262 ;
      RECT 8.262 3.038 8.586 3.082 ;
      RECT 8.262 2.588 8.586 2.632 ;
      RECT 8.262 2.408 8.586 2.452 ;
      RECT 8.262 1.958 8.586 2.002 ;
      RECT 8.262 1.778 8.586 1.822 ;
      RECT 8.262 1.328 8.586 1.372 ;
      RECT 8.262 0.518 8.586 0.562 ;
      RECT 8.262 0.068 8.586 0.112 ;
      RECT 8.714 9.608 8.782 9.922 ;
      RECT 8.714 8.978 8.782 9.292 ;
      RECT 8.714 8.348 8.782 8.662 ;
      RECT 8.714 7.718 8.782 8.032 ;
      RECT 8.714 7.088 8.782 7.402 ;
      RECT 8.714 6.458 8.782 6.772 ;
      RECT 8.714 5.828 8.782 6.142 ;
      RECT 8.714 5.198 8.782 5.512 ;
      RECT 8.714 4.568 8.782 4.882 ;
      RECT 8.714 3.938 8.782 4.252 ;
      RECT 8.714 3.308 8.782 3.622 ;
      RECT 8.714 2.678 8.782 2.992 ;
      RECT 8.714 2.048 8.782 2.362 ;
      RECT 8.714 1.418 8.782 1.732 ;
      RECT 8.714 0.788 8.782 1.102 ;
      RECT 8.714 0.158 8.782 0.472 ;
      RECT 8.822 9.608 8.89 9.922 ;
      RECT 8.822 8.978 8.89 9.292 ;
      RECT 8.822 8.348 8.89 8.662 ;
      RECT 8.822 7.718 8.89 8.032 ;
      RECT 8.822 7.088 8.89 7.402 ;
      RECT 8.822 6.458 8.89 6.772 ;
      RECT 8.822 5.828 8.89 6.142 ;
      RECT 8.822 5.198 8.89 5.512 ;
      RECT 8.822 4.568 8.89 4.882 ;
      RECT 8.822 3.938 8.89 4.252 ;
      RECT 8.822 3.308 8.89 3.622 ;
      RECT 8.822 2.678 8.89 2.992 ;
      RECT 8.822 2.048 8.89 2.362 ;
      RECT 8.822 1.418 8.89 1.732 ;
      RECT 8.822 0.788 8.89 1.102 ;
      RECT 8.822 0.158 8.89 0.472 ;
      RECT 8.93 9.608 8.998 9.922 ;
      RECT 8.93 8.978 8.998 9.292 ;
      RECT 8.93 8.348 8.998 8.662 ;
      RECT 8.93 7.718 8.998 8.032 ;
      RECT 8.93 7.088 8.998 7.402 ;
      RECT 8.93 6.458 8.998 6.772 ;
      RECT 8.93 5.828 8.998 6.142 ;
      RECT 8.93 5.198 8.998 5.512 ;
      RECT 8.93 4.568 8.998 4.882 ;
      RECT 8.93 3.938 8.998 4.252 ;
      RECT 8.93 3.308 8.998 3.622 ;
      RECT 8.93 2.678 8.998 2.992 ;
      RECT 8.93 2.048 8.998 2.362 ;
      RECT 8.93 1.418 8.998 1.732 ;
      RECT 8.93 0.788 8.998 1.102 ;
      RECT 8.93 0.158 8.998 0.472 ;
      RECT 8.694 9.968 9.018 10.012 ;
      RECT 8.694 9.518 9.018 9.562 ;
      RECT 8.694 9.338 9.018 9.382 ;
      RECT 8.694 8.888 9.018 8.932 ;
      RECT 8.694 8.708 9.018 8.752 ;
      RECT 8.694 8.258 9.018 8.302 ;
      RECT 8.694 8.078 9.018 8.122 ;
      RECT 8.694 7.628 9.018 7.672 ;
      RECT 8.694 7.448 9.018 7.492 ;
      RECT 8.694 6.998 9.018 7.042 ;
      RECT 8.694 6.818 9.018 6.862 ;
      RECT 8.694 6.368 9.018 6.412 ;
      RECT 8.694 6.188 9.018 6.232 ;
      RECT 8.694 5.738 9.018 5.782 ;
      RECT 8.694 5.558 9.018 5.602 ;
      RECT 8.694 5.108 9.018 5.152 ;
      RECT 8.694 4.928 9.018 4.972 ;
      RECT 8.694 4.478 9.018 4.522 ;
      RECT 8.694 4.298 9.018 4.342 ;
      RECT 8.694 3.848 9.018 3.892 ;
      RECT 8.694 3.668 9.018 3.712 ;
      RECT 8.694 3.218 9.018 3.262 ;
      RECT 8.694 3.038 9.018 3.082 ;
      RECT 8.694 2.588 9.018 2.632 ;
      RECT 8.694 2.408 9.018 2.452 ;
      RECT 8.694 1.958 9.018 2.002 ;
      RECT 8.694 1.778 9.018 1.822 ;
      RECT 8.694 1.328 9.018 1.372 ;
      RECT 8.694 1.148 9.018 1.192 ;
      RECT 8.694 0.698 9.018 0.742 ;
      RECT 8.694 0.518 9.018 0.562 ;
      RECT 8.694 0.068 9.018 0.112 ;
      RECT 9.146 9.608 9.214 9.922 ;
      RECT 9.146 8.978 9.214 9.292 ;
      RECT 9.146 8.348 9.214 8.662 ;
      RECT 9.146 7.718 9.214 8.032 ;
      RECT 9.146 7.088 9.214 7.402 ;
      RECT 9.146 6.458 9.214 6.772 ;
      RECT 9.146 5.828 9.214 6.142 ;
      RECT 9.146 5.198 9.214 5.512 ;
      RECT 9.146 4.568 9.214 4.882 ;
      RECT 9.146 3.938 9.214 4.252 ;
      RECT 9.146 3.308 9.214 3.622 ;
      RECT 9.146 2.678 9.214 2.992 ;
      RECT 9.146 2.048 9.214 2.362 ;
      RECT 9.146 1.418 9.214 1.732 ;
      RECT 9.146 0.788 9.214 1.102 ;
      RECT 9.146 0.158 9.214 0.472 ;
      RECT 9.254 9.608 9.322 9.922 ;
      RECT 9.254 8.978 9.322 9.292 ;
      RECT 9.254 8.348 9.322 8.662 ;
      RECT 9.254 7.718 9.322 8.032 ;
      RECT 9.254 7.088 9.322 7.402 ;
      RECT 9.254 6.458 9.322 6.772 ;
      RECT 9.254 5.828 9.322 6.142 ;
      RECT 9.254 5.198 9.322 5.512 ;
      RECT 9.254 4.568 9.322 4.882 ;
      RECT 9.254 3.938 9.322 4.252 ;
      RECT 9.254 3.308 9.322 3.622 ;
      RECT 9.254 2.678 9.322 2.992 ;
      RECT 9.254 2.048 9.322 2.362 ;
      RECT 9.254 1.418 9.322 1.732 ;
      RECT 9.254 0.788 9.322 1.102 ;
      RECT 9.254 0.158 9.322 0.472 ;
      RECT 9.362 9.608 9.43 9.922 ;
      RECT 9.362 8.978 9.43 9.292 ;
      RECT 9.362 8.348 9.43 8.662 ;
      RECT 9.362 7.718 9.43 8.032 ;
      RECT 9.362 7.088 9.43 7.402 ;
      RECT 9.362 6.458 9.43 6.772 ;
      RECT 9.362 5.828 9.43 6.142 ;
      RECT 9.362 5.198 9.43 5.512 ;
      RECT 9.362 4.568 9.43 4.882 ;
      RECT 9.362 3.938 9.43 4.252 ;
      RECT 9.362 3.308 9.43 3.622 ;
      RECT 9.362 2.678 9.43 2.992 ;
      RECT 9.362 2.048 9.43 2.362 ;
      RECT 9.362 1.418 9.43 1.732 ;
      RECT 9.362 0.788 9.43 1.102 ;
      RECT 9.362 0.158 9.43 0.472 ;
      RECT 9.126 9.968 9.45 10.012 ;
      RECT 9.126 9.518 9.45 9.562 ;
      RECT 9.126 9.338 9.45 9.382 ;
      RECT 9.126 8.888 9.45 8.932 ;
      RECT 9.126 8.708 9.45 8.752 ;
      RECT 9.126 8.258 9.45 8.302 ;
      RECT 9.126 8.078 9.45 8.122 ;
      RECT 9.126 7.628 9.45 7.672 ;
      RECT 9.126 7.448 9.45 7.492 ;
      RECT 9.126 6.998 9.45 7.042 ;
      RECT 9.126 6.818 9.45 6.862 ;
      RECT 9.126 6.368 9.45 6.412 ;
      RECT 9.126 6.188 9.45 6.232 ;
      RECT 9.126 5.738 9.45 5.782 ;
      RECT 9.126 5.558 9.45 5.602 ;
      RECT 9.126 5.108 9.45 5.152 ;
      RECT 9.126 4.928 9.45 4.972 ;
      RECT 9.126 4.478 9.45 4.522 ;
      RECT 9.126 4.298 9.45 4.342 ;
      RECT 9.126 3.848 9.45 3.892 ;
      RECT 9.126 3.668 9.45 3.712 ;
      RECT 9.126 3.218 9.45 3.262 ;
      RECT 9.126 3.038 9.45 3.082 ;
      RECT 9.126 2.588 9.45 2.632 ;
      RECT 9.126 2.408 9.45 2.452 ;
      RECT 9.126 1.958 9.45 2.002 ;
      RECT 9.126 1.778 9.45 1.822 ;
      RECT 9.126 1.328 9.45 1.372 ;
      RECT 9.126 1.148 9.45 1.192 ;
      RECT 9.126 0.698 9.45 0.742 ;
      RECT 9.126 0.518 9.45 0.562 ;
      RECT 9.126 0.068 9.45 0.112 ;
    LAYER v0 ;
      RECT 9.362 0.068 9.43 0.112 ;
      RECT 9.362 0.518 9.43 0.562 ;
      RECT 9.362 0.698 9.43 0.742 ;
      RECT 9.362 1.148 9.43 1.192 ;
      RECT 9.362 1.328 9.43 1.372 ;
      RECT 9.362 1.778 9.43 1.822 ;
      RECT 9.362 1.958 9.43 2.002 ;
      RECT 9.362 2.408 9.43 2.452 ;
      RECT 9.362 2.588 9.43 2.632 ;
      RECT 9.362 3.038 9.43 3.082 ;
      RECT 9.362 3.218 9.43 3.262 ;
      RECT 9.362 3.668 9.43 3.712 ;
      RECT 9.362 3.848 9.43 3.892 ;
      RECT 9.362 4.298 9.43 4.342 ;
      RECT 9.362 4.478 9.43 4.522 ;
      RECT 9.362 4.928 9.43 4.972 ;
      RECT 9.362 5.108 9.43 5.152 ;
      RECT 9.362 5.558 9.43 5.602 ;
      RECT 9.362 5.738 9.43 5.782 ;
      RECT 9.362 6.188 9.43 6.232 ;
      RECT 9.362 6.368 9.43 6.412 ;
      RECT 9.362 6.818 9.43 6.862 ;
      RECT 9.362 6.998 9.43 7.042 ;
      RECT 9.362 7.448 9.43 7.492 ;
      RECT 9.362 7.628 9.43 7.672 ;
      RECT 9.362 8.078 9.43 8.122 ;
      RECT 9.362 8.258 9.43 8.302 ;
      RECT 9.362 8.708 9.43 8.752 ;
      RECT 9.362 8.888 9.43 8.932 ;
      RECT 9.362 9.338 9.43 9.382 ;
      RECT 9.362 9.518 9.43 9.562 ;
      RECT 9.362 9.968 9.43 10.012 ;
      RECT 9.146 0.068 9.214 0.112 ;
      RECT 9.146 0.518 9.214 0.562 ;
      RECT 9.146 0.698 9.214 0.742 ;
      RECT 9.146 1.148 9.214 1.192 ;
      RECT 9.146 1.328 9.214 1.372 ;
      RECT 9.146 1.778 9.214 1.822 ;
      RECT 9.146 1.958 9.214 2.002 ;
      RECT 9.146 2.408 9.214 2.452 ;
      RECT 9.146 2.588 9.214 2.632 ;
      RECT 9.146 3.038 9.214 3.082 ;
      RECT 9.146 3.218 9.214 3.262 ;
      RECT 9.146 3.668 9.214 3.712 ;
      RECT 9.146 3.848 9.214 3.892 ;
      RECT 9.146 4.298 9.214 4.342 ;
      RECT 9.146 4.478 9.214 4.522 ;
      RECT 9.146 4.928 9.214 4.972 ;
      RECT 9.146 5.108 9.214 5.152 ;
      RECT 9.146 5.558 9.214 5.602 ;
      RECT 9.146 5.738 9.214 5.782 ;
      RECT 9.146 6.188 9.214 6.232 ;
      RECT 9.146 6.368 9.214 6.412 ;
      RECT 9.146 6.818 9.214 6.862 ;
      RECT 9.146 6.998 9.214 7.042 ;
      RECT 9.146 7.448 9.214 7.492 ;
      RECT 9.146 7.628 9.214 7.672 ;
      RECT 9.146 8.078 9.214 8.122 ;
      RECT 9.146 8.258 9.214 8.302 ;
      RECT 9.146 8.708 9.214 8.752 ;
      RECT 9.146 8.888 9.214 8.932 ;
      RECT 9.146 9.338 9.214 9.382 ;
      RECT 9.146 9.518 9.214 9.562 ;
      RECT 9.146 9.968 9.214 10.012 ;
      RECT 8.93 0.068 8.998 0.112 ;
      RECT 8.93 0.518 8.998 0.562 ;
      RECT 8.93 0.698 8.998 0.742 ;
      RECT 8.93 1.148 8.998 1.192 ;
      RECT 8.93 1.328 8.998 1.372 ;
      RECT 8.93 1.778 8.998 1.822 ;
      RECT 8.93 1.958 8.998 2.002 ;
      RECT 8.93 2.408 8.998 2.452 ;
      RECT 8.93 2.588 8.998 2.632 ;
      RECT 8.93 3.038 8.998 3.082 ;
      RECT 8.93 3.218 8.998 3.262 ;
      RECT 8.93 3.668 8.998 3.712 ;
      RECT 8.93 3.848 8.998 3.892 ;
      RECT 8.93 4.298 8.998 4.342 ;
      RECT 8.93 4.478 8.998 4.522 ;
      RECT 8.93 4.928 8.998 4.972 ;
      RECT 8.93 5.108 8.998 5.152 ;
      RECT 8.93 5.558 8.998 5.602 ;
      RECT 8.93 5.738 8.998 5.782 ;
      RECT 8.93 6.188 8.998 6.232 ;
      RECT 8.93 6.368 8.998 6.412 ;
      RECT 8.93 6.818 8.998 6.862 ;
      RECT 8.93 6.998 8.998 7.042 ;
      RECT 8.93 7.448 8.998 7.492 ;
      RECT 8.93 7.628 8.998 7.672 ;
      RECT 8.93 8.078 8.998 8.122 ;
      RECT 8.93 8.258 8.998 8.302 ;
      RECT 8.93 8.708 8.998 8.752 ;
      RECT 8.93 8.888 8.998 8.932 ;
      RECT 8.93 9.338 8.998 9.382 ;
      RECT 8.93 9.518 8.998 9.562 ;
      RECT 8.93 9.968 8.998 10.012 ;
      RECT 8.714 0.068 8.782 0.112 ;
      RECT 8.714 0.518 8.782 0.562 ;
      RECT 8.714 0.698 8.782 0.742 ;
      RECT 8.714 1.148 8.782 1.192 ;
      RECT 8.714 1.328 8.782 1.372 ;
      RECT 8.714 1.778 8.782 1.822 ;
      RECT 8.714 1.958 8.782 2.002 ;
      RECT 8.714 2.408 8.782 2.452 ;
      RECT 8.714 2.588 8.782 2.632 ;
      RECT 8.714 3.038 8.782 3.082 ;
      RECT 8.714 3.218 8.782 3.262 ;
      RECT 8.714 3.668 8.782 3.712 ;
      RECT 8.714 3.848 8.782 3.892 ;
      RECT 8.714 4.298 8.782 4.342 ;
      RECT 8.714 4.478 8.782 4.522 ;
      RECT 8.714 4.928 8.782 4.972 ;
      RECT 8.714 5.108 8.782 5.152 ;
      RECT 8.714 5.558 8.782 5.602 ;
      RECT 8.714 5.738 8.782 5.782 ;
      RECT 8.714 6.188 8.782 6.232 ;
      RECT 8.714 6.368 8.782 6.412 ;
      RECT 8.714 6.818 8.782 6.862 ;
      RECT 8.714 6.998 8.782 7.042 ;
      RECT 8.714 7.448 8.782 7.492 ;
      RECT 8.714 7.628 8.782 7.672 ;
      RECT 8.714 8.078 8.782 8.122 ;
      RECT 8.714 8.258 8.782 8.302 ;
      RECT 8.714 8.708 8.782 8.752 ;
      RECT 8.714 8.888 8.782 8.932 ;
      RECT 8.714 9.338 8.782 9.382 ;
      RECT 8.714 9.518 8.782 9.562 ;
      RECT 8.714 9.968 8.782 10.012 ;
      RECT 8.498 0.068 8.566 0.112 ;
      RECT 8.498 0.518 8.566 0.562 ;
      RECT 8.498 1.328 8.566 1.372 ;
      RECT 8.498 1.778 8.566 1.822 ;
      RECT 8.498 1.958 8.566 2.002 ;
      RECT 8.498 2.408 8.566 2.452 ;
      RECT 8.498 2.588 8.566 2.632 ;
      RECT 8.498 3.038 8.566 3.082 ;
      RECT 8.498 3.218 8.566 3.262 ;
      RECT 8.498 3.668 8.566 3.712 ;
      RECT 8.498 3.848 8.566 3.892 ;
      RECT 8.498 4.298 8.566 4.342 ;
      RECT 8.498 4.478 8.566 4.522 ;
      RECT 8.498 4.928 8.566 4.972 ;
      RECT 8.498 5.108 8.566 5.152 ;
      RECT 8.498 5.558 8.566 5.602 ;
      RECT 8.498 5.738 8.566 5.782 ;
      RECT 8.498 6.188 8.566 6.232 ;
      RECT 8.498 6.368 8.566 6.412 ;
      RECT 8.498 6.818 8.566 6.862 ;
      RECT 8.498 6.998 8.566 7.042 ;
      RECT 8.498 7.448 8.566 7.492 ;
      RECT 8.498 7.628 8.566 7.672 ;
      RECT 8.498 8.078 8.566 8.122 ;
      RECT 8.498 8.258 8.566 8.302 ;
      RECT 8.498 8.708 8.566 8.752 ;
      RECT 8.498 9.518 8.566 9.562 ;
      RECT 8.498 9.968 8.566 10.012 ;
      RECT 8.282 0.068 8.35 0.112 ;
      RECT 8.282 0.518 8.35 0.562 ;
      RECT 8.282 1.328 8.35 1.372 ;
      RECT 8.282 1.778 8.35 1.822 ;
      RECT 8.282 1.958 8.35 2.002 ;
      RECT 8.282 2.408 8.35 2.452 ;
      RECT 8.282 2.588 8.35 2.632 ;
      RECT 8.282 3.038 8.35 3.082 ;
      RECT 8.282 3.218 8.35 3.262 ;
      RECT 8.282 3.668 8.35 3.712 ;
      RECT 8.282 3.848 8.35 3.892 ;
      RECT 8.282 4.298 8.35 4.342 ;
      RECT 8.282 4.478 8.35 4.522 ;
      RECT 8.282 4.928 8.35 4.972 ;
      RECT 8.282 5.108 8.35 5.152 ;
      RECT 8.282 5.558 8.35 5.602 ;
      RECT 8.282 5.738 8.35 5.782 ;
      RECT 8.282 6.188 8.35 6.232 ;
      RECT 8.282 6.368 8.35 6.412 ;
      RECT 8.282 6.818 8.35 6.862 ;
      RECT 8.282 6.998 8.35 7.042 ;
      RECT 8.282 7.448 8.35 7.492 ;
      RECT 8.282 7.628 8.35 7.672 ;
      RECT 8.282 8.078 8.35 8.122 ;
      RECT 8.282 8.258 8.35 8.302 ;
      RECT 8.282 8.708 8.35 8.752 ;
      RECT 8.282 9.518 8.35 9.562 ;
      RECT 8.282 9.968 8.35 10.012 ;
      RECT 8.066 0.068 8.134 0.112 ;
      RECT 8.066 0.518 8.134 0.562 ;
      RECT 8.066 1.958 8.134 2.002 ;
      RECT 8.066 2.408 8.134 2.452 ;
      RECT 8.066 2.588 8.134 2.632 ;
      RECT 8.066 3.038 8.134 3.082 ;
      RECT 8.066 3.218 8.134 3.262 ;
      RECT 8.066 3.668 8.134 3.712 ;
      RECT 8.066 3.848 8.134 3.892 ;
      RECT 8.066 4.298 8.134 4.342 ;
      RECT 8.066 4.478 8.134 4.522 ;
      RECT 8.066 4.928 8.134 4.972 ;
      RECT 8.066 5.108 8.134 5.152 ;
      RECT 8.066 5.558 8.134 5.602 ;
      RECT 8.066 5.738 8.134 5.782 ;
      RECT 8.066 6.188 8.134 6.232 ;
      RECT 8.066 6.368 8.134 6.412 ;
      RECT 8.066 6.818 8.134 6.862 ;
      RECT 8.066 6.998 8.134 7.042 ;
      RECT 8.066 7.448 8.134 7.492 ;
      RECT 8.066 7.628 8.134 7.672 ;
      RECT 8.066 8.078 8.134 8.122 ;
      RECT 8.066 9.518 8.134 9.562 ;
      RECT 8.066 9.968 8.134 10.012 ;
      RECT 7.85 0.068 7.918 0.112 ;
      RECT 7.85 0.518 7.918 0.562 ;
      RECT 7.85 1.958 7.918 2.002 ;
      RECT 7.85 2.408 7.918 2.452 ;
      RECT 7.85 2.588 7.918 2.632 ;
      RECT 7.85 3.038 7.918 3.082 ;
      RECT 7.85 3.218 7.918 3.262 ;
      RECT 7.85 3.668 7.918 3.712 ;
      RECT 7.85 3.848 7.918 3.892 ;
      RECT 7.85 4.298 7.918 4.342 ;
      RECT 7.85 4.478 7.918 4.522 ;
      RECT 7.85 4.928 7.918 4.972 ;
      RECT 7.85 5.108 7.918 5.152 ;
      RECT 7.85 5.558 7.918 5.602 ;
      RECT 7.85 5.738 7.918 5.782 ;
      RECT 7.85 6.188 7.918 6.232 ;
      RECT 7.85 6.368 7.918 6.412 ;
      RECT 7.85 6.818 7.918 6.862 ;
      RECT 7.85 6.998 7.918 7.042 ;
      RECT 7.85 7.448 7.918 7.492 ;
      RECT 7.85 7.628 7.918 7.672 ;
      RECT 7.85 8.078 7.918 8.122 ;
      RECT 7.85 9.518 7.918 9.562 ;
      RECT 7.85 9.968 7.918 10.012 ;
      RECT 7.634 0.068 7.702 0.112 ;
      RECT 7.634 0.518 7.702 0.562 ;
      RECT 7.634 2.588 7.702 2.632 ;
      RECT 7.634 3.038 7.702 3.082 ;
      RECT 7.634 3.218 7.702 3.262 ;
      RECT 7.634 3.668 7.702 3.712 ;
      RECT 7.634 3.848 7.702 3.892 ;
      RECT 7.634 4.298 7.702 4.342 ;
      RECT 7.634 4.478 7.702 4.522 ;
      RECT 7.634 4.928 7.702 4.972 ;
      RECT 7.634 5.108 7.702 5.152 ;
      RECT 7.634 5.558 7.702 5.602 ;
      RECT 7.634 5.738 7.702 5.782 ;
      RECT 7.634 6.188 7.702 6.232 ;
      RECT 7.634 6.368 7.702 6.412 ;
      RECT 7.634 6.818 7.702 6.862 ;
      RECT 7.634 6.998 7.702 7.042 ;
      RECT 7.634 7.448 7.702 7.492 ;
      RECT 7.634 9.518 7.702 9.562 ;
      RECT 7.634 9.968 7.702 10.012 ;
      RECT 7.418 0.068 7.486 0.112 ;
      RECT 7.418 0.518 7.486 0.562 ;
      RECT 7.418 2.588 7.486 2.632 ;
      RECT 7.418 3.038 7.486 3.082 ;
      RECT 7.418 3.218 7.486 3.262 ;
      RECT 7.418 3.668 7.486 3.712 ;
      RECT 7.418 3.848 7.486 3.892 ;
      RECT 7.418 4.298 7.486 4.342 ;
      RECT 7.418 4.478 7.486 4.522 ;
      RECT 7.418 4.928 7.486 4.972 ;
      RECT 7.418 5.108 7.486 5.152 ;
      RECT 7.418 5.558 7.486 5.602 ;
      RECT 7.418 5.738 7.486 5.782 ;
      RECT 7.418 6.188 7.486 6.232 ;
      RECT 7.418 6.368 7.486 6.412 ;
      RECT 7.418 6.818 7.486 6.862 ;
      RECT 7.418 6.998 7.486 7.042 ;
      RECT 7.418 7.448 7.486 7.492 ;
      RECT 7.418 9.518 7.486 9.562 ;
      RECT 7.418 9.968 7.486 10.012 ;
      RECT 7.202 0.068 7.27 0.112 ;
      RECT 7.202 0.518 7.27 0.562 ;
      RECT 7.202 0.698 7.27 0.742 ;
      RECT 7.202 1.148 7.27 1.192 ;
      RECT 7.202 3.218 7.27 3.262 ;
      RECT 7.202 3.668 7.27 3.712 ;
      RECT 7.202 3.848 7.27 3.892 ;
      RECT 7.202 4.298 7.27 4.342 ;
      RECT 7.202 4.478 7.27 4.522 ;
      RECT 7.202 4.928 7.27 4.972 ;
      RECT 7.202 5.108 7.27 5.152 ;
      RECT 7.202 5.558 7.27 5.602 ;
      RECT 7.202 5.738 7.27 5.782 ;
      RECT 7.202 6.188 7.27 6.232 ;
      RECT 7.202 6.368 7.27 6.412 ;
      RECT 7.202 6.818 7.27 6.862 ;
      RECT 7.202 8.888 7.27 8.932 ;
      RECT 7.202 9.338 7.27 9.382 ;
      RECT 7.202 9.518 7.27 9.562 ;
      RECT 7.202 9.968 7.27 10.012 ;
      RECT 6.986 0.068 7.054 0.112 ;
      RECT 6.986 0.518 7.054 0.562 ;
      RECT 6.986 0.698 7.054 0.742 ;
      RECT 6.986 1.148 7.054 1.192 ;
      RECT 6.986 3.218 7.054 3.262 ;
      RECT 6.986 3.668 7.054 3.712 ;
      RECT 6.986 3.848 7.054 3.892 ;
      RECT 6.986 4.298 7.054 4.342 ;
      RECT 6.986 4.478 7.054 4.522 ;
      RECT 6.986 4.928 7.054 4.972 ;
      RECT 6.986 5.108 7.054 5.152 ;
      RECT 6.986 5.558 7.054 5.602 ;
      RECT 6.986 5.738 7.054 5.782 ;
      RECT 6.986 6.188 7.054 6.232 ;
      RECT 6.986 6.368 7.054 6.412 ;
      RECT 6.986 6.818 7.054 6.862 ;
      RECT 6.986 8.888 7.054 8.932 ;
      RECT 6.986 9.338 7.054 9.382 ;
      RECT 6.986 9.518 7.054 9.562 ;
      RECT 6.986 9.968 7.054 10.012 ;
      RECT 6.77 0.068 6.838 0.112 ;
      RECT 6.77 0.518 6.838 0.562 ;
      RECT 6.77 0.698 6.838 0.742 ;
      RECT 6.77 1.148 6.838 1.192 ;
      RECT 6.77 1.328 6.838 1.372 ;
      RECT 6.77 1.778 6.838 1.822 ;
      RECT 6.77 3.848 6.838 3.892 ;
      RECT 6.77 4.298 6.838 4.342 ;
      RECT 6.77 4.478 6.838 4.522 ;
      RECT 6.77 4.928 6.838 4.972 ;
      RECT 6.77 5.108 6.838 5.152 ;
      RECT 6.77 5.558 6.838 5.602 ;
      RECT 6.77 5.738 6.838 5.782 ;
      RECT 6.77 6.188 6.838 6.232 ;
      RECT 6.77 8.258 6.838 8.302 ;
      RECT 6.77 8.708 6.838 8.752 ;
      RECT 6.77 8.888 6.838 8.932 ;
      RECT 6.77 9.338 6.838 9.382 ;
      RECT 6.77 9.518 6.838 9.562 ;
      RECT 6.77 9.968 6.838 10.012 ;
      RECT 6.554 0.068 6.622 0.112 ;
      RECT 6.554 0.518 6.622 0.562 ;
      RECT 6.554 0.698 6.622 0.742 ;
      RECT 6.554 1.148 6.622 1.192 ;
      RECT 6.554 1.328 6.622 1.372 ;
      RECT 6.554 1.778 6.622 1.822 ;
      RECT 6.554 3.848 6.622 3.892 ;
      RECT 6.554 4.298 6.622 4.342 ;
      RECT 6.554 4.478 6.622 4.522 ;
      RECT 6.554 4.928 6.622 4.972 ;
      RECT 6.554 5.108 6.622 5.152 ;
      RECT 6.554 5.558 6.622 5.602 ;
      RECT 6.554 5.738 6.622 5.782 ;
      RECT 6.554 6.188 6.622 6.232 ;
      RECT 6.554 8.258 6.622 8.302 ;
      RECT 6.554 8.708 6.622 8.752 ;
      RECT 6.554 8.888 6.622 8.932 ;
      RECT 6.554 9.338 6.622 9.382 ;
      RECT 6.554 9.518 6.622 9.562 ;
      RECT 6.554 9.968 6.622 10.012 ;
      RECT 6.338 0.068 6.406 0.112 ;
      RECT 6.338 0.518 6.406 0.562 ;
      RECT 6.338 0.698 6.406 0.742 ;
      RECT 6.338 1.148 6.406 1.192 ;
      RECT 6.338 1.328 6.406 1.372 ;
      RECT 6.338 1.778 6.406 1.822 ;
      RECT 6.338 1.958 6.406 2.002 ;
      RECT 6.338 2.408 6.406 2.452 ;
      RECT 6.338 4.478 6.406 4.522 ;
      RECT 6.338 4.928 6.406 4.972 ;
      RECT 6.338 5.108 6.406 5.152 ;
      RECT 6.338 5.558 6.406 5.602 ;
      RECT 6.338 7.628 6.406 7.672 ;
      RECT 6.338 8.078 6.406 8.122 ;
      RECT 6.338 8.258 6.406 8.302 ;
      RECT 6.338 8.708 6.406 8.752 ;
      RECT 6.338 8.888 6.406 8.932 ;
      RECT 6.338 9.338 6.406 9.382 ;
      RECT 6.338 9.518 6.406 9.562 ;
      RECT 6.338 9.968 6.406 10.012 ;
      RECT 6.122 0.068 6.19 0.112 ;
      RECT 6.122 0.518 6.19 0.562 ;
      RECT 6.122 0.698 6.19 0.742 ;
      RECT 6.122 1.148 6.19 1.192 ;
      RECT 6.122 1.328 6.19 1.372 ;
      RECT 6.122 1.778 6.19 1.822 ;
      RECT 6.122 1.958 6.19 2.002 ;
      RECT 6.122 2.408 6.19 2.452 ;
      RECT 6.122 4.478 6.19 4.522 ;
      RECT 6.122 4.928 6.19 4.972 ;
      RECT 6.122 5.108 6.19 5.152 ;
      RECT 6.122 5.558 6.19 5.602 ;
      RECT 6.122 7.628 6.19 7.672 ;
      RECT 6.122 8.078 6.19 8.122 ;
      RECT 6.122 8.258 6.19 8.302 ;
      RECT 6.122 8.708 6.19 8.752 ;
      RECT 6.122 8.888 6.19 8.932 ;
      RECT 6.122 9.338 6.19 9.382 ;
      RECT 6.122 9.518 6.19 9.562 ;
      RECT 6.122 9.968 6.19 10.012 ;
      RECT 5.906 0.068 5.974 0.112 ;
      RECT 5.906 0.518 5.974 0.562 ;
      RECT 5.906 0.698 5.974 0.742 ;
      RECT 5.906 1.148 5.974 1.192 ;
      RECT 5.906 1.328 5.974 1.372 ;
      RECT 5.906 1.778 5.974 1.822 ;
      RECT 5.906 1.958 5.974 2.002 ;
      RECT 5.906 2.408 5.974 2.452 ;
      RECT 5.906 2.588 5.974 2.632 ;
      RECT 5.906 3.038 5.974 3.082 ;
      RECT 5.906 4.478 5.974 4.522 ;
      RECT 5.906 4.928 5.974 4.972 ;
      RECT 5.906 5.108 5.974 5.152 ;
      RECT 5.906 5.558 5.974 5.602 ;
      RECT 5.906 6.998 5.974 7.042 ;
      RECT 5.906 7.448 5.974 7.492 ;
      RECT 5.906 7.628 5.974 7.672 ;
      RECT 5.906 8.078 5.974 8.122 ;
      RECT 5.906 8.258 5.974 8.302 ;
      RECT 5.906 8.708 5.974 8.752 ;
      RECT 5.906 8.888 5.974 8.932 ;
      RECT 5.906 9.338 5.974 9.382 ;
      RECT 5.906 9.518 5.974 9.562 ;
      RECT 5.906 9.968 5.974 10.012 ;
      RECT 5.69 0.068 5.758 0.112 ;
      RECT 5.69 0.518 5.758 0.562 ;
      RECT 5.69 0.698 5.758 0.742 ;
      RECT 5.69 1.148 5.758 1.192 ;
      RECT 5.69 1.328 5.758 1.372 ;
      RECT 5.69 1.778 5.758 1.822 ;
      RECT 5.69 1.958 5.758 2.002 ;
      RECT 5.69 2.408 5.758 2.452 ;
      RECT 5.69 2.588 5.758 2.632 ;
      RECT 5.69 3.038 5.758 3.082 ;
      RECT 5.69 4.478 5.758 4.522 ;
      RECT 5.69 4.928 5.758 4.972 ;
      RECT 5.69 5.108 5.758 5.152 ;
      RECT 5.69 5.558 5.758 5.602 ;
      RECT 5.69 6.998 5.758 7.042 ;
      RECT 5.69 7.448 5.758 7.492 ;
      RECT 5.69 7.628 5.758 7.672 ;
      RECT 5.69 8.078 5.758 8.122 ;
      RECT 5.69 8.258 5.758 8.302 ;
      RECT 5.69 8.708 5.758 8.752 ;
      RECT 5.69 8.888 5.758 8.932 ;
      RECT 5.69 9.338 5.758 9.382 ;
      RECT 5.69 9.518 5.758 9.562 ;
      RECT 5.69 9.968 5.758 10.012 ;
      RECT 5.474 0.068 5.542 0.112 ;
      RECT 5.474 0.518 5.542 0.562 ;
      RECT 5.474 0.698 5.542 0.742 ;
      RECT 5.474 1.148 5.542 1.192 ;
      RECT 5.474 1.328 5.542 1.372 ;
      RECT 5.474 1.778 5.542 1.822 ;
      RECT 5.474 1.958 5.542 2.002 ;
      RECT 5.474 2.408 5.542 2.452 ;
      RECT 5.474 2.588 5.542 2.632 ;
      RECT 5.474 3.038 5.542 3.082 ;
      RECT 5.474 3.218 5.542 3.262 ;
      RECT 5.474 3.668 5.542 3.712 ;
      RECT 5.474 6.368 5.542 6.412 ;
      RECT 5.474 6.818 5.542 6.862 ;
      RECT 5.474 6.998 5.542 7.042 ;
      RECT 5.474 7.448 5.542 7.492 ;
      RECT 5.474 7.628 5.542 7.672 ;
      RECT 5.474 8.078 5.542 8.122 ;
      RECT 5.474 8.258 5.542 8.302 ;
      RECT 5.474 8.708 5.542 8.752 ;
      RECT 5.474 8.888 5.542 8.932 ;
      RECT 5.474 9.338 5.542 9.382 ;
      RECT 5.474 9.518 5.542 9.562 ;
      RECT 5.474 9.968 5.542 10.012 ;
      RECT 5.258 0.068 5.326 0.112 ;
      RECT 5.258 0.518 5.326 0.562 ;
      RECT 5.258 0.698 5.326 0.742 ;
      RECT 5.258 1.148 5.326 1.192 ;
      RECT 5.258 1.328 5.326 1.372 ;
      RECT 5.258 1.778 5.326 1.822 ;
      RECT 5.258 1.958 5.326 2.002 ;
      RECT 5.258 2.408 5.326 2.452 ;
      RECT 5.258 2.588 5.326 2.632 ;
      RECT 5.258 3.038 5.326 3.082 ;
      RECT 5.258 3.218 5.326 3.262 ;
      RECT 5.258 3.668 5.326 3.712 ;
      RECT 5.258 6.368 5.326 6.412 ;
      RECT 5.258 6.818 5.326 6.862 ;
      RECT 5.258 6.998 5.326 7.042 ;
      RECT 5.258 7.448 5.326 7.492 ;
      RECT 5.258 7.628 5.326 7.672 ;
      RECT 5.258 8.078 5.326 8.122 ;
      RECT 5.258 8.258 5.326 8.302 ;
      RECT 5.258 8.708 5.326 8.752 ;
      RECT 5.258 8.888 5.326 8.932 ;
      RECT 5.258 9.338 5.326 9.382 ;
      RECT 5.258 9.518 5.326 9.562 ;
      RECT 5.258 9.968 5.326 10.012 ;
      RECT 5.042 0.068 5.11 0.112 ;
      RECT 5.042 0.518 5.11 0.562 ;
      RECT 5.042 0.698 5.11 0.742 ;
      RECT 5.042 1.148 5.11 1.192 ;
      RECT 5.042 1.328 5.11 1.372 ;
      RECT 5.042 1.778 5.11 1.822 ;
      RECT 5.042 1.958 5.11 2.002 ;
      RECT 5.042 2.408 5.11 2.452 ;
      RECT 5.042 2.588 5.11 2.632 ;
      RECT 5.042 3.038 5.11 3.082 ;
      RECT 5.042 3.218 5.11 3.262 ;
      RECT 5.042 3.668 5.11 3.712 ;
      RECT 5.042 3.848 5.11 3.892 ;
      RECT 5.042 4.298 5.11 4.342 ;
      RECT 5.042 5.738 5.11 5.782 ;
      RECT 5.042 6.188 5.11 6.232 ;
      RECT 5.042 6.368 5.11 6.412 ;
      RECT 5.042 6.818 5.11 6.862 ;
      RECT 5.042 6.998 5.11 7.042 ;
      RECT 5.042 7.448 5.11 7.492 ;
      RECT 5.042 7.628 5.11 7.672 ;
      RECT 5.042 8.078 5.11 8.122 ;
      RECT 5.042 8.258 5.11 8.302 ;
      RECT 5.042 8.708 5.11 8.752 ;
      RECT 5.042 8.888 5.11 8.932 ;
      RECT 5.042 9.338 5.11 9.382 ;
      RECT 5.042 9.518 5.11 9.562 ;
      RECT 5.042 9.968 5.11 10.012 ;
      RECT 4.826 0.068 4.894 0.112 ;
      RECT 4.826 0.518 4.894 0.562 ;
      RECT 4.826 0.698 4.894 0.742 ;
      RECT 4.826 1.148 4.894 1.192 ;
      RECT 4.826 1.328 4.894 1.372 ;
      RECT 4.826 1.778 4.894 1.822 ;
      RECT 4.826 1.958 4.894 2.002 ;
      RECT 4.826 2.408 4.894 2.452 ;
      RECT 4.826 2.588 4.894 2.632 ;
      RECT 4.826 3.038 4.894 3.082 ;
      RECT 4.826 3.218 4.894 3.262 ;
      RECT 4.826 3.668 4.894 3.712 ;
      RECT 4.826 3.848 4.894 3.892 ;
      RECT 4.826 4.298 4.894 4.342 ;
      RECT 4.826 5.738 4.894 5.782 ;
      RECT 4.826 6.188 4.894 6.232 ;
      RECT 4.826 6.368 4.894 6.412 ;
      RECT 4.826 6.818 4.894 6.862 ;
      RECT 4.826 6.998 4.894 7.042 ;
      RECT 4.826 7.448 4.894 7.492 ;
      RECT 4.826 7.628 4.894 7.672 ;
      RECT 4.826 8.078 4.894 8.122 ;
      RECT 4.826 8.258 4.894 8.302 ;
      RECT 4.826 8.708 4.894 8.752 ;
      RECT 4.826 8.888 4.894 8.932 ;
      RECT 4.826 9.338 4.894 9.382 ;
      RECT 4.826 9.518 4.894 9.562 ;
      RECT 4.826 9.968 4.894 10.012 ;
      RECT 4.61 0.068 4.678 0.112 ;
      RECT 4.61 0.518 4.678 0.562 ;
      RECT 4.61 0.698 4.678 0.742 ;
      RECT 4.61 1.148 4.678 1.192 ;
      RECT 4.61 1.328 4.678 1.372 ;
      RECT 4.61 1.778 4.678 1.822 ;
      RECT 4.61 1.958 4.678 2.002 ;
      RECT 4.61 2.408 4.678 2.452 ;
      RECT 4.61 2.588 4.678 2.632 ;
      RECT 4.61 3.038 4.678 3.082 ;
      RECT 4.61 3.218 4.678 3.262 ;
      RECT 4.61 3.668 4.678 3.712 ;
      RECT 4.61 3.848 4.678 3.892 ;
      RECT 4.61 4.298 4.678 4.342 ;
      RECT 4.61 5.738 4.678 5.782 ;
      RECT 4.61 6.188 4.678 6.232 ;
      RECT 4.61 6.368 4.678 6.412 ;
      RECT 4.61 6.818 4.678 6.862 ;
      RECT 4.61 6.998 4.678 7.042 ;
      RECT 4.61 7.448 4.678 7.492 ;
      RECT 4.61 7.628 4.678 7.672 ;
      RECT 4.61 8.078 4.678 8.122 ;
      RECT 4.61 8.258 4.678 8.302 ;
      RECT 4.61 8.708 4.678 8.752 ;
      RECT 4.61 8.888 4.678 8.932 ;
      RECT 4.61 9.338 4.678 9.382 ;
      RECT 4.61 9.518 4.678 9.562 ;
      RECT 4.61 9.968 4.678 10.012 ;
      RECT 4.394 0.068 4.462 0.112 ;
      RECT 4.394 0.518 4.462 0.562 ;
      RECT 4.394 0.698 4.462 0.742 ;
      RECT 4.394 1.148 4.462 1.192 ;
      RECT 4.394 1.328 4.462 1.372 ;
      RECT 4.394 1.778 4.462 1.822 ;
      RECT 4.394 1.958 4.462 2.002 ;
      RECT 4.394 2.408 4.462 2.452 ;
      RECT 4.394 2.588 4.462 2.632 ;
      RECT 4.394 3.038 4.462 3.082 ;
      RECT 4.394 3.218 4.462 3.262 ;
      RECT 4.394 3.668 4.462 3.712 ;
      RECT 4.394 3.848 4.462 3.892 ;
      RECT 4.394 4.298 4.462 4.342 ;
      RECT 4.394 5.738 4.462 5.782 ;
      RECT 4.394 6.188 4.462 6.232 ;
      RECT 4.394 6.368 4.462 6.412 ;
      RECT 4.394 6.818 4.462 6.862 ;
      RECT 4.394 6.998 4.462 7.042 ;
      RECT 4.394 7.448 4.462 7.492 ;
      RECT 4.394 7.628 4.462 7.672 ;
      RECT 4.394 8.078 4.462 8.122 ;
      RECT 4.394 8.258 4.462 8.302 ;
      RECT 4.394 8.708 4.462 8.752 ;
      RECT 4.394 8.888 4.462 8.932 ;
      RECT 4.394 9.338 4.462 9.382 ;
      RECT 4.394 9.518 4.462 9.562 ;
      RECT 4.394 9.968 4.462 10.012 ;
      RECT 4.178 0.068 4.246 0.112 ;
      RECT 4.178 0.518 4.246 0.562 ;
      RECT 4.178 0.698 4.246 0.742 ;
      RECT 4.178 1.148 4.246 1.192 ;
      RECT 4.178 1.328 4.246 1.372 ;
      RECT 4.178 1.778 4.246 1.822 ;
      RECT 4.178 1.958 4.246 2.002 ;
      RECT 4.178 2.408 4.246 2.452 ;
      RECT 4.178 2.588 4.246 2.632 ;
      RECT 4.178 3.038 4.246 3.082 ;
      RECT 4.178 3.218 4.246 3.262 ;
      RECT 4.178 3.668 4.246 3.712 ;
      RECT 4.178 6.368 4.246 6.412 ;
      RECT 4.178 6.818 4.246 6.862 ;
      RECT 4.178 6.998 4.246 7.042 ;
      RECT 4.178 7.448 4.246 7.492 ;
      RECT 4.178 7.628 4.246 7.672 ;
      RECT 4.178 8.078 4.246 8.122 ;
      RECT 4.178 8.258 4.246 8.302 ;
      RECT 4.178 8.708 4.246 8.752 ;
      RECT 4.178 8.888 4.246 8.932 ;
      RECT 4.178 9.338 4.246 9.382 ;
      RECT 4.178 9.518 4.246 9.562 ;
      RECT 4.178 9.968 4.246 10.012 ;
      RECT 3.962 0.068 4.03 0.112 ;
      RECT 3.962 0.518 4.03 0.562 ;
      RECT 3.962 0.698 4.03 0.742 ;
      RECT 3.962 1.148 4.03 1.192 ;
      RECT 3.962 1.328 4.03 1.372 ;
      RECT 3.962 1.778 4.03 1.822 ;
      RECT 3.962 1.958 4.03 2.002 ;
      RECT 3.962 2.408 4.03 2.452 ;
      RECT 3.962 2.588 4.03 2.632 ;
      RECT 3.962 3.038 4.03 3.082 ;
      RECT 3.962 3.218 4.03 3.262 ;
      RECT 3.962 3.668 4.03 3.712 ;
      RECT 3.962 6.368 4.03 6.412 ;
      RECT 3.962 6.818 4.03 6.862 ;
      RECT 3.962 6.998 4.03 7.042 ;
      RECT 3.962 7.448 4.03 7.492 ;
      RECT 3.962 7.628 4.03 7.672 ;
      RECT 3.962 8.078 4.03 8.122 ;
      RECT 3.962 8.258 4.03 8.302 ;
      RECT 3.962 8.708 4.03 8.752 ;
      RECT 3.962 8.888 4.03 8.932 ;
      RECT 3.962 9.338 4.03 9.382 ;
      RECT 3.962 9.518 4.03 9.562 ;
      RECT 3.962 9.968 4.03 10.012 ;
      RECT 3.746 0.068 3.814 0.112 ;
      RECT 3.746 0.518 3.814 0.562 ;
      RECT 3.746 0.698 3.814 0.742 ;
      RECT 3.746 1.148 3.814 1.192 ;
      RECT 3.746 1.328 3.814 1.372 ;
      RECT 3.746 1.778 3.814 1.822 ;
      RECT 3.746 1.958 3.814 2.002 ;
      RECT 3.746 2.408 3.814 2.452 ;
      RECT 3.746 2.588 3.814 2.632 ;
      RECT 3.746 3.038 3.814 3.082 ;
      RECT 3.746 4.478 3.814 4.522 ;
      RECT 3.746 4.928 3.814 4.972 ;
      RECT 3.746 5.108 3.814 5.152 ;
      RECT 3.746 5.558 3.814 5.602 ;
      RECT 3.746 6.998 3.814 7.042 ;
      RECT 3.746 7.448 3.814 7.492 ;
      RECT 3.746 7.628 3.814 7.672 ;
      RECT 3.746 8.078 3.814 8.122 ;
      RECT 3.746 8.258 3.814 8.302 ;
      RECT 3.746 8.708 3.814 8.752 ;
      RECT 3.746 8.888 3.814 8.932 ;
      RECT 3.746 9.338 3.814 9.382 ;
      RECT 3.746 9.518 3.814 9.562 ;
      RECT 3.746 9.968 3.814 10.012 ;
      RECT 3.53 0.068 3.598 0.112 ;
      RECT 3.53 0.518 3.598 0.562 ;
      RECT 3.53 0.698 3.598 0.742 ;
      RECT 3.53 1.148 3.598 1.192 ;
      RECT 3.53 1.328 3.598 1.372 ;
      RECT 3.53 1.778 3.598 1.822 ;
      RECT 3.53 1.958 3.598 2.002 ;
      RECT 3.53 2.408 3.598 2.452 ;
      RECT 3.53 2.588 3.598 2.632 ;
      RECT 3.53 3.038 3.598 3.082 ;
      RECT 3.53 4.478 3.598 4.522 ;
      RECT 3.53 4.928 3.598 4.972 ;
      RECT 3.53 5.108 3.598 5.152 ;
      RECT 3.53 5.558 3.598 5.602 ;
      RECT 3.53 6.998 3.598 7.042 ;
      RECT 3.53 7.448 3.598 7.492 ;
      RECT 3.53 7.628 3.598 7.672 ;
      RECT 3.53 8.078 3.598 8.122 ;
      RECT 3.53 8.258 3.598 8.302 ;
      RECT 3.53 8.708 3.598 8.752 ;
      RECT 3.53 8.888 3.598 8.932 ;
      RECT 3.53 9.338 3.598 9.382 ;
      RECT 3.53 9.518 3.598 9.562 ;
      RECT 3.53 9.968 3.598 10.012 ;
      RECT 3.314 0.068 3.382 0.112 ;
      RECT 3.314 0.518 3.382 0.562 ;
      RECT 3.314 0.698 3.382 0.742 ;
      RECT 3.314 1.148 3.382 1.192 ;
      RECT 3.314 1.328 3.382 1.372 ;
      RECT 3.314 1.778 3.382 1.822 ;
      RECT 3.314 1.958 3.382 2.002 ;
      RECT 3.314 2.408 3.382 2.452 ;
      RECT 3.314 4.478 3.382 4.522 ;
      RECT 3.314 4.928 3.382 4.972 ;
      RECT 3.314 5.108 3.382 5.152 ;
      RECT 3.314 5.558 3.382 5.602 ;
      RECT 3.314 7.628 3.382 7.672 ;
      RECT 3.314 8.078 3.382 8.122 ;
      RECT 3.314 8.258 3.382 8.302 ;
      RECT 3.314 8.708 3.382 8.752 ;
      RECT 3.314 8.888 3.382 8.932 ;
      RECT 3.314 9.338 3.382 9.382 ;
      RECT 3.314 9.518 3.382 9.562 ;
      RECT 3.314 9.968 3.382 10.012 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 3.098 0.518 3.166 0.562 ;
      RECT 3.098 0.698 3.166 0.742 ;
      RECT 3.098 1.148 3.166 1.192 ;
      RECT 3.098 1.328 3.166 1.372 ;
      RECT 3.098 1.778 3.166 1.822 ;
      RECT 3.098 1.958 3.166 2.002 ;
      RECT 3.098 2.408 3.166 2.452 ;
      RECT 3.098 4.478 3.166 4.522 ;
      RECT 3.098 4.928 3.166 4.972 ;
      RECT 3.098 5.108 3.166 5.152 ;
      RECT 3.098 5.558 3.166 5.602 ;
      RECT 3.098 7.628 3.166 7.672 ;
      RECT 3.098 8.078 3.166 8.122 ;
      RECT 3.098 8.258 3.166 8.302 ;
      RECT 3.098 8.708 3.166 8.752 ;
      RECT 3.098 8.888 3.166 8.932 ;
      RECT 3.098 9.338 3.166 9.382 ;
      RECT 3.098 9.518 3.166 9.562 ;
      RECT 3.098 9.968 3.166 10.012 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.882 0.518 2.95 0.562 ;
      RECT 2.882 0.698 2.95 0.742 ;
      RECT 2.882 1.148 2.95 1.192 ;
      RECT 2.882 1.328 2.95 1.372 ;
      RECT 2.882 1.778 2.95 1.822 ;
      RECT 2.882 3.848 2.95 3.892 ;
      RECT 2.882 4.298 2.95 4.342 ;
      RECT 2.882 4.478 2.95 4.522 ;
      RECT 2.882 4.928 2.95 4.972 ;
      RECT 2.882 5.108 2.95 5.152 ;
      RECT 2.882 5.558 2.95 5.602 ;
      RECT 2.882 5.738 2.95 5.782 ;
      RECT 2.882 6.188 2.95 6.232 ;
      RECT 2.882 8.258 2.95 8.302 ;
      RECT 2.882 8.708 2.95 8.752 ;
      RECT 2.882 8.888 2.95 8.932 ;
      RECT 2.882 9.338 2.95 9.382 ;
      RECT 2.882 9.518 2.95 9.562 ;
      RECT 2.882 9.968 2.95 10.012 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.666 0.698 2.734 0.742 ;
      RECT 2.666 1.148 2.734 1.192 ;
      RECT 2.666 1.328 2.734 1.372 ;
      RECT 2.666 1.778 2.734 1.822 ;
      RECT 2.666 3.848 2.734 3.892 ;
      RECT 2.666 4.298 2.734 4.342 ;
      RECT 2.666 4.478 2.734 4.522 ;
      RECT 2.666 4.928 2.734 4.972 ;
      RECT 2.666 5.108 2.734 5.152 ;
      RECT 2.666 5.558 2.734 5.602 ;
      RECT 2.666 5.738 2.734 5.782 ;
      RECT 2.666 6.188 2.734 6.232 ;
      RECT 2.666 8.258 2.734 8.302 ;
      RECT 2.666 8.708 2.734 8.752 ;
      RECT 2.666 8.888 2.734 8.932 ;
      RECT 2.666 9.338 2.734 9.382 ;
      RECT 2.666 9.518 2.734 9.562 ;
      RECT 2.666 9.968 2.734 10.012 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.45 0.518 2.518 0.562 ;
      RECT 2.45 0.698 2.518 0.742 ;
      RECT 2.45 1.148 2.518 1.192 ;
      RECT 2.45 3.218 2.518 3.262 ;
      RECT 2.45 3.668 2.518 3.712 ;
      RECT 2.45 3.848 2.518 3.892 ;
      RECT 2.45 4.298 2.518 4.342 ;
      RECT 2.45 4.478 2.518 4.522 ;
      RECT 2.45 4.928 2.518 4.972 ;
      RECT 2.45 5.108 2.518 5.152 ;
      RECT 2.45 5.558 2.518 5.602 ;
      RECT 2.45 5.738 2.518 5.782 ;
      RECT 2.45 6.188 2.518 6.232 ;
      RECT 2.45 6.368 2.518 6.412 ;
      RECT 2.45 6.818 2.518 6.862 ;
      RECT 2.45 8.888 2.518 8.932 ;
      RECT 2.45 9.338 2.518 9.382 ;
      RECT 2.45 9.518 2.518 9.562 ;
      RECT 2.45 9.968 2.518 10.012 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.234 0.698 2.302 0.742 ;
      RECT 2.234 1.148 2.302 1.192 ;
      RECT 2.234 3.218 2.302 3.262 ;
      RECT 2.234 3.668 2.302 3.712 ;
      RECT 2.234 3.848 2.302 3.892 ;
      RECT 2.234 4.298 2.302 4.342 ;
      RECT 2.234 4.478 2.302 4.522 ;
      RECT 2.234 4.928 2.302 4.972 ;
      RECT 2.234 5.108 2.302 5.152 ;
      RECT 2.234 5.558 2.302 5.602 ;
      RECT 2.234 5.738 2.302 5.782 ;
      RECT 2.234 6.188 2.302 6.232 ;
      RECT 2.234 6.368 2.302 6.412 ;
      RECT 2.234 6.818 2.302 6.862 ;
      RECT 2.234 8.888 2.302 8.932 ;
      RECT 2.234 9.338 2.302 9.382 ;
      RECT 2.234 9.518 2.302 9.562 ;
      RECT 2.234 9.968 2.302 10.012 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 2.018 2.588 2.086 2.632 ;
      RECT 2.018 3.038 2.086 3.082 ;
      RECT 2.018 3.218 2.086 3.262 ;
      RECT 2.018 3.668 2.086 3.712 ;
      RECT 2.018 3.848 2.086 3.892 ;
      RECT 2.018 4.298 2.086 4.342 ;
      RECT 2.018 4.478 2.086 4.522 ;
      RECT 2.018 4.928 2.086 4.972 ;
      RECT 2.018 5.108 2.086 5.152 ;
      RECT 2.018 5.558 2.086 5.602 ;
      RECT 2.018 5.738 2.086 5.782 ;
      RECT 2.018 6.188 2.086 6.232 ;
      RECT 2.018 6.368 2.086 6.412 ;
      RECT 2.018 6.818 2.086 6.862 ;
      RECT 2.018 6.998 2.086 7.042 ;
      RECT 2.018 7.448 2.086 7.492 ;
      RECT 2.018 9.518 2.086 9.562 ;
      RECT 2.018 9.968 2.086 10.012 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.802 2.588 1.87 2.632 ;
      RECT 1.802 3.038 1.87 3.082 ;
      RECT 1.802 3.218 1.87 3.262 ;
      RECT 1.802 3.668 1.87 3.712 ;
      RECT 1.802 3.848 1.87 3.892 ;
      RECT 1.802 4.298 1.87 4.342 ;
      RECT 1.802 4.478 1.87 4.522 ;
      RECT 1.802 4.928 1.87 4.972 ;
      RECT 1.802 5.108 1.87 5.152 ;
      RECT 1.802 5.558 1.87 5.602 ;
      RECT 1.802 5.738 1.87 5.782 ;
      RECT 1.802 6.188 1.87 6.232 ;
      RECT 1.802 6.368 1.87 6.412 ;
      RECT 1.802 6.818 1.87 6.862 ;
      RECT 1.802 6.998 1.87 7.042 ;
      RECT 1.802 7.448 1.87 7.492 ;
      RECT 1.802 9.518 1.87 9.562 ;
      RECT 1.802 9.968 1.87 10.012 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.586 1.958 1.654 2.002 ;
      RECT 1.586 2.408 1.654 2.452 ;
      RECT 1.586 2.588 1.654 2.632 ;
      RECT 1.586 3.038 1.654 3.082 ;
      RECT 1.586 3.218 1.654 3.262 ;
      RECT 1.586 3.668 1.654 3.712 ;
      RECT 1.586 3.848 1.654 3.892 ;
      RECT 1.586 4.298 1.654 4.342 ;
      RECT 1.586 4.478 1.654 4.522 ;
      RECT 1.586 4.928 1.654 4.972 ;
      RECT 1.586 5.108 1.654 5.152 ;
      RECT 1.586 5.558 1.654 5.602 ;
      RECT 1.586 5.738 1.654 5.782 ;
      RECT 1.586 6.188 1.654 6.232 ;
      RECT 1.586 6.368 1.654 6.412 ;
      RECT 1.586 6.818 1.654 6.862 ;
      RECT 1.586 6.998 1.654 7.042 ;
      RECT 1.586 7.448 1.654 7.492 ;
      RECT 1.586 7.628 1.654 7.672 ;
      RECT 1.586 8.078 1.654 8.122 ;
      RECT 1.586 9.518 1.654 9.562 ;
      RECT 1.586 9.968 1.654 10.012 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.37 1.958 1.438 2.002 ;
      RECT 1.37 2.408 1.438 2.452 ;
      RECT 1.37 2.588 1.438 2.632 ;
      RECT 1.37 3.038 1.438 3.082 ;
      RECT 1.37 3.218 1.438 3.262 ;
      RECT 1.37 3.668 1.438 3.712 ;
      RECT 1.37 3.848 1.438 3.892 ;
      RECT 1.37 4.298 1.438 4.342 ;
      RECT 1.37 4.478 1.438 4.522 ;
      RECT 1.37 4.928 1.438 4.972 ;
      RECT 1.37 5.108 1.438 5.152 ;
      RECT 1.37 5.558 1.438 5.602 ;
      RECT 1.37 5.738 1.438 5.782 ;
      RECT 1.37 6.188 1.438 6.232 ;
      RECT 1.37 6.368 1.438 6.412 ;
      RECT 1.37 6.818 1.438 6.862 ;
      RECT 1.37 6.998 1.438 7.042 ;
      RECT 1.37 7.448 1.438 7.492 ;
      RECT 1.37 7.628 1.438 7.672 ;
      RECT 1.37 8.078 1.438 8.122 ;
      RECT 1.37 9.518 1.438 9.562 ;
      RECT 1.37 9.968 1.438 10.012 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.154 1.328 1.222 1.372 ;
      RECT 1.154 1.778 1.222 1.822 ;
      RECT 1.154 1.958 1.222 2.002 ;
      RECT 1.154 2.408 1.222 2.452 ;
      RECT 1.154 2.588 1.222 2.632 ;
      RECT 1.154 3.038 1.222 3.082 ;
      RECT 1.154 3.218 1.222 3.262 ;
      RECT 1.154 3.668 1.222 3.712 ;
      RECT 1.154 3.848 1.222 3.892 ;
      RECT 1.154 4.298 1.222 4.342 ;
      RECT 1.154 4.478 1.222 4.522 ;
      RECT 1.154 4.928 1.222 4.972 ;
      RECT 1.154 5.108 1.222 5.152 ;
      RECT 1.154 5.558 1.222 5.602 ;
      RECT 1.154 5.738 1.222 5.782 ;
      RECT 1.154 6.188 1.222 6.232 ;
      RECT 1.154 6.368 1.222 6.412 ;
      RECT 1.154 6.818 1.222 6.862 ;
      RECT 1.154 6.998 1.222 7.042 ;
      RECT 1.154 7.448 1.222 7.492 ;
      RECT 1.154 7.628 1.222 7.672 ;
      RECT 1.154 8.078 1.222 8.122 ;
      RECT 1.154 8.258 1.222 8.302 ;
      RECT 1.154 8.708 1.222 8.752 ;
      RECT 1.154 9.518 1.222 9.562 ;
      RECT 1.154 9.968 1.222 10.012 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.938 1.328 1.006 1.372 ;
      RECT 0.938 1.778 1.006 1.822 ;
      RECT 0.938 1.958 1.006 2.002 ;
      RECT 0.938 2.408 1.006 2.452 ;
      RECT 0.938 2.588 1.006 2.632 ;
      RECT 0.938 3.038 1.006 3.082 ;
      RECT 0.938 3.218 1.006 3.262 ;
      RECT 0.938 3.668 1.006 3.712 ;
      RECT 0.938 3.848 1.006 3.892 ;
      RECT 0.938 4.298 1.006 4.342 ;
      RECT 0.938 4.478 1.006 4.522 ;
      RECT 0.938 4.928 1.006 4.972 ;
      RECT 0.938 5.108 1.006 5.152 ;
      RECT 0.938 5.558 1.006 5.602 ;
      RECT 0.938 5.738 1.006 5.782 ;
      RECT 0.938 6.188 1.006 6.232 ;
      RECT 0.938 6.368 1.006 6.412 ;
      RECT 0.938 6.818 1.006 6.862 ;
      RECT 0.938 6.998 1.006 7.042 ;
      RECT 0.938 7.448 1.006 7.492 ;
      RECT 0.938 7.628 1.006 7.672 ;
      RECT 0.938 8.078 1.006 8.122 ;
      RECT 0.938 8.258 1.006 8.302 ;
      RECT 0.938 8.708 1.006 8.752 ;
      RECT 0.938 9.518 1.006 9.562 ;
      RECT 0.938 9.968 1.006 10.012 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.722 0.698 0.79 0.742 ;
      RECT 0.722 1.148 0.79 1.192 ;
      RECT 0.722 1.328 0.79 1.372 ;
      RECT 0.722 1.778 0.79 1.822 ;
      RECT 0.722 1.958 0.79 2.002 ;
      RECT 0.722 2.408 0.79 2.452 ;
      RECT 0.722 2.588 0.79 2.632 ;
      RECT 0.722 3.038 0.79 3.082 ;
      RECT 0.722 3.218 0.79 3.262 ;
      RECT 0.722 3.668 0.79 3.712 ;
      RECT 0.722 3.848 0.79 3.892 ;
      RECT 0.722 4.298 0.79 4.342 ;
      RECT 0.722 4.478 0.79 4.522 ;
      RECT 0.722 4.928 0.79 4.972 ;
      RECT 0.722 5.108 0.79 5.152 ;
      RECT 0.722 5.558 0.79 5.602 ;
      RECT 0.722 5.738 0.79 5.782 ;
      RECT 0.722 6.188 0.79 6.232 ;
      RECT 0.722 6.368 0.79 6.412 ;
      RECT 0.722 6.818 0.79 6.862 ;
      RECT 0.722 6.998 0.79 7.042 ;
      RECT 0.722 7.448 0.79 7.492 ;
      RECT 0.722 7.628 0.79 7.672 ;
      RECT 0.722 8.078 0.79 8.122 ;
      RECT 0.722 8.258 0.79 8.302 ;
      RECT 0.722 8.708 0.79 8.752 ;
      RECT 0.722 8.888 0.79 8.932 ;
      RECT 0.722 9.338 0.79 9.382 ;
      RECT 0.722 9.518 0.79 9.562 ;
      RECT 0.722 9.968 0.79 10.012 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.506 0.698 0.574 0.742 ;
      RECT 0.506 1.148 0.574 1.192 ;
      RECT 0.506 1.328 0.574 1.372 ;
      RECT 0.506 1.778 0.574 1.822 ;
      RECT 0.506 1.958 0.574 2.002 ;
      RECT 0.506 2.408 0.574 2.452 ;
      RECT 0.506 2.588 0.574 2.632 ;
      RECT 0.506 3.038 0.574 3.082 ;
      RECT 0.506 3.218 0.574 3.262 ;
      RECT 0.506 3.668 0.574 3.712 ;
      RECT 0.506 3.848 0.574 3.892 ;
      RECT 0.506 4.298 0.574 4.342 ;
      RECT 0.506 4.478 0.574 4.522 ;
      RECT 0.506 4.928 0.574 4.972 ;
      RECT 0.506 5.108 0.574 5.152 ;
      RECT 0.506 5.558 0.574 5.602 ;
      RECT 0.506 5.738 0.574 5.782 ;
      RECT 0.506 6.188 0.574 6.232 ;
      RECT 0.506 6.368 0.574 6.412 ;
      RECT 0.506 6.818 0.574 6.862 ;
      RECT 0.506 6.998 0.574 7.042 ;
      RECT 0.506 7.448 0.574 7.492 ;
      RECT 0.506 7.628 0.574 7.672 ;
      RECT 0.506 8.078 0.574 8.122 ;
      RECT 0.506 8.258 0.574 8.302 ;
      RECT 0.506 8.708 0.574 8.752 ;
      RECT 0.506 8.888 0.574 8.932 ;
      RECT 0.506 9.338 0.574 9.382 ;
      RECT 0.506 9.518 0.574 9.562 ;
      RECT 0.506 9.968 0.574 10.012 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.29 0.698 0.358 0.742 ;
      RECT 0.29 1.148 0.358 1.192 ;
      RECT 0.29 1.328 0.358 1.372 ;
      RECT 0.29 1.778 0.358 1.822 ;
      RECT 0.29 1.958 0.358 2.002 ;
      RECT 0.29 2.408 0.358 2.452 ;
      RECT 0.29 2.588 0.358 2.632 ;
      RECT 0.29 3.038 0.358 3.082 ;
      RECT 0.29 3.218 0.358 3.262 ;
      RECT 0.29 3.668 0.358 3.712 ;
      RECT 0.29 3.848 0.358 3.892 ;
      RECT 0.29 4.298 0.358 4.342 ;
      RECT 0.29 4.478 0.358 4.522 ;
      RECT 0.29 4.928 0.358 4.972 ;
      RECT 0.29 5.108 0.358 5.152 ;
      RECT 0.29 5.558 0.358 5.602 ;
      RECT 0.29 5.738 0.358 5.782 ;
      RECT 0.29 6.188 0.358 6.232 ;
      RECT 0.29 6.368 0.358 6.412 ;
      RECT 0.29 6.818 0.358 6.862 ;
      RECT 0.29 6.998 0.358 7.042 ;
      RECT 0.29 7.448 0.358 7.492 ;
      RECT 0.29 7.628 0.358 7.672 ;
      RECT 0.29 8.078 0.358 8.122 ;
      RECT 0.29 8.258 0.358 8.302 ;
      RECT 0.29 8.708 0.358 8.752 ;
      RECT 0.29 8.888 0.358 8.932 ;
      RECT 0.29 9.338 0.358 9.382 ;
      RECT 0.29 9.518 0.358 9.562 ;
      RECT 0.29 9.968 0.358 10.012 ;
      RECT 0.074 0.068 0.142 0.112 ;
      RECT 0.074 0.518 0.142 0.562 ;
      RECT 0.074 0.698 0.142 0.742 ;
      RECT 0.074 1.148 0.142 1.192 ;
      RECT 0.074 1.328 0.142 1.372 ;
      RECT 0.074 1.778 0.142 1.822 ;
      RECT 0.074 1.958 0.142 2.002 ;
      RECT 0.074 2.408 0.142 2.452 ;
      RECT 0.074 2.588 0.142 2.632 ;
      RECT 0.074 3.038 0.142 3.082 ;
      RECT 0.074 3.218 0.142 3.262 ;
      RECT 0.074 3.668 0.142 3.712 ;
      RECT 0.074 3.848 0.142 3.892 ;
      RECT 0.074 4.298 0.142 4.342 ;
      RECT 0.074 4.478 0.142 4.522 ;
      RECT 0.074 4.928 0.142 4.972 ;
      RECT 0.074 5.108 0.142 5.152 ;
      RECT 0.074 5.558 0.142 5.602 ;
      RECT 0.074 5.738 0.142 5.782 ;
      RECT 0.074 6.188 0.142 6.232 ;
      RECT 0.074 6.368 0.142 6.412 ;
      RECT 0.074 6.818 0.142 6.862 ;
      RECT 0.074 6.998 0.142 7.042 ;
      RECT 0.074 7.448 0.142 7.492 ;
      RECT 0.074 7.628 0.142 7.672 ;
      RECT 0.074 8.078 0.142 8.122 ;
      RECT 0.074 8.258 0.142 8.302 ;
      RECT 0.074 8.708 0.142 8.752 ;
      RECT 0.074 8.888 0.142 8.932 ;
      RECT 0.074 9.338 0.142 9.382 ;
      RECT 0.074 9.518 0.142 9.562 ;
      RECT 0.074 9.968 0.142 10.012 ;
  END
END b15qfdglban1v00x5

MACRO b15qgbao4an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbao4an1n05x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    ANTENNADIFFAREA 0.0918 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 5.2144445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 5.2144445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.292 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.068 0.592 0.112 ;
      LAYER v1 ;
        RECT 0.078 0.068 0.138 0.112 ;
        RECT 0.51 0.068 0.57 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.506 0.088 0.574 0.132 ;
    END
  END o1
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END d
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
      LAYER v0 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 1.37 0.498 1.438 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
        RECT 1.586 0.088 1.654 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.518 1.688 0.562 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
    LAYER v1 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.158 0.518 1.218 0.562 ;
      RECT 0.51 0.518 0.57 0.562 ;
    LAYER v0 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.068 1.438 0.292 ;
  END
END b15qgbao4an1n05x5

MACRO b15qgbar1an1n04x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbar1an1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.29 0.068 0.358 0.292 ;
    LAYER v0 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.293 0.25 0.337 ;
      RECT 0.074 0.088 0.142 0.132 ;
      RECT 0.074 0.498 0.142 0.542 ;
  END
END b15qgbar1an1n04x5

MACRO b15qgbar1an1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbar1an1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.29 0.068 0.358 0.292 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
    LAYER v0 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.293 0.25 0.337 ;
      RECT 0.074 0.088 0.142 0.132 ;
      RECT 0.074 0.498 0.142 0.542 ;
  END
END b15qgbar1an1n08x5

MACRO b15qgbar1an1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbar1an1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.29 0.068 0.358 0.292 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.586 0.068 1.654 0.292 ;
    LAYER v0 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.293 0.25 0.337 ;
      RECT 0.074 0.088 0.142 0.132 ;
      RECT 0.074 0.498 0.142 0.542 ;
  END
END b15qgbar1an1n16x5

MACRO b15qgbar1an1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbar1an1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.29 0.068 0.358 0.292 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.586 0.068 1.654 0.292 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.666 0.068 2.734 0.292 ;
      RECT 2.774 0.068 2.842 0.562 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 3.098 0.068 3.166 0.292 ;
      RECT 3.206 0.068 3.274 0.562 ;
      RECT 3.314 0.338 3.382 0.562 ;
      RECT 3.314 0.068 3.382 0.292 ;
    LAYER v0 ;
      RECT 3.314 0.088 3.382 0.132 ;
      RECT 3.314 0.498 3.382 0.542 ;
      RECT 3.206 0.293 3.274 0.337 ;
      RECT 3.098 0.088 3.166 0.132 ;
      RECT 3.098 0.498 3.166 0.542 ;
      RECT 2.882 0.088 2.95 0.132 ;
      RECT 2.882 0.498 2.95 0.542 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.666 0.088 2.734 0.132 ;
      RECT 2.666 0.498 2.734 0.542 ;
      RECT 2.45 0.088 2.518 0.132 ;
      RECT 2.45 0.498 2.518 0.542 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.234 0.088 2.302 0.132 ;
      RECT 2.234 0.498 2.302 0.542 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 2.018 0.498 2.086 0.542 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.293 0.25 0.337 ;
      RECT 0.074 0.088 0.142 0.132 ;
      RECT 0.074 0.498 0.142 0.542 ;
  END
END b15qgbar1an1n32x5

MACRO b15qgbar1an1n64x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbar1an1n64x5 0 0 ;
  SIZE 6.912 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.946 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.946 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.29 0.068 0.358 0.292 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.586 0.068 1.654 0.292 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.666 0.068 2.734 0.292 ;
      RECT 2.774 0.068 2.842 0.562 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 3.098 0.068 3.166 0.292 ;
      RECT 3.206 0.068 3.274 0.562 ;
      RECT 3.314 0.338 3.382 0.562 ;
      RECT 3.314 0.068 3.382 0.292 ;
      RECT 3.53 0.338 3.598 0.562 ;
      RECT 3.53 0.068 3.598 0.292 ;
      RECT 3.638 0.068 3.706 0.562 ;
      RECT 3.746 0.338 3.814 0.562 ;
      RECT 3.746 0.068 3.814 0.292 ;
      RECT 3.962 0.338 4.03 0.562 ;
      RECT 3.962 0.068 4.03 0.292 ;
      RECT 4.07 0.068 4.138 0.562 ;
      RECT 4.178 0.338 4.246 0.562 ;
      RECT 4.178 0.068 4.246 0.292 ;
      RECT 4.394 0.338 4.462 0.562 ;
      RECT 4.394 0.068 4.462 0.292 ;
      RECT 4.502 0.068 4.57 0.562 ;
      RECT 4.61 0.338 4.678 0.562 ;
      RECT 4.61 0.068 4.678 0.292 ;
      RECT 4.826 0.338 4.894 0.562 ;
      RECT 4.826 0.068 4.894 0.292 ;
      RECT 4.934 0.068 5.002 0.562 ;
      RECT 5.042 0.338 5.11 0.562 ;
      RECT 5.042 0.068 5.11 0.292 ;
      RECT 5.258 0.338 5.326 0.562 ;
      RECT 5.258 0.068 5.326 0.292 ;
      RECT 5.366 0.068 5.434 0.562 ;
      RECT 5.474 0.338 5.542 0.562 ;
      RECT 5.474 0.068 5.542 0.292 ;
      RECT 5.69 0.338 5.758 0.562 ;
      RECT 5.69 0.068 5.758 0.292 ;
      RECT 5.798 0.068 5.866 0.562 ;
      RECT 5.906 0.338 5.974 0.562 ;
      RECT 5.906 0.068 5.974 0.292 ;
      RECT 6.122 0.338 6.19 0.562 ;
      RECT 6.122 0.068 6.19 0.292 ;
      RECT 6.23 0.068 6.298 0.562 ;
      RECT 6.338 0.338 6.406 0.562 ;
      RECT 6.338 0.068 6.406 0.292 ;
      RECT 6.554 0.338 6.622 0.562 ;
      RECT 6.554 0.068 6.622 0.292 ;
      RECT 6.662 0.068 6.73 0.562 ;
      RECT 6.77 0.338 6.838 0.562 ;
      RECT 6.77 0.068 6.838 0.292 ;
    LAYER v0 ;
      RECT 6.77 0.088 6.838 0.132 ;
      RECT 6.77 0.498 6.838 0.542 ;
      RECT 6.662 0.293 6.73 0.337 ;
      RECT 6.554 0.088 6.622 0.132 ;
      RECT 6.554 0.498 6.622 0.542 ;
      RECT 6.338 0.088 6.406 0.132 ;
      RECT 6.338 0.498 6.406 0.542 ;
      RECT 6.23 0.293 6.298 0.337 ;
      RECT 6.122 0.088 6.19 0.132 ;
      RECT 6.122 0.498 6.19 0.542 ;
      RECT 5.906 0.088 5.974 0.132 ;
      RECT 5.906 0.498 5.974 0.542 ;
      RECT 5.798 0.293 5.866 0.337 ;
      RECT 5.69 0.088 5.758 0.132 ;
      RECT 5.69 0.498 5.758 0.542 ;
      RECT 5.474 0.088 5.542 0.132 ;
      RECT 5.474 0.498 5.542 0.542 ;
      RECT 5.366 0.293 5.434 0.337 ;
      RECT 5.258 0.088 5.326 0.132 ;
      RECT 5.258 0.498 5.326 0.542 ;
      RECT 5.042 0.088 5.11 0.132 ;
      RECT 5.042 0.498 5.11 0.542 ;
      RECT 4.934 0.293 5.002 0.337 ;
      RECT 4.826 0.088 4.894 0.132 ;
      RECT 4.826 0.498 4.894 0.542 ;
      RECT 4.61 0.088 4.678 0.132 ;
      RECT 4.61 0.498 4.678 0.542 ;
      RECT 4.502 0.293 4.57 0.337 ;
      RECT 4.394 0.088 4.462 0.132 ;
      RECT 4.394 0.498 4.462 0.542 ;
      RECT 4.178 0.088 4.246 0.132 ;
      RECT 4.178 0.498 4.246 0.542 ;
      RECT 4.07 0.293 4.138 0.337 ;
      RECT 3.962 0.088 4.03 0.132 ;
      RECT 3.962 0.498 4.03 0.542 ;
      RECT 3.746 0.088 3.814 0.132 ;
      RECT 3.746 0.498 3.814 0.542 ;
      RECT 3.638 0.293 3.706 0.337 ;
      RECT 3.53 0.088 3.598 0.132 ;
      RECT 3.53 0.498 3.598 0.542 ;
      RECT 3.314 0.088 3.382 0.132 ;
      RECT 3.314 0.498 3.382 0.542 ;
      RECT 3.206 0.293 3.274 0.337 ;
      RECT 3.098 0.088 3.166 0.132 ;
      RECT 3.098 0.498 3.166 0.542 ;
      RECT 2.882 0.088 2.95 0.132 ;
      RECT 2.882 0.498 2.95 0.542 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.666 0.088 2.734 0.132 ;
      RECT 2.666 0.498 2.734 0.542 ;
      RECT 2.45 0.088 2.518 0.132 ;
      RECT 2.45 0.498 2.518 0.542 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.234 0.088 2.302 0.132 ;
      RECT 2.234 0.498 2.302 0.542 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 2.018 0.498 2.086 0.542 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.293 0.25 0.337 ;
      RECT 0.074 0.088 0.142 0.132 ;
      RECT 0.074 0.498 0.142 0.542 ;
  END
END b15qgbar1an1n64x5

MACRO b15qgbar1an1n72x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbar1an1n72x5 0 0 ;
  SIZE 7.776 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 7.81 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 7.81 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.29 0.068 0.358 0.292 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.586 0.068 1.654 0.292 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.666 0.068 2.734 0.292 ;
      RECT 2.774 0.068 2.842 0.562 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 3.098 0.068 3.166 0.292 ;
      RECT 3.206 0.068 3.274 0.562 ;
      RECT 3.314 0.338 3.382 0.562 ;
      RECT 3.314 0.068 3.382 0.292 ;
      RECT 3.53 0.338 3.598 0.562 ;
      RECT 3.53 0.068 3.598 0.292 ;
      RECT 3.638 0.068 3.706 0.562 ;
      RECT 3.746 0.338 3.814 0.562 ;
      RECT 3.746 0.068 3.814 0.292 ;
      RECT 3.962 0.338 4.03 0.562 ;
      RECT 3.962 0.068 4.03 0.292 ;
      RECT 4.07 0.068 4.138 0.562 ;
      RECT 4.178 0.338 4.246 0.562 ;
      RECT 4.178 0.068 4.246 0.292 ;
      RECT 4.394 0.338 4.462 0.562 ;
      RECT 4.394 0.068 4.462 0.292 ;
      RECT 4.502 0.068 4.57 0.562 ;
      RECT 4.61 0.338 4.678 0.562 ;
      RECT 4.61 0.068 4.678 0.292 ;
      RECT 4.826 0.338 4.894 0.562 ;
      RECT 4.826 0.068 4.894 0.292 ;
      RECT 4.934 0.068 5.002 0.562 ;
      RECT 5.042 0.338 5.11 0.562 ;
      RECT 5.042 0.068 5.11 0.292 ;
      RECT 5.258 0.338 5.326 0.562 ;
      RECT 5.258 0.068 5.326 0.292 ;
      RECT 5.366 0.068 5.434 0.562 ;
      RECT 5.474 0.338 5.542 0.562 ;
      RECT 5.474 0.068 5.542 0.292 ;
      RECT 5.69 0.338 5.758 0.562 ;
      RECT 5.69 0.068 5.758 0.292 ;
      RECT 5.798 0.068 5.866 0.562 ;
      RECT 5.906 0.338 5.974 0.562 ;
      RECT 5.906 0.068 5.974 0.292 ;
      RECT 6.122 0.338 6.19 0.562 ;
      RECT 6.122 0.068 6.19 0.292 ;
      RECT 6.23 0.068 6.298 0.562 ;
      RECT 6.338 0.338 6.406 0.562 ;
      RECT 6.338 0.068 6.406 0.292 ;
      RECT 6.554 0.338 6.622 0.562 ;
      RECT 6.554 0.068 6.622 0.292 ;
      RECT 6.662 0.068 6.73 0.562 ;
      RECT 6.77 0.338 6.838 0.562 ;
      RECT 6.77 0.068 6.838 0.292 ;
      RECT 6.986 0.338 7.054 0.562 ;
      RECT 6.986 0.068 7.054 0.292 ;
      RECT 7.094 0.068 7.162 0.562 ;
      RECT 7.202 0.338 7.27 0.562 ;
      RECT 7.202 0.068 7.27 0.292 ;
      RECT 7.418 0.338 7.486 0.562 ;
      RECT 7.418 0.068 7.486 0.292 ;
      RECT 7.526 0.068 7.594 0.562 ;
      RECT 7.634 0.338 7.702 0.562 ;
      RECT 7.634 0.068 7.702 0.292 ;
    LAYER v0 ;
      RECT 7.634 0.088 7.702 0.132 ;
      RECT 7.634 0.498 7.702 0.542 ;
      RECT 7.526 0.293 7.594 0.337 ;
      RECT 7.418 0.088 7.486 0.132 ;
      RECT 7.418 0.498 7.486 0.542 ;
      RECT 7.202 0.088 7.27 0.132 ;
      RECT 7.202 0.498 7.27 0.542 ;
      RECT 7.094 0.293 7.162 0.337 ;
      RECT 6.986 0.088 7.054 0.132 ;
      RECT 6.986 0.498 7.054 0.542 ;
      RECT 6.77 0.088 6.838 0.132 ;
      RECT 6.77 0.498 6.838 0.542 ;
      RECT 6.662 0.293 6.73 0.337 ;
      RECT 6.554 0.088 6.622 0.132 ;
      RECT 6.554 0.498 6.622 0.542 ;
      RECT 6.338 0.088 6.406 0.132 ;
      RECT 6.338 0.498 6.406 0.542 ;
      RECT 6.23 0.293 6.298 0.337 ;
      RECT 6.122 0.088 6.19 0.132 ;
      RECT 6.122 0.498 6.19 0.542 ;
      RECT 5.906 0.088 5.974 0.132 ;
      RECT 5.906 0.498 5.974 0.542 ;
      RECT 5.798 0.293 5.866 0.337 ;
      RECT 5.69 0.088 5.758 0.132 ;
      RECT 5.69 0.498 5.758 0.542 ;
      RECT 5.474 0.088 5.542 0.132 ;
      RECT 5.474 0.498 5.542 0.542 ;
      RECT 5.366 0.293 5.434 0.337 ;
      RECT 5.258 0.088 5.326 0.132 ;
      RECT 5.258 0.498 5.326 0.542 ;
      RECT 5.042 0.088 5.11 0.132 ;
      RECT 5.042 0.498 5.11 0.542 ;
      RECT 4.934 0.293 5.002 0.337 ;
      RECT 4.826 0.088 4.894 0.132 ;
      RECT 4.826 0.498 4.894 0.542 ;
      RECT 4.61 0.088 4.678 0.132 ;
      RECT 4.61 0.498 4.678 0.542 ;
      RECT 4.502 0.293 4.57 0.337 ;
      RECT 4.394 0.088 4.462 0.132 ;
      RECT 4.394 0.498 4.462 0.542 ;
      RECT 4.178 0.088 4.246 0.132 ;
      RECT 4.178 0.498 4.246 0.542 ;
      RECT 4.07 0.293 4.138 0.337 ;
      RECT 3.962 0.088 4.03 0.132 ;
      RECT 3.962 0.498 4.03 0.542 ;
      RECT 3.746 0.088 3.814 0.132 ;
      RECT 3.746 0.498 3.814 0.542 ;
      RECT 3.638 0.293 3.706 0.337 ;
      RECT 3.53 0.088 3.598 0.132 ;
      RECT 3.53 0.498 3.598 0.542 ;
      RECT 3.314 0.088 3.382 0.132 ;
      RECT 3.314 0.498 3.382 0.542 ;
      RECT 3.206 0.293 3.274 0.337 ;
      RECT 3.098 0.088 3.166 0.132 ;
      RECT 3.098 0.498 3.166 0.542 ;
      RECT 2.882 0.088 2.95 0.132 ;
      RECT 2.882 0.498 2.95 0.542 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.666 0.088 2.734 0.132 ;
      RECT 2.666 0.498 2.734 0.542 ;
      RECT 2.45 0.088 2.518 0.132 ;
      RECT 2.45 0.498 2.518 0.542 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.234 0.088 2.302 0.132 ;
      RECT 2.234 0.498 2.302 0.542 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 2.018 0.498 2.086 0.542 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.182 0.293 0.25 0.337 ;
      RECT 0.074 0.088 0.142 0.132 ;
      RECT 0.074 0.498 0.142 0.542 ;
  END
END b15qgbar1an1n72x5

MACRO b15qgbbd2an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbbd2an1n05x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER m2 ;
        RECT 0.596 0.518 1.132 0.562 ;
      LAYER v1 ;
        RECT 0.618 0.518 0.678 0.562 ;
        RECT 1.05 0.518 1.11 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.088 0.142 0.132 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
        RECT 0.506 0.088 0.574 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.068 1.256 0.112 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.154 0.068 1.222 0.562 ;
    LAYER v1 ;
      RECT 1.158 0.068 1.218 0.112 ;
      RECT 0.186 0.068 0.246 0.112 ;
    LAYER v0 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.182 0.293 0.25 0.337 ;
    LAYER m1 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.338 0.938 0.382 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
  END
END b15qgbbd2an1n05x5

MACRO b15qgbbd4an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbbd4an1n05x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.498 2.518 0.542 ;
        RECT 2.45 0.088 2.518 0.132 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
        RECT 1.37 0.498 1.438 0.542 ;
        RECT 2.234 0.498 2.302 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 1.154 0.088 1.222 0.132 ;
        RECT 1.37 0.088 1.438 0.132 ;
        RECT 2.234 0.088 2.302 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.068 1.132 0.112 ;
      RECT 0.488 0.518 1.996 0.562 ;
      RECT 2 0.068 2.428 0.112 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.068 1.654 0.292 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.018 0.068 2.086 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
    LAYER v1 ;
      RECT 2.346 0.068 2.406 0.112 ;
      RECT 2.022 0.068 2.082 0.112 ;
      RECT 1.914 0.518 1.974 0.562 ;
      RECT 1.482 0.518 1.542 0.562 ;
      RECT 1.05 0.068 1.11 0.112 ;
      RECT 0.618 0.068 0.678 0.112 ;
      RECT 0.51 0.518 0.57 0.562 ;
      RECT 0.294 0.068 0.354 0.112 ;
    LAYER v0 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 2.018 0.498 2.086 0.542 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.338 0.938 0.382 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.654 0.248 1.802 0.292 ;
      RECT 1.802 0.068 1.87 0.292 ;
  END
END b15qgbbd4an1n05x5

MACRO b15qgbbf1an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbbf1an1n05x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.722 0.088 0.79 0.132 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.506 0.088 0.574 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.068 0.7 0.112 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
    LAYER v1 ;
      RECT 0.618 0.068 0.678 0.112 ;
      RECT 0.294 0.068 0.354 0.112 ;
    LAYER v0 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
  END
END b15qgbbf1an1n05x5

MACRO b15qgbbf1an1n15x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbbf1an1n15x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    ANTENNADIFFAREA 0.153 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 1.438 0.562 ;
        RECT 0.938 0.068 1.006 0.562 ;
        RECT 0.722 0.338 1.006 0.382 ;
        RECT 0.722 0.068 0.79 0.562 ;
      LAYER m2 ;
        RECT 0.92 0.428 1.456 0.472 ;
      LAYER v1 ;
        RECT 0.942 0.428 1.002 0.472 ;
        RECT 1.374 0.428 1.434 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 0.938 0.088 1.006 0.132 ;
        RECT 1.37 0.498 1.438 0.542 ;
        RECT 1.37 0.088 1.438 0.132 ;
    END
  END o
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
        RECT 1.586 0.498 1.654 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 1.154 0.088 1.222 0.132 ;
        RECT 1.586 0.088 1.654 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.068 1.564 0.112 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.478 0.068 1.546 0.562 ;
    LAYER v1 ;
      RECT 1.482 0.068 1.542 0.112 ;
      RECT 1.05 0.068 1.11 0.112 ;
      RECT 0.618 0.068 0.678 0.112 ;
      RECT 0.294 0.068 0.354 0.112 ;
    LAYER v0 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.79 0.338 0.938 0.382 ;
      RECT 0.938 0.068 1.006 0.562 ;
  END
END b15qgbbf1an1n15x5

MACRO b15qgbbf1an1n30x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbbf1an1n30x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER m2 ;
        RECT 0.164 0.428 0.7 0.472 ;
      LAYER v1 ;
        RECT 0.186 0.428 0.246 0.472 ;
        RECT 0.618 0.428 0.678 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    ANTENNADIFFAREA 0.2754 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.068 3.166 0.562 ;
        RECT 2.882 0.338 3.166 0.382 ;
        RECT 2.882 0.068 2.95 0.562 ;
        RECT 2.45 0.068 2.518 0.562 ;
        RECT 1.802 0.068 1.87 0.562 ;
        RECT 1.37 0.068 1.438 0.562 ;
        RECT 1.154 0.338 1.438 0.382 ;
        RECT 1.154 0.068 1.222 0.562 ;
      LAYER m2 ;
        RECT 1.352 0.428 2.968 0.472 ;
      LAYER v1 ;
        RECT 1.374 0.428 1.434 0.472 ;
        RECT 1.806 0.428 1.866 0.472 ;
        RECT 2.454 0.428 2.514 0.472 ;
        RECT 2.886 0.428 2.946 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.498 1.222 0.542 ;
        RECT 1.154 0.088 1.222 0.132 ;
        RECT 1.37 0.498 1.438 0.542 ;
        RECT 1.37 0.088 1.438 0.132 ;
        RECT 1.802 0.498 1.87 0.542 ;
        RECT 1.802 0.088 1.87 0.132 ;
        RECT 2.45 0.498 2.518 0.542 ;
        RECT 2.45 0.088 2.518 0.132 ;
        RECT 2.882 0.498 2.95 0.542 ;
        RECT 2.882 0.088 2.95 0.132 ;
        RECT 3.098 0.498 3.166 0.542 ;
        RECT 3.098 0.088 3.166 0.132 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 1.586 0.498 1.654 0.542 ;
        RECT 2.018 0.498 2.086 0.542 ;
        RECT 2.234 0.498 2.302 0.542 ;
        RECT 2.666 0.498 2.734 0.542 ;
        RECT 3.314 0.498 3.382 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 0.938 0.088 1.006 0.132 ;
        RECT 1.586 0.088 1.654 0.132 ;
        RECT 2.018 0.088 2.086 0.132 ;
        RECT 2.234 0.088 2.302 0.132 ;
        RECT 2.666 0.088 2.734 0.132 ;
        RECT 3.314 0.088 3.382 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.068 3.292 0.112 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 2.882 0.068 2.95 0.562 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 2.774 0.068 2.842 0.562 ;
      RECT 3.206 0.068 3.274 0.562 ;
    LAYER v1 ;
      RECT 3.21 0.068 3.27 0.112 ;
      RECT 2.778 0.068 2.838 0.112 ;
      RECT 2.346 0.068 2.406 0.112 ;
      RECT 1.914 0.068 1.974 0.112 ;
      RECT 1.482 0.068 1.542 0.112 ;
      RECT 1.05 0.068 1.11 0.112 ;
      RECT 0.51 0.068 0.57 0.112 ;
    LAYER v0 ;
      RECT 3.206 0.293 3.274 0.337 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 2.95 0.338 3.098 0.382 ;
      RECT 3.098 0.068 3.166 0.562 ;
  END
END b15qgbbf1an1n30x5

MACRO b15qgbdcpan1n04x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbdcpan1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.29 0.498 0.358 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.182 -0.022 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.202 ;
      RECT 0.29 0.068 0.358 0.202 ;
    LAYER v0 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.074 0.088 0.142 0.132 ;
  END
END b15qgbdcpan1n04x5

MACRO b15qgbdcpan1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbdcpan1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 0.722 0.498 0.79 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.382 ;
        RECT 0.182 -0.022 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.202 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.722 0.068 0.79 0.202 ;
    LAYER v0 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.074 0.088 0.142 0.132 ;
  END
END b15qgbdcpan1n08x5

MACRO b15qgbdcpan1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbdcpan1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
        RECT 1.37 0.498 1.438 0.542 ;
        RECT 1.586 0.498 1.654 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.382 ;
        RECT 1.046 -0.022 1.114 0.382 ;
        RECT 0.614 -0.022 0.682 0.382 ;
        RECT 0.182 -0.022 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.614 0.293 0.682 0.337 ;
        RECT 1.046 0.293 1.114 0.337 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.202 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.154 0.068 1.222 0.202 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.586 0.068 1.654 0.202 ;
    LAYER v0 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.074 0.088 0.142 0.132 ;
  END
END b15qgbdcpan1n16x5

MACRO b15qgbdcpan1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbdcpan1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
        RECT 1.37 0.498 1.438 0.542 ;
        RECT 1.586 0.498 1.654 0.542 ;
        RECT 1.802 0.498 1.87 0.542 ;
        RECT 2.018 0.498 2.086 0.542 ;
        RECT 2.234 0.498 2.302 0.542 ;
        RECT 2.45 0.498 2.518 0.542 ;
        RECT 2.666 0.498 2.734 0.542 ;
        RECT 2.882 0.498 2.95 0.542 ;
        RECT 3.098 0.498 3.166 0.542 ;
        RECT 3.314 0.498 3.382 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.206 -0.022 3.274 0.382 ;
        RECT 2.774 -0.022 2.842 0.382 ;
        RECT 2.342 -0.022 2.41 0.382 ;
        RECT 1.91 -0.022 1.978 0.382 ;
        RECT 1.478 -0.022 1.546 0.382 ;
        RECT 1.046 -0.022 1.114 0.382 ;
        RECT 0.614 -0.022 0.682 0.382 ;
        RECT 0.182 -0.022 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.614 0.293 0.682 0.337 ;
        RECT 1.046 0.293 1.114 0.337 ;
        RECT 1.478 0.293 1.546 0.337 ;
        RECT 1.91 0.293 1.978 0.337 ;
        RECT 2.342 0.293 2.41 0.337 ;
        RECT 2.774 0.293 2.842 0.337 ;
        RECT 3.206 0.293 3.274 0.337 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.202 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.154 0.068 1.222 0.202 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.586 0.068 1.654 0.202 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 2.018 0.068 2.086 0.202 ;
      RECT 2.234 0.068 2.302 0.202 ;
      RECT 2.45 0.068 2.518 0.202 ;
      RECT 2.666 0.068 2.734 0.202 ;
      RECT 2.882 0.068 2.95 0.202 ;
      RECT 3.098 0.068 3.166 0.202 ;
      RECT 3.314 0.068 3.382 0.202 ;
    LAYER v0 ;
      RECT 3.314 0.088 3.382 0.132 ;
      RECT 3.098 0.088 3.166 0.132 ;
      RECT 2.882 0.088 2.95 0.132 ;
      RECT 2.666 0.088 2.734 0.132 ;
      RECT 2.45 0.088 2.518 0.132 ;
      RECT 2.234 0.088 2.302 0.132 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.074 0.088 0.142 0.132 ;
  END
END b15qgbdcpan1n32x5

MACRO b15qgbdcpan1n64x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbdcpan1n64x5 0 0 ;
  SIZE 6.912 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.946 0.652 ;
        RECT 6.77 0.428 6.838 0.652 ;
        RECT 6.554 0.428 6.622 0.652 ;
        RECT 6.338 0.428 6.406 0.652 ;
        RECT 6.122 0.428 6.19 0.652 ;
        RECT 5.906 0.428 5.974 0.652 ;
        RECT 5.69 0.428 5.758 0.652 ;
        RECT 5.474 0.428 5.542 0.652 ;
        RECT 5.258 0.428 5.326 0.652 ;
        RECT 5.042 0.428 5.11 0.652 ;
        RECT 4.826 0.428 4.894 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 4.394 0.428 4.462 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
        RECT 1.37 0.498 1.438 0.542 ;
        RECT 1.586 0.498 1.654 0.542 ;
        RECT 1.802 0.498 1.87 0.542 ;
        RECT 2.018 0.498 2.086 0.542 ;
        RECT 2.234 0.498 2.302 0.542 ;
        RECT 2.45 0.498 2.518 0.542 ;
        RECT 2.666 0.498 2.734 0.542 ;
        RECT 2.882 0.498 2.95 0.542 ;
        RECT 3.098 0.498 3.166 0.542 ;
        RECT 3.314 0.498 3.382 0.542 ;
        RECT 3.53 0.498 3.598 0.542 ;
        RECT 3.746 0.498 3.814 0.542 ;
        RECT 3.962 0.498 4.03 0.542 ;
        RECT 4.178 0.498 4.246 0.542 ;
        RECT 4.394 0.498 4.462 0.542 ;
        RECT 4.61 0.498 4.678 0.542 ;
        RECT 4.826 0.498 4.894 0.542 ;
        RECT 5.042 0.498 5.11 0.542 ;
        RECT 5.258 0.498 5.326 0.542 ;
        RECT 5.474 0.498 5.542 0.542 ;
        RECT 5.69 0.498 5.758 0.542 ;
        RECT 5.906 0.498 5.974 0.542 ;
        RECT 6.122 0.498 6.19 0.542 ;
        RECT 6.338 0.498 6.406 0.542 ;
        RECT 6.554 0.498 6.622 0.542 ;
        RECT 6.77 0.498 6.838 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.946 0.022 ;
        RECT 6.662 -0.022 6.73 0.382 ;
        RECT 6.23 -0.022 6.298 0.382 ;
        RECT 5.798 -0.022 5.866 0.382 ;
        RECT 5.366 -0.022 5.434 0.382 ;
        RECT 4.934 -0.022 5.002 0.382 ;
        RECT 4.502 -0.022 4.57 0.382 ;
        RECT 4.07 -0.022 4.138 0.382 ;
        RECT 3.638 -0.022 3.706 0.382 ;
        RECT 3.206 -0.022 3.274 0.382 ;
        RECT 2.774 -0.022 2.842 0.382 ;
        RECT 2.342 -0.022 2.41 0.382 ;
        RECT 1.91 -0.022 1.978 0.382 ;
        RECT 1.478 -0.022 1.546 0.382 ;
        RECT 1.046 -0.022 1.114 0.382 ;
        RECT 0.614 -0.022 0.682 0.382 ;
        RECT 0.182 -0.022 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.614 0.293 0.682 0.337 ;
        RECT 1.046 0.293 1.114 0.337 ;
        RECT 1.478 0.293 1.546 0.337 ;
        RECT 1.91 0.293 1.978 0.337 ;
        RECT 2.342 0.293 2.41 0.337 ;
        RECT 2.774 0.293 2.842 0.337 ;
        RECT 3.206 0.293 3.274 0.337 ;
        RECT 3.638 0.293 3.706 0.337 ;
        RECT 4.07 0.293 4.138 0.337 ;
        RECT 4.502 0.293 4.57 0.337 ;
        RECT 4.934 0.293 5.002 0.337 ;
        RECT 5.366 0.293 5.434 0.337 ;
        RECT 5.798 0.293 5.866 0.337 ;
        RECT 6.23 0.293 6.298 0.337 ;
        RECT 6.662 0.293 6.73 0.337 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.202 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.154 0.068 1.222 0.202 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.586 0.068 1.654 0.202 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 2.018 0.068 2.086 0.202 ;
      RECT 2.234 0.068 2.302 0.202 ;
      RECT 2.45 0.068 2.518 0.202 ;
      RECT 2.666 0.068 2.734 0.202 ;
      RECT 2.882 0.068 2.95 0.202 ;
      RECT 3.098 0.068 3.166 0.202 ;
      RECT 3.314 0.068 3.382 0.202 ;
      RECT 3.53 0.068 3.598 0.202 ;
      RECT 3.746 0.068 3.814 0.202 ;
      RECT 3.962 0.068 4.03 0.202 ;
      RECT 4.178 0.068 4.246 0.202 ;
      RECT 4.394 0.068 4.462 0.202 ;
      RECT 4.61 0.068 4.678 0.202 ;
      RECT 4.826 0.068 4.894 0.202 ;
      RECT 5.042 0.068 5.11 0.202 ;
      RECT 5.258 0.068 5.326 0.202 ;
      RECT 5.474 0.068 5.542 0.202 ;
      RECT 5.69 0.068 5.758 0.202 ;
      RECT 5.906 0.068 5.974 0.202 ;
      RECT 6.122 0.068 6.19 0.202 ;
      RECT 6.338 0.068 6.406 0.202 ;
      RECT 6.554 0.068 6.622 0.202 ;
      RECT 6.77 0.068 6.838 0.202 ;
    LAYER v0 ;
      RECT 6.77 0.088 6.838 0.132 ;
      RECT 6.554 0.088 6.622 0.132 ;
      RECT 6.338 0.088 6.406 0.132 ;
      RECT 6.122 0.088 6.19 0.132 ;
      RECT 5.906 0.088 5.974 0.132 ;
      RECT 5.69 0.088 5.758 0.132 ;
      RECT 5.474 0.088 5.542 0.132 ;
      RECT 5.258 0.088 5.326 0.132 ;
      RECT 5.042 0.088 5.11 0.132 ;
      RECT 4.826 0.088 4.894 0.132 ;
      RECT 4.61 0.088 4.678 0.132 ;
      RECT 4.394 0.088 4.462 0.132 ;
      RECT 4.178 0.088 4.246 0.132 ;
      RECT 3.962 0.088 4.03 0.132 ;
      RECT 3.746 0.088 3.814 0.132 ;
      RECT 3.53 0.088 3.598 0.132 ;
      RECT 3.314 0.088 3.382 0.132 ;
      RECT 3.098 0.088 3.166 0.132 ;
      RECT 2.882 0.088 2.95 0.132 ;
      RECT 2.666 0.088 2.734 0.132 ;
      RECT 2.45 0.088 2.518 0.132 ;
      RECT 2.234 0.088 2.302 0.132 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.074 0.088 0.142 0.132 ;
  END
END b15qgbdcpan1n64x5

MACRO b15qgbdp1an1n00x5
  CLASS CORE ANTENNACELL ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbdp1an1n00x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN dpd1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END dpd1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.29 0.498 0.358 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.182 0.158 0.25 0.562 ;
        RECT 0.074 0.158 0.25 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END vssx
END b15qgbdp1an1n00x5

MACRO b15qgbff4an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbff4an1n05x5 0 0 ;
  SIZE 7.776 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 6.662 0.068 6.73 0.562 ;
        RECT 3.206 0.068 3.274 0.562 ;
      LAYER m2 ;
        RECT 3.188 0.338 6.748 0.382 ;
      LAYER v1 ;
        RECT 3.21 0.338 3.27 0.382 ;
        RECT 6.666 0.338 6.726 0.382 ;
      LAYER v0 ;
        RECT 3.206 0.293 3.274 0.337 ;
        RECT 6.662 0.293 6.73 0.337 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 6.23 0.068 6.298 0.562 ;
        RECT 4.502 0.068 4.57 0.562 ;
      LAYER m2 ;
        RECT 4.484 0.518 6.316 0.562 ;
      LAYER v1 ;
        RECT 4.506 0.518 4.566 0.562 ;
        RECT 6.234 0.518 6.294 0.562 ;
      LAYER v0 ;
        RECT 4.502 0.293 4.57 0.337 ;
        RECT 6.23 0.293 6.298 0.337 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 7.634 0.068 7.702 0.562 ;
      LAYER v0 ;
        RECT 7.634 0.498 7.702 0.542 ;
        RECT 7.634 0.088 7.702 0.132 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 7.81 0.652 ;
        RECT 7.418 0.428 7.486 0.652 ;
        RECT 6.986 0.428 7.054 0.652 ;
        RECT 6.77 0.428 6.838 0.652 ;
        RECT 6.338 0.428 6.406 0.652 ;
        RECT 5.906 0.428 5.974 0.652 ;
        RECT 4.394 0.428 4.462 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
        RECT 1.37 0.498 1.438 0.542 ;
        RECT 2.882 0.498 2.95 0.542 ;
        RECT 3.314 0.498 3.382 0.542 ;
        RECT 3.53 0.498 3.598 0.542 ;
        RECT 4.394 0.498 4.462 0.542 ;
        RECT 5.906 0.498 5.974 0.542 ;
        RECT 6.338 0.498 6.406 0.542 ;
        RECT 6.77 0.498 6.838 0.542 ;
        RECT 6.986 0.498 7.054 0.542 ;
        RECT 7.418 0.498 7.486 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 7.81 0.022 ;
        RECT 7.418 -0.022 7.486 0.202 ;
        RECT 6.554 -0.022 6.622 0.202 ;
        RECT 6.338 -0.022 6.406 0.202 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.53 -0.022 3.598 0.202 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 2.882 -0.022 2.95 0.292 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 1.154 0.088 1.222 0.132 ;
        RECT 1.37 0.088 1.438 0.132 ;
        RECT 2.882 0.088 2.95 0.132 ;
        RECT 3.314 0.088 3.382 0.132 ;
        RECT 3.53 0.088 3.598 0.132 ;
        RECT 4.178 0.088 4.246 0.132 ;
        RECT 6.338 0.088 6.406 0.132 ;
        RECT 6.554 0.088 6.622 0.132 ;
        RECT 7.418 0.088 7.486 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.518 1.564 0.562 ;
      RECT 1.568 0.248 2.552 0.292 ;
      RECT 1.784 0.158 2.752 0.202 ;
      RECT 3.08 0.158 3.848 0.202 ;
      RECT 2.216 0.518 4.156 0.562 ;
      RECT 3.928 0.158 4.48 0.202 ;
      RECT 0.596 0.428 5.036 0.472 ;
      RECT 0.704 0.068 5.452 0.112 ;
      RECT 2.632 0.248 5.56 0.292 ;
      RECT 4.808 0.158 5.884 0.202 ;
      RECT 5.78 0.068 7.288 0.112 ;
      RECT 5.116 0.428 7.736 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.938 0.068 1.006 0.562 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 2.018 0.068 2.086 0.562 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 3.746 0.338 3.814 0.562 ;
      RECT 2.666 0.068 2.734 0.202 ;
      RECT 2.774 0.068 2.842 0.562 ;
      RECT 3.098 0.068 3.166 0.562 ;
      RECT 3.206 0.068 3.274 0.562 ;
      RECT 3.638 0.158 3.706 0.562 ;
      RECT 3.746 0.068 3.814 0.292 ;
      RECT 4.61 0.068 4.678 0.562 ;
      RECT 4.07 0.158 4.138 0.562 ;
      RECT 4.178 0.248 4.246 0.562 ;
      RECT 4.394 0.068 4.462 0.202 ;
      RECT 4.502 0.068 4.57 0.562 ;
      RECT 5.042 0.068 5.11 0.562 ;
      RECT 4.826 0.068 4.894 0.292 ;
      RECT 4.934 0.158 5.002 0.562 ;
      RECT 5.474 0.338 5.542 0.562 ;
      RECT 5.366 0.068 5.434 0.472 ;
      RECT 5.474 0.068 5.542 0.292 ;
      RECT 5.906 0.068 5.974 0.292 ;
      RECT 5.69 0.068 5.758 0.202 ;
      RECT 5.798 0.068 5.866 0.562 ;
      RECT 6.122 0.338 6.19 0.562 ;
      RECT 6.446 0.068 6.514 0.382 ;
      RECT 6.23 0.068 6.298 0.562 ;
      RECT 6.77 0.068 6.838 0.292 ;
      RECT 6.662 0.068 6.73 0.562 ;
      RECT 7.094 0.068 7.162 0.562 ;
      RECT 7.202 0.068 7.27 0.562 ;
      RECT 7.526 0.068 7.594 0.562 ;
    LAYER v1 ;
      RECT 7.53 0.428 7.59 0.472 ;
      RECT 7.206 0.068 7.266 0.112 ;
      RECT 7.098 0.428 7.158 0.472 ;
      RECT 6.45 0.068 6.51 0.112 ;
      RECT 6.126 0.428 6.186 0.472 ;
      RECT 5.802 0.068 5.862 0.112 ;
      RECT 5.694 0.158 5.754 0.202 ;
      RECT 5.478 0.248 5.538 0.292 ;
      RECT 5.37 0.068 5.43 0.112 ;
      RECT 5.262 0.428 5.322 0.472 ;
      RECT 4.938 0.428 4.998 0.472 ;
      RECT 4.83 0.158 4.89 0.202 ;
      RECT 4.614 0.248 4.674 0.292 ;
      RECT 4.398 0.158 4.458 0.202 ;
      RECT 4.182 0.248 4.242 0.292 ;
      RECT 4.074 0.518 4.134 0.562 ;
      RECT 3.966 0.158 4.026 0.202 ;
      RECT 3.642 0.158 3.702 0.202 ;
      RECT 3.102 0.158 3.162 0.202 ;
      RECT 2.778 0.248 2.838 0.292 ;
      RECT 2.67 0.158 2.73 0.202 ;
      RECT 2.454 0.248 2.514 0.292 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.238 0.518 2.298 0.562 ;
      RECT 1.914 0.068 1.974 0.112 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 1.59 0.248 1.65 0.292 ;
      RECT 1.482 0.518 1.542 0.562 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.726 0.068 0.786 0.112 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.294 0.518 0.354 0.562 ;
    LAYER v0 ;
      RECT 7.526 0.293 7.594 0.337 ;
      RECT 7.202 0.088 7.27 0.132 ;
      RECT 7.202 0.498 7.27 0.542 ;
      RECT 7.094 0.293 7.162 0.337 ;
      RECT 6.986 0.088 7.054 0.132 ;
      RECT 6.77 0.088 6.838 0.132 ;
      RECT 6.554 0.498 6.622 0.542 ;
      RECT 6.122 0.088 6.19 0.132 ;
      RECT 6.122 0.498 6.19 0.542 ;
      RECT 5.906 0.088 5.974 0.132 ;
      RECT 5.798 0.293 5.866 0.337 ;
      RECT 5.69 0.088 5.758 0.132 ;
      RECT 5.69 0.498 5.758 0.542 ;
      RECT 5.474 0.088 5.542 0.132 ;
      RECT 5.474 0.498 5.542 0.542 ;
      RECT 5.366 0.293 5.434 0.337 ;
      RECT 5.258 0.088 5.326 0.132 ;
      RECT 5.258 0.498 5.326 0.542 ;
      RECT 5.042 0.088 5.11 0.132 ;
      RECT 5.042 0.498 5.11 0.542 ;
      RECT 4.934 0.293 5.002 0.337 ;
      RECT 4.826 0.088 4.894 0.132 ;
      RECT 4.826 0.498 4.894 0.542 ;
      RECT 4.61 0.088 4.678 0.132 ;
      RECT 4.61 0.498 4.678 0.542 ;
      RECT 4.394 0.088 4.462 0.132 ;
      RECT 4.178 0.498 4.246 0.542 ;
      RECT 4.07 0.293 4.138 0.337 ;
      RECT 3.962 0.088 4.03 0.132 ;
      RECT 3.962 0.498 4.03 0.542 ;
      RECT 3.746 0.088 3.814 0.132 ;
      RECT 3.746 0.498 3.814 0.542 ;
      RECT 3.638 0.293 3.706 0.337 ;
      RECT 3.098 0.088 3.166 0.132 ;
      RECT 3.098 0.498 3.166 0.542 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.666 0.088 2.734 0.132 ;
      RECT 2.666 0.498 2.734 0.542 ;
      RECT 2.45 0.088 2.518 0.132 ;
      RECT 2.45 0.498 2.518 0.542 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.234 0.088 2.302 0.132 ;
      RECT 2.234 0.498 2.302 0.542 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 2.018 0.498 2.086 0.542 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 2.086 0.338 2.234 0.382 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.518 0.338 2.666 0.382 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 3.814 0.338 3.962 0.382 ;
      RECT 3.962 0.338 4.03 0.562 ;
      RECT 3.814 0.248 3.962 0.292 ;
      RECT 3.962 0.068 4.03 0.292 ;
      RECT 4.678 0.338 4.826 0.382 ;
      RECT 4.826 0.338 4.894 0.562 ;
      RECT 5.11 0.338 5.258 0.382 ;
      RECT 5.258 0.068 5.326 0.562 ;
      RECT 5.542 0.338 5.69 0.382 ;
      RECT 5.69 0.338 5.758 0.562 ;
      RECT 5.974 0.248 6.122 0.292 ;
      RECT 6.122 0.068 6.19 0.292 ;
      RECT 6.514 0.338 6.554 0.382 ;
      RECT 6.554 0.338 6.622 0.562 ;
      RECT 6.838 0.248 6.986 0.292 ;
      RECT 6.986 0.068 7.054 0.292 ;
  END
END b15qgbff4an1n05x5

MACRO b15qgbin1an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbin1an1n05x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
    END
  END vssx
END b15qgbin1an1n05x5

MACRO b15qgbin1an1n15x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbin1an1n15x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER m2 ;
        RECT 0.164 0.068 1.132 0.112 ;
      LAYER v1 ;
        RECT 0.186 0.068 0.246 0.112 ;
        RECT 0.618 0.068 0.678 0.112 ;
        RECT 1.05 0.068 1.11 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.614 0.293 0.682 0.337 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    ANTENNADIFFAREA 0.153 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.562 ;
        RECT 0.506 0.068 0.574 0.562 ;
        RECT 0.29 0.338 0.574 0.382 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.518 1.024 0.562 ;
      LAYER v1 ;
        RECT 0.51 0.518 0.57 0.562 ;
        RECT 0.942 0.518 1.002 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.088 0.358 0.132 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 0.938 0.088 1.006 0.132 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 1.154 0.088 1.222 0.132 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.938 0.068 1.006 0.562 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.068 0.574 0.562 ;
  END
END b15qgbin1an1n15x5

MACRO b15qgbin1an1n40x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbin1an1n40x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.068 3.274 0.562 ;
        RECT 2.774 0.068 2.842 0.562 ;
        RECT 2.342 0.068 2.41 0.562 ;
        RECT 1.91 0.068 1.978 0.562 ;
        RECT 1.478 0.068 1.546 0.562 ;
        RECT 1.046 0.068 1.114 0.562 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER m2 ;
        RECT 0.164 0.518 3.292 0.562 ;
      LAYER v1 ;
        RECT 0.186 0.518 0.246 0.562 ;
        RECT 0.618 0.518 0.678 0.562 ;
        RECT 1.05 0.518 1.11 0.562 ;
        RECT 1.482 0.518 1.542 0.562 ;
        RECT 1.914 0.518 1.974 0.562 ;
        RECT 2.346 0.518 2.406 0.562 ;
        RECT 2.778 0.518 2.838 0.562 ;
        RECT 3.21 0.518 3.27 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.614 0.293 0.682 0.337 ;
        RECT 1.046 0.293 1.114 0.337 ;
        RECT 1.478 0.293 1.546 0.337 ;
        RECT 1.91 0.293 1.978 0.337 ;
        RECT 2.342 0.293 2.41 0.337 ;
        RECT 2.774 0.293 2.842 0.337 ;
        RECT 3.206 0.293 3.274 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    ANTENNADIFFAREA 0.3672 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.919111 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.919111 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.068 3.166 0.562 ;
        RECT 2.882 0.338 3.166 0.382 ;
        RECT 2.882 0.068 2.95 0.562 ;
        RECT 2.234 0.068 2.302 0.562 ;
        RECT 2.018 0.338 2.302 0.382 ;
        RECT 2.018 0.068 2.086 0.562 ;
        RECT 1.37 0.068 1.438 0.562 ;
        RECT 1.154 0.338 1.438 0.382 ;
        RECT 1.154 0.068 1.222 0.562 ;
        RECT 0.506 0.068 0.574 0.562 ;
        RECT 0.29 0.338 0.574 0.382 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER m2 ;
        RECT 0.272 0.068 2.968 0.112 ;
      LAYER v1 ;
        RECT 0.294 0.068 0.354 0.112 ;
        RECT 0.51 0.068 0.57 0.112 ;
        RECT 1.158 0.068 1.218 0.112 ;
        RECT 1.374 0.068 1.434 0.112 ;
        RECT 2.022 0.068 2.082 0.112 ;
        RECT 2.238 0.068 2.298 0.112 ;
        RECT 2.886 0.068 2.946 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.088 0.358 0.132 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 1.154 0.498 1.222 0.542 ;
        RECT 1.154 0.088 1.222 0.132 ;
        RECT 1.37 0.498 1.438 0.542 ;
        RECT 1.37 0.088 1.438 0.132 ;
        RECT 2.018 0.498 2.086 0.542 ;
        RECT 2.018 0.088 2.086 0.132 ;
        RECT 2.234 0.498 2.302 0.542 ;
        RECT 2.234 0.088 2.302 0.132 ;
        RECT 2.882 0.498 2.95 0.542 ;
        RECT 2.882 0.088 2.95 0.132 ;
        RECT 3.098 0.498 3.166 0.542 ;
        RECT 3.098 0.088 3.166 0.132 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.314 0.338 3.382 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.586 0.338 1.654 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 1.586 0.498 1.654 0.542 ;
        RECT 1.802 0.498 1.87 0.542 ;
        RECT 2.45 0.498 2.518 0.542 ;
        RECT 2.666 0.498 2.734 0.542 ;
        RECT 3.314 0.498 3.382 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.314 -0.022 3.382 0.292 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 0.938 -0.022 1.006 0.292 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 0.938 0.088 1.006 0.132 ;
        RECT 1.586 0.088 1.654 0.132 ;
        RECT 1.802 0.088 1.87 0.132 ;
        RECT 2.45 0.088 2.518 0.132 ;
        RECT 2.666 0.088 2.734 0.132 ;
        RECT 3.314 0.088 3.382 0.132 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 2.018 0.068 2.086 0.562 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.882 0.068 2.95 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.774 0.068 2.842 0.562 ;
      RECT 3.206 0.068 3.274 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 2.086 0.338 2.234 0.382 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.95 0.338 3.098 0.382 ;
      RECT 3.098 0.068 3.166 0.562 ;
  END
END b15qgbin1an1n40x5

MACRO b15qgblf4an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgblf4an1n05x5 0 0 ;
  SIZE 3.888 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER m2 ;
        RECT 0.596 0.158 1.148 0.202 ;
      LAYER v1 ;
        RECT 0.618 0.158 0.678 0.202 ;
        RECT 1.05 0.158 1.11 0.202 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.068 3.814 0.562 ;
      LAYER v0 ;
        RECT 3.746 0.498 3.814 0.542 ;
        RECT 3.746 0.088 3.814 0.132 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.068 3.274 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.293 3.274 0.337 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.922 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.098 0.338 3.166 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 2.018 0.498 2.086 0.542 ;
        RECT 2.45 0.498 2.518 0.542 ;
        RECT 2.882 0.498 2.95 0.542 ;
        RECT 3.098 0.498 3.166 0.542 ;
        RECT 3.53 0.498 3.598 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.922 0.022 ;
        RECT 3.53 -0.022 3.598 0.202 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.938 0.088 1.006 0.132 ;
        RECT 2.45 0.088 2.518 0.132 ;
        RECT 3.314 0.088 3.382 0.132 ;
        RECT 3.53 0.088 3.598 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.068 0.608 0.112 ;
      RECT 0.04 0.518 1.456 0.562 ;
      RECT 1.228 0.158 1.564 0.202 ;
      RECT 0.688 0.068 1.996 0.112 ;
      RECT 1.784 0.518 2.86 0.562 ;
      RECT 0.488 0.248 3.848 0.292 ;
    LAYER m1 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.29 0.068 0.358 0.292 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 2.666 0.068 2.734 0.562 ;
      RECT 2.774 0.068 2.842 0.562 ;
      RECT 3.314 0.248 3.382 0.562 ;
      RECT 3.638 0.068 3.706 0.562 ;
    LAYER v1 ;
      RECT 3.642 0.248 3.702 0.292 ;
      RECT 3.426 0.248 3.486 0.292 ;
      RECT 2.778 0.518 2.838 0.562 ;
      RECT 2.67 0.248 2.73 0.292 ;
      RECT 2.238 0.518 2.298 0.562 ;
      RECT 1.914 0.068 1.974 0.112 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.59 0.068 1.65 0.112 ;
      RECT 1.482 0.158 1.542 0.202 ;
      RECT 1.374 0.248 1.434 0.292 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 0.726 0.068 0.786 0.112 ;
      RECT 0.51 0.068 0.57 0.112 ;
      RECT 0.51 0.248 0.57 0.292 ;
      RECT 0.294 0.068 0.354 0.112 ;
      RECT 0.294 0.518 0.354 0.562 ;
    LAYER v0 ;
      RECT 3.638 0.293 3.706 0.337 ;
      RECT 3.314 0.498 3.382 0.542 ;
      RECT 3.098 0.088 3.166 0.132 ;
      RECT 2.882 0.088 2.95 0.132 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.666 0.088 2.734 0.132 ;
      RECT 2.666 0.498 2.734 0.542 ;
      RECT 2.234 0.088 2.302 0.132 ;
      RECT 2.234 0.498 2.302 0.542 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.222 0.158 1.33 0.202 ;
      RECT 2.086 0.248 2.234 0.292 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.95 0.248 3.098 0.292 ;
      RECT 3.098 0.068 3.166 0.292 ;
      RECT 3.382 0.248 3.422 0.292 ;
      RECT 3.422 0.068 3.49 0.292 ;
  END
END b15qgblf4an1n05x5

MACRO b15qgbmx2an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbmx2an1n05x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER m2 ;
        RECT 0.164 0.518 1.256 0.562 ;
      LAYER v1 ;
        RECT 0.186 0.518 0.246 0.562 ;
        RECT 1.05 0.518 1.11 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END sa
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.293 1.978 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.498 2.518 0.542 ;
        RECT 2.45 0.088 2.518 0.132 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 2.018 0.498 2.086 0.542 ;
        RECT 2.234 0.498 2.302 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 2.018 0.088 2.086 0.132 ;
        RECT 2.234 0.088 2.302 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.068 1.564 0.112 ;
      RECT 0.704 0.338 1.672 0.382 ;
      RECT 0.92 0.428 1.888 0.472 ;
      RECT 1.336 0.518 2.428 0.562 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.586 0.068 1.654 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
    LAYER v1 ;
      RECT 2.346 0.518 2.406 0.562 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.482 0.068 1.542 0.112 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.294 0.068 0.354 0.112 ;
    LAYER v0 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.654 0.248 1.802 0.292 ;
      RECT 1.802 0.068 1.87 0.562 ;
  END
END b15qgbmx2an1n05x5

MACRO b15qgbmx2an1n10x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbmx2an1n10x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER m2 ;
        RECT 0.164 0.518 1.256 0.562 ;
      LAYER v1 ;
        RECT 0.186 0.518 0.246 0.562 ;
        RECT 1.05 0.518 1.11 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END sa
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.293 1.978 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.562 ;
        RECT 2.45 0.338 2.734 0.382 ;
        RECT 2.45 0.068 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.498 2.518 0.542 ;
        RECT 2.45 0.088 2.518 0.132 ;
        RECT 2.666 0.498 2.734 0.542 ;
        RECT 2.666 0.088 2.734 0.132 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 2.018 0.498 2.086 0.542 ;
        RECT 2.234 0.498 2.302 0.542 ;
        RECT 2.882 0.498 2.95 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 2.018 0.088 2.086 0.132 ;
        RECT 2.234 0.088 2.302 0.132 ;
        RECT 2.882 0.088 2.95 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.068 1.564 0.112 ;
      RECT 0.704 0.338 1.672 0.382 ;
      RECT 0.92 0.428 1.888 0.472 ;
      RECT 1.336 0.518 2.86 0.562 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.586 0.068 1.654 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.774 0.068 2.842 0.562 ;
    LAYER v1 ;
      RECT 2.778 0.518 2.838 0.562 ;
      RECT 2.346 0.518 2.406 0.562 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.482 0.068 1.542 0.112 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.294 0.068 0.354 0.112 ;
    LAYER v0 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.654 0.248 1.802 0.292 ;
      RECT 1.802 0.068 1.87 0.562 ;
  END
END b15qgbmx2an1n10x5

MACRO b15qgbna2an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbna2an1n05x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    ANTENNADIFFAREA 0.0918 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 5.2144445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 5.2144445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.428 0.592 0.472 ;
      LAYER v1 ;
        RECT 0.078 0.428 0.138 0.472 ;
        RECT 0.51 0.428 0.57 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END o1
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.722 0.498 0.79 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.088 0.79 0.132 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.506 0.338 0.574 0.562 ;
    LAYER v0 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.29 0.088 0.358 0.132 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.292 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
  END
END b15qgbna2an1n05x5

MACRO b15qgbna2an1n10x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbna2an1n10x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER m2 ;
        RECT 0.164 0.518 0.7 0.562 ;
      LAYER v1 ;
        RECT 0.186 0.518 0.246 0.562 ;
        RECT 0.618 0.518 0.678 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.562 ;
        RECT 1.046 0.068 1.114 0.562 ;
      LAYER m2 ;
        RECT 1.028 0.518 1.564 0.562 ;
      LAYER v1 ;
        RECT 1.05 0.518 1.11 0.562 ;
        RECT 1.482 0.518 1.542 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    ANTENNADIFFAREA 0.1377 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.338 1.438 0.562 ;
        RECT 1.154 0.338 1.438 0.382 ;
        RECT 1.154 0.338 1.222 0.562 ;
        RECT 0.506 0.068 0.574 0.562 ;
        RECT 0.29 0.248 0.574 0.292 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.428 1.24 0.472 ;
      LAYER v1 ;
        RECT 0.51 0.428 0.57 0.472 ;
        RECT 1.158 0.428 1.218 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.088 0.358 0.132 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 1.154 0.498 1.222 0.542 ;
        RECT 1.37 0.498 1.438 0.542 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.338 1.654 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 1.586 0.498 1.654 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 0.938 -0.022 1.006 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.088 1.006 0.132 ;
        RECT 1.586 0.088 1.654 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.068 1.24 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
    LAYER v1 ;
      RECT 1.158 0.068 1.218 0.112 ;
      RECT 0.726 0.068 0.786 0.112 ;
      RECT 0.078 0.068 0.138 0.112 ;
    LAYER v0 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.074 0.088 0.142 0.132 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.068 1.438 0.292 ;
  END
END b15qgbna2an1n10x5

MACRO b15qgbna3an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbna3an1n05x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    ANTENNADIFFAREA 0.1071 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 5.5904445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 1.106 LAYER m1 ;
      ANTENNAMAXAREACAR 5.2144445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 1.006 0.562 ;
        RECT 0.722 0.338 1.006 0.382 ;
        RECT 0.722 0.338 0.79 0.562 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.428 0.808 0.472 ;
      LAYER v1 ;
        RECT 0.078 0.428 0.138 0.472 ;
        RECT 0.726 0.428 0.786 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.938 0.498 1.006 0.542 ;
    END
  END o1
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END c
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.088 1.222 0.132 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
    LAYER v0 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.29 0.088 0.358 0.132 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.292 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.79 0.338 0.938 0.382 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
  END
END b15qgbna3an1n05x5

MACRO b15qgbno2an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbno2an1n05x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    ANTENNADIFFAREA 0.0918 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 5.2144445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 5.2144445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.292 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.158 0.592 0.202 ;
      LAYER v1 ;
        RECT 0.078 0.158 0.138 0.202 ;
        RECT 0.51 0.158 0.57 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.506 0.088 0.574 0.132 ;
    END
  END o1
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
      LAYER v0 ;
        RECT 0.722 0.498 0.79 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
        RECT 0.722 0.088 0.79 0.132 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.506 0.068 0.574 0.292 ;
    LAYER v0 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.338 0.574 0.562 ;
  END
END b15qgbno2an1n05x5

MACRO b15qgbno2an1n10x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbno2an1n10x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER m2 ;
        RECT 0.164 0.518 0.7 0.562 ;
      LAYER v1 ;
        RECT 0.186 0.518 0.246 0.562 ;
        RECT 0.618 0.518 0.678 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.562 ;
        RECT 1.046 0.068 1.114 0.562 ;
      LAYER m2 ;
        RECT 1.028 0.518 1.564 0.562 ;
      LAYER v1 ;
        RECT 1.05 0.518 1.11 0.562 ;
        RECT 1.482 0.518 1.542 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    ANTENNADIFFAREA 0.1377 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.438 0.292 ;
        RECT 1.37 0.068 1.438 0.292 ;
        RECT 1.154 0.068 1.222 0.292 ;
        RECT 0.506 0.068 0.574 0.562 ;
        RECT 0.29 0.248 0.574 0.292 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.068 1.24 0.112 ;
      LAYER v1 ;
        RECT 0.51 0.068 0.57 0.112 ;
        RECT 1.158 0.068 1.218 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.088 0.358 0.132 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 1.154 0.088 1.222 0.132 ;
        RECT 1.37 0.088 1.438 0.132 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.338 1.654 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
      LAYER v0 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 1.586 0.498 1.654 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 0.938 -0.022 1.006 0.292 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 0.938 0.088 1.006 0.132 ;
        RECT 1.586 0.088 1.654 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.428 1.24 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
    LAYER v1 ;
      RECT 1.158 0.428 1.218 0.472 ;
      RECT 0.726 0.428 0.786 0.472 ;
      RECT 0.078 0.428 0.138 0.472 ;
    LAYER v0 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.068 1.438 0.292 ;
  END
END b15qgbno2an1n10x5

MACRO b15qgbno3an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbno3an1n05x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    ANTENNADIFFAREA 0.1071 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 1.106 LAYER m1 ;
      ANTENNAMAXAREACAR 5.2144445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 5.5904445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 1.006 0.292 ;
        RECT 0.938 0.068 1.006 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.158 0.808 0.202 ;
      LAYER v1 ;
        RECT 0.078 0.158 0.138 0.202 ;
        RECT 0.726 0.158 0.786 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 0.938 0.088 1.006 0.132 ;
    END
  END o1
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END c
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
      LAYER v0 ;
        RECT 1.154 0.498 1.222 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 1.154 0.088 1.222 0.132 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
    LAYER v0 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.79 0.338 0.938 0.382 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
  END
END b15qgbno3an1n05x5

MACRO b15qgboa4an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgboa4an1n05x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
        RECT 0.29 0.338 0.574 0.382 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.088 0.358 0.132 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.938 0.498 1.006 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 0.938 0.088 1.006 0.132 ;
        RECT 1.586 0.088 1.654 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.158 1.24 0.202 ;
      RECT 0.704 0.428 1.688 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.586 0.338 1.654 0.562 ;
    LAYER v1 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.158 0.158 1.218 0.202 ;
      RECT 0.726 0.158 0.786 0.202 ;
      RECT 0.726 0.428 0.786 0.472 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.074 0.088 0.142 0.132 ;
    LAYER m1 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.068 1.438 0.292 ;
  END
END b15qgboa4an1n05x5

MACRO b15qgbth1an1n00x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbth1an1n00x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.182 0.158 0.25 0.562 ;
        RECT 0.074 0.158 0.25 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.382 0.358 0.562 ;
      RECT 0.29 0.068 0.358 0.112 ;
  END
END b15qgbth1an1n00x5

MACRO b15qgbtl1an1n00x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbtl1an1n00x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.29 0.498 0.358 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.182 0.158 0.25 0.562 ;
        RECT 0.074 0.158 0.25 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.0215 0.358 0.112 ;
  END
END b15qgbtl1an1n00x5

MACRO b15qgbxo2an1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbxo2an1n05x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER m2 ;
        RECT 0.164 0.338 1.132 0.382 ;
      LAYER v1 ;
        RECT 0.186 0.338 0.246 0.382 ;
        RECT 1.05 0.338 1.11 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.562 ;
        RECT 1.91 0.068 1.978 0.562 ;
      LAYER m2 ;
        RECT 1.892 0.428 2.428 0.472 ;
      LAYER v1 ;
        RECT 1.914 0.428 1.974 0.472 ;
        RECT 2.346 0.428 2.406 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.293 1.978 0.337 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.562 ;
        RECT 0.722 0.338 1.006 0.382 ;
        RECT 0.722 0.068 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 0.938 0.088 1.006 0.132 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 1.586 0.498 1.654 0.542 ;
        RECT 2.018 0.498 2.086 0.542 ;
        RECT 2.45 0.498 2.518 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 1.586 0.088 1.654 0.132 ;
        RECT 2.018 0.088 2.086 0.132 ;
        RECT 2.45 0.088 2.518 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.428 0.7 0.472 ;
      RECT 0.488 0.158 1.456 0.202 ;
      RECT 0.38 0.068 2.32 0.112 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
    LAYER v1 ;
      RECT 2.238 0.068 2.298 0.112 ;
      RECT 1.806 0.068 1.866 0.112 ;
      RECT 1.482 0.068 1.542 0.112 ;
      RECT 1.374 0.158 1.434 0.202 ;
      RECT 1.158 0.068 1.218 0.112 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.51 0.158 0.57 0.202 ;
      RECT 0.402 0.068 0.462 0.112 ;
      RECT 0.294 0.428 0.354 0.472 ;
    LAYER v0 ;
      RECT 2.234 0.088 2.302 0.132 ;
      RECT 2.234 0.498 2.302 0.542 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.088 1.438 0.132 ;
      RECT 1.37 0.498 1.438 0.542 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.466 0.338 0.506 0.382 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.068 1.438 0.562 ;
  END
END b15qgbxo2an1n05x5

MACRO b15qgbxo2an1n10x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qgbxo2an1n10x5 0 0 ;
  SIZE 4.32 BY 0.63 ;
  SYMMETRY X ;
  SITE bonuscore ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.562 ;
        RECT 1.478 0.068 1.546 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER m2 ;
        RECT 0.164 0.158 1.996 0.202 ;
      LAYER v1 ;
        RECT 0.186 0.158 0.246 0.202 ;
        RECT 1.482 0.158 1.542 0.202 ;
        RECT 1.914 0.158 1.974 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 1.478 0.293 1.546 0.337 ;
        RECT 1.91 0.293 1.978 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 4.2644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.068 4.138 0.562 ;
        RECT 3.638 0.068 3.706 0.562 ;
        RECT 3.206 0.068 3.274 0.562 ;
      LAYER m2 ;
        RECT 3.188 0.158 4.156 0.202 ;
      LAYER v1 ;
        RECT 3.21 0.158 3.27 0.202 ;
        RECT 3.642 0.158 3.702 0.202 ;
        RECT 4.074 0.158 4.134 0.202 ;
      LAYER v0 ;
        RECT 3.206 0.293 3.274 0.337 ;
        RECT 3.638 0.293 3.706 0.337 ;
        RECT 4.07 0.293 4.138 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    ANTENNADIFFAREA 0.1836 LAYER m2 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.919111 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.482 LAYER m1 ;
      ANTENNAMAXAREACAR 9.6704445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.919111 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.068 2.086 0.562 ;
        RECT 1.37 0.068 1.438 0.562 ;
        RECT 1.154 0.248 1.438 0.292 ;
        RECT 1.154 0.068 1.222 0.562 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.428 2.104 0.472 ;
      LAYER v1 ;
        RECT 0.51 0.428 0.57 0.472 ;
        RECT 1.158 0.428 1.218 0.472 ;
        RECT 1.374 0.428 1.434 0.472 ;
        RECT 2.022 0.428 2.082 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 1.154 0.498 1.222 0.542 ;
        RECT 1.154 0.088 1.222 0.132 ;
        RECT 1.37 0.498 1.438 0.542 ;
        RECT 1.37 0.088 1.438 0.132 ;
        RECT 2.018 0.498 2.086 0.542 ;
        RECT 2.018 0.088 2.086 0.132 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.354 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 2.234 0.498 2.302 0.542 ;
        RECT 2.882 0.498 2.95 0.542 ;
        RECT 3.098 0.498 3.166 0.542 ;
        RECT 3.746 0.498 3.814 0.542 ;
        RECT 4.178 0.498 4.246 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.354 0.022 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 2.234 0.088 2.302 0.132 ;
        RECT 2.882 0.088 2.95 0.132 ;
        RECT 3.098 0.088 3.166 0.132 ;
        RECT 3.746 0.088 3.814 0.132 ;
        RECT 4.178 0.088 4.246 0.132 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.248 1.132 0.292 ;
      RECT 0.92 0.068 2.536 0.112 ;
      RECT 0.92 0.338 4.048 0.382 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 1.802 0.068 1.87 0.382 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.018 0.068 2.086 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 3.314 0.068 3.382 0.562 ;
      RECT 2.774 0.068 2.842 0.562 ;
      RECT 3.206 0.068 3.274 0.562 ;
      RECT 3.638 0.068 3.706 0.562 ;
      RECT 3.962 0.068 4.03 0.562 ;
      RECT 4.07 0.068 4.138 0.562 ;
    LAYER v1 ;
      RECT 3.966 0.338 4.026 0.382 ;
      RECT 3.318 0.338 3.378 0.382 ;
      RECT 2.778 0.338 2.838 0.382 ;
      RECT 2.454 0.068 2.514 0.112 ;
      RECT 2.346 0.338 2.406 0.382 ;
      RECT 1.806 0.338 1.866 0.382 ;
      RECT 1.698 0.068 1.758 0.112 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.05 0.248 1.11 0.292 ;
      RECT 0.942 0.068 1.002 0.112 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.618 0.248 0.678 0.292 ;
      RECT 0.294 0.248 0.354 0.292 ;
    LAYER v0 ;
      RECT 3.962 0.088 4.03 0.132 ;
      RECT 3.962 0.498 4.03 0.542 ;
      RECT 3.53 0.088 3.598 0.132 ;
      RECT 3.53 0.498 3.598 0.542 ;
      RECT 3.314 0.088 3.382 0.132 ;
      RECT 3.314 0.498 3.382 0.542 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.666 0.088 2.734 0.132 ;
      RECT 2.666 0.498 2.734 0.542 ;
      RECT 2.45 0.088 2.518 0.132 ;
      RECT 2.45 0.498 2.518 0.542 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 1.802 0.088 1.87 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.722 0.088 0.79 0.132 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.428 0.938 0.472 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.654 0.428 1.694 0.472 ;
      RECT 1.694 0.068 1.762 0.472 ;
      RECT 1.762 0.428 1.802 0.472 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 2.518 0.338 2.666 0.382 ;
      RECT 2.666 0.068 2.734 0.562 ;
      RECT 3.382 0.338 3.53 0.382 ;
      RECT 3.53 0.068 3.598 0.562 ;
  END
END b15qgbxo2an1n10x5

MACRO b15qolcutan1nm1x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qolcutan1nm1x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
    END
  END a
  PIN b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
    END
  END b
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.202 ;
      RECT 0.29 0.068 0.358 0.202 ;
    LAYER v0 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.182 0.138 0.25 0.182 ;
    LAYER m1 ;
      RECT 0.142 0.3375 0.182 0.3825 ;
      RECT 0.182 0.338 0.358 0.382 ;
      RECT 0.358 0.3375 0.398 0.3825 ;
  END
END b15qolcutan1nm1x5

MACRO b15qolmppan1nm1x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qolmppan1nm1x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.074 0.158 0.466 0.202 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.076 0.408 0.14 0.452 ;
        RECT 0.076 0.268 0.14 0.312 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.4 0.2365 0.464 0.2805 ;
        RECT 0.4 0.088 0.464 0.132 ;
    END
  END a
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
    END
  END vssx
END b15qolmppan1nm1x5

MACRO b15qolspwan1nm1x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15qolspwan1nm1x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.0915 0.142 0.1355 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.29 0.0915 0.358 0.1355 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.358 0.562 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.4945 0.142 0.5385 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.29 0.4945 0.358 0.5385 ;
    END
  END b
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
    END
  END vssx
END b15qolspwan1nm1x5

MACRO b15revid0an1nm1x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15revid0an1nm1x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
        RECT 0.074 0.248 0.25 0.292 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.1135 0.142 0.1575 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.202 ;
    LAYER v0 ;
      RECT 0.182 0.1135 0.25 0.1575 ;
    LAYER m1 ;
      RECT 0.074 0.2015 0.142 0.292 ;
      RECT 0.142 0.248 0.182 0.292 ;
  END
END b15revid0an1nm1x5

MACRO b15revid1an1nm1x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15revid1an1nm1x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.1135 0.25 0.1575 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.1135 0.142 0.1575 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.248 ;
  END
END b15revid1an1nm1x5

MACRO b15tihi00an1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15tihi00an1n03x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.202 ;
  END
END b15tihi00an1n03x5

MACRO b15tilo00an1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15tilo00an1n03x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.182 -0.022 0.25 0.112 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.1115 0.25 0.202 ;
  END
END b15tilo00an1n03x5

MACRO b15ydp151an1n03x5
  CLASS CORE ANTENNACELL ;
  ORIGIN 0 0 ;
  FOREIGN b15ydp151an1n03x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN dpd1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.00306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
    END
  END dpd1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
    END
  END vssx
END b15ydp151an1n03x5

MACRO b15ydp251an1n03x5
  CLASS CORE ANTENNACELL ;
  ORIGIN 0 0 ;
  FOREIGN b15ydp251an1n03x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN dpd1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.00306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END dpd1
  PIN dpd2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.00306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END dpd2
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
    END
  END vssx
END b15ydp251an1n03x5

MACRO b15ygnc01an1d03x5
  CLASS CORE ANTENNACELL ;
  ORIGIN 0 0 ;
  FOREIGN b15ygnc01an1d03x5 0 0 ;
  SIZE 0.324 BY 1.26 ;
  SYMMETRY Y ;
  SITE core ;
  PIN gnac1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.00306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.968 0.25 1.192 ;
      LAYER v0 ;
        RECT 0.182 1.058 0.25 1.102 ;
    END
  END gnac1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.608 0.142 0.742 ;
      LAYER v0 ;
        RECT 0.076 0.678 0.14 0.722 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
        RECT -0.034 1.238 0.358 1.282 ;
        RECT 0.074 1.148 0.142 1.282 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.074 1.168 0.142 1.212 ;
    END
  END vssx
END b15ygnc01an1d03x5

MACRO b15zdcf11an1n04x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf11an1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END vssx
END b15zdcf11an1n04x5

MACRO b15zdcf11an1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf11an1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END vssx
END b15zdcf11an1n08x5

MACRO b15zdcf11an1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf11an1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.654 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.222 0.472 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.382 ;
        RECT 1.37 0.158 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.382 ;
        RECT 1.154 -0.022 1.222 0.382 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.382 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
        RECT 0.938 0.293 1.006 0.337 ;
        RECT 1.154 0.293 1.222 0.337 ;
        RECT 1.37 0.293 1.438 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
    END
  END vssx
END b15zdcf11an1n16x5

MACRO b15zdcf11an1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf11an1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.382 0.472 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.95 0.472 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.518 0.472 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 2.086 0.472 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.654 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.222 0.472 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.316 0.538 3.38 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.314 -0.022 3.382 0.382 ;
        RECT 3.098 0.158 3.382 0.202 ;
        RECT 3.098 -0.022 3.166 0.382 ;
        RECT 2.882 -0.022 2.95 0.382 ;
        RECT 2.666 0.158 2.95 0.202 ;
        RECT 2.666 -0.022 2.734 0.382 ;
        RECT 2.45 -0.022 2.518 0.382 ;
        RECT 2.234 0.158 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.382 ;
        RECT 2.018 -0.022 2.086 0.382 ;
        RECT 1.802 0.158 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.382 ;
        RECT 1.586 -0.022 1.654 0.382 ;
        RECT 1.37 0.158 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.382 ;
        RECT 1.154 -0.022 1.222 0.382 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.382 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
        RECT 0.938 0.293 1.006 0.337 ;
        RECT 1.154 0.293 1.222 0.337 ;
        RECT 1.37 0.293 1.438 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
        RECT 1.802 0.293 1.87 0.337 ;
        RECT 2.018 0.293 2.086 0.337 ;
        RECT 2.234 0.293 2.302 0.337 ;
        RECT 2.45 0.293 2.518 0.337 ;
        RECT 2.666 0.293 2.734 0.337 ;
        RECT 2.882 0.293 2.95 0.337 ;
        RECT 3.098 0.293 3.166 0.337 ;
        RECT 3.314 0.293 3.382 0.337 ;
    END
  END vssx
END b15zdcf11an1n32x5

MACRO b15zdcf11an1n64x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf11an1n64x5 0 0 ;
  SIZE 6.912 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.946 0.652 ;
        RECT 6.77 0.428 6.838 0.652 ;
        RECT 6.554 0.428 6.838 0.472 ;
        RECT 6.554 0.428 6.622 0.652 ;
        RECT 6.338 0.428 6.406 0.652 ;
        RECT 6.122 0.428 6.406 0.472 ;
        RECT 6.122 0.428 6.19 0.652 ;
        RECT 5.906 0.428 5.974 0.652 ;
        RECT 5.69 0.428 5.974 0.472 ;
        RECT 5.69 0.428 5.758 0.652 ;
        RECT 5.474 0.428 5.542 0.652 ;
        RECT 5.258 0.428 5.542 0.472 ;
        RECT 5.258 0.428 5.326 0.652 ;
        RECT 5.042 0.428 5.11 0.652 ;
        RECT 4.826 0.428 5.11 0.472 ;
        RECT 4.826 0.428 4.894 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 4.394 0.428 4.678 0.472 ;
        RECT 4.394 0.428 4.462 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.962 0.428 4.246 0.472 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.53 0.428 3.814 0.472 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.382 0.472 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.95 0.472 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.518 0.472 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 2.086 0.472 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.654 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.222 0.472 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
        RECT 3.638 0.428 3.706 0.472 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 4.07 0.428 4.138 0.472 ;
        RECT 4.18 0.538 4.244 0.582 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 4.502 0.428 4.57 0.472 ;
        RECT 4.612 0.538 4.676 0.582 ;
        RECT 4.828 0.538 4.892 0.582 ;
        RECT 4.934 0.428 5.002 0.472 ;
        RECT 5.044 0.538 5.108 0.582 ;
        RECT 5.26 0.538 5.324 0.582 ;
        RECT 5.366 0.428 5.434 0.472 ;
        RECT 5.476 0.538 5.54 0.582 ;
        RECT 5.692 0.538 5.756 0.582 ;
        RECT 5.798 0.428 5.866 0.472 ;
        RECT 5.908 0.538 5.972 0.582 ;
        RECT 6.124 0.538 6.188 0.582 ;
        RECT 6.23 0.428 6.298 0.472 ;
        RECT 6.34 0.538 6.404 0.582 ;
        RECT 6.556 0.538 6.62 0.582 ;
        RECT 6.662 0.428 6.73 0.472 ;
        RECT 6.772 0.538 6.836 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.946 0.022 ;
        RECT 6.77 -0.022 6.838 0.382 ;
        RECT 6.554 0.158 6.838 0.202 ;
        RECT 6.554 -0.022 6.622 0.382 ;
        RECT 6.338 -0.022 6.406 0.382 ;
        RECT 6.122 0.158 6.406 0.202 ;
        RECT 6.122 -0.022 6.19 0.382 ;
        RECT 5.906 -0.022 5.974 0.382 ;
        RECT 5.69 0.158 5.974 0.202 ;
        RECT 5.69 -0.022 5.758 0.382 ;
        RECT 5.474 -0.022 5.542 0.382 ;
        RECT 5.258 0.158 5.542 0.202 ;
        RECT 5.258 -0.022 5.326 0.382 ;
        RECT 5.042 -0.022 5.11 0.382 ;
        RECT 4.826 0.158 5.11 0.202 ;
        RECT 4.826 -0.022 4.894 0.382 ;
        RECT 4.61 -0.022 4.678 0.382 ;
        RECT 4.394 0.158 4.678 0.202 ;
        RECT 4.394 -0.022 4.462 0.382 ;
        RECT 4.178 -0.022 4.246 0.382 ;
        RECT 3.962 0.158 4.246 0.202 ;
        RECT 3.962 -0.022 4.03 0.382 ;
        RECT 3.746 -0.022 3.814 0.382 ;
        RECT 3.53 0.158 3.814 0.202 ;
        RECT 3.53 -0.022 3.598 0.382 ;
        RECT 3.314 -0.022 3.382 0.382 ;
        RECT 3.098 0.158 3.382 0.202 ;
        RECT 3.098 -0.022 3.166 0.382 ;
        RECT 2.882 -0.022 2.95 0.382 ;
        RECT 2.666 0.158 2.95 0.202 ;
        RECT 2.666 -0.022 2.734 0.382 ;
        RECT 2.45 -0.022 2.518 0.382 ;
        RECT 2.234 0.158 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.382 ;
        RECT 2.018 -0.022 2.086 0.382 ;
        RECT 1.802 0.158 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.382 ;
        RECT 1.586 -0.022 1.654 0.382 ;
        RECT 1.37 0.158 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.382 ;
        RECT 1.154 -0.022 1.222 0.382 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.382 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
        RECT 0.938 0.293 1.006 0.337 ;
        RECT 1.154 0.293 1.222 0.337 ;
        RECT 1.37 0.293 1.438 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
        RECT 1.802 0.293 1.87 0.337 ;
        RECT 2.018 0.293 2.086 0.337 ;
        RECT 2.234 0.293 2.302 0.337 ;
        RECT 2.45 0.293 2.518 0.337 ;
        RECT 2.666 0.293 2.734 0.337 ;
        RECT 2.882 0.293 2.95 0.337 ;
        RECT 3.098 0.293 3.166 0.337 ;
        RECT 3.314 0.293 3.382 0.337 ;
        RECT 3.53 0.293 3.598 0.337 ;
        RECT 3.746 0.293 3.814 0.337 ;
        RECT 3.962 0.293 4.03 0.337 ;
        RECT 4.178 0.293 4.246 0.337 ;
        RECT 4.394 0.293 4.462 0.337 ;
        RECT 4.61 0.293 4.678 0.337 ;
        RECT 4.826 0.293 4.894 0.337 ;
        RECT 5.042 0.293 5.11 0.337 ;
        RECT 5.258 0.293 5.326 0.337 ;
        RECT 5.474 0.293 5.542 0.337 ;
        RECT 5.69 0.293 5.758 0.337 ;
        RECT 5.906 0.293 5.974 0.337 ;
        RECT 6.122 0.293 6.19 0.337 ;
        RECT 6.338 0.293 6.406 0.337 ;
        RECT 6.554 0.293 6.622 0.337 ;
        RECT 6.77 0.293 6.838 0.337 ;
    END
  END vssx
END b15zdcf11an1n64x5

MACRO b15zdcf33an1n04x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf33an1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END vssx
END b15zdcf33an1n04x5

MACRO b15zdcf33an1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf33an1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END vssx
END b15zdcf33an1n08x5

MACRO b15zdcf33an1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf33an1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.654 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.222 0.472 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.382 ;
        RECT 1.37 0.158 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.382 ;
        RECT 1.154 -0.022 1.222 0.382 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.382 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
        RECT 0.938 0.293 1.006 0.337 ;
        RECT 1.154 0.293 1.222 0.337 ;
        RECT 1.37 0.293 1.438 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
    END
  END vssx
END b15zdcf33an1n16x5

MACRO b15zdcf33an1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf33an1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.382 0.472 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.95 0.472 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.518 0.472 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 2.086 0.472 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.654 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.222 0.472 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.316 0.538 3.38 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.314 -0.022 3.382 0.382 ;
        RECT 3.098 0.158 3.382 0.202 ;
        RECT 3.098 -0.022 3.166 0.382 ;
        RECT 2.882 -0.022 2.95 0.382 ;
        RECT 2.666 0.158 2.95 0.202 ;
        RECT 2.666 -0.022 2.734 0.382 ;
        RECT 2.45 -0.022 2.518 0.382 ;
        RECT 2.234 0.158 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.382 ;
        RECT 2.018 -0.022 2.086 0.382 ;
        RECT 1.802 0.158 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.382 ;
        RECT 1.586 -0.022 1.654 0.382 ;
        RECT 1.37 0.158 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.382 ;
        RECT 1.154 -0.022 1.222 0.382 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.382 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
        RECT 0.938 0.293 1.006 0.337 ;
        RECT 1.154 0.293 1.222 0.337 ;
        RECT 1.37 0.293 1.438 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
        RECT 1.802 0.293 1.87 0.337 ;
        RECT 2.018 0.293 2.086 0.337 ;
        RECT 2.234 0.293 2.302 0.337 ;
        RECT 2.45 0.293 2.518 0.337 ;
        RECT 2.666 0.293 2.734 0.337 ;
        RECT 2.882 0.293 2.95 0.337 ;
        RECT 3.098 0.293 3.166 0.337 ;
        RECT 3.314 0.293 3.382 0.337 ;
    END
  END vssx
END b15zdcf33an1n32x5

MACRO b15zdcf33an1n64x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf33an1n64x5 0 0 ;
  SIZE 6.912 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.946 0.652 ;
        RECT 6.77 0.428 6.838 0.652 ;
        RECT 6.554 0.428 6.838 0.472 ;
        RECT 6.554 0.428 6.622 0.652 ;
        RECT 6.338 0.428 6.406 0.652 ;
        RECT 6.122 0.428 6.406 0.472 ;
        RECT 6.122 0.428 6.19 0.652 ;
        RECT 5.906 0.428 5.974 0.652 ;
        RECT 5.69 0.428 5.974 0.472 ;
        RECT 5.69 0.428 5.758 0.652 ;
        RECT 5.474 0.428 5.542 0.652 ;
        RECT 5.258 0.428 5.542 0.472 ;
        RECT 5.258 0.428 5.326 0.652 ;
        RECT 5.042 0.428 5.11 0.652 ;
        RECT 4.826 0.428 5.11 0.472 ;
        RECT 4.826 0.428 4.894 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 4.394 0.428 4.678 0.472 ;
        RECT 4.394 0.428 4.462 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.962 0.428 4.246 0.472 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.53 0.428 3.814 0.472 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.382 0.472 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.95 0.472 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.518 0.472 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 2.086 0.472 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.654 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.222 0.472 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
        RECT 3.638 0.428 3.706 0.472 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 4.07 0.428 4.138 0.472 ;
        RECT 4.18 0.538 4.244 0.582 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 4.502 0.428 4.57 0.472 ;
        RECT 4.612 0.538 4.676 0.582 ;
        RECT 4.828 0.538 4.892 0.582 ;
        RECT 4.934 0.428 5.002 0.472 ;
        RECT 5.044 0.538 5.108 0.582 ;
        RECT 5.26 0.538 5.324 0.582 ;
        RECT 5.366 0.428 5.434 0.472 ;
        RECT 5.476 0.538 5.54 0.582 ;
        RECT 5.692 0.538 5.756 0.582 ;
        RECT 5.798 0.428 5.866 0.472 ;
        RECT 5.908 0.538 5.972 0.582 ;
        RECT 6.124 0.538 6.188 0.582 ;
        RECT 6.23 0.428 6.298 0.472 ;
        RECT 6.34 0.538 6.404 0.582 ;
        RECT 6.556 0.538 6.62 0.582 ;
        RECT 6.662 0.428 6.73 0.472 ;
        RECT 6.772 0.538 6.836 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.946 0.022 ;
        RECT 6.77 -0.022 6.838 0.382 ;
        RECT 6.554 0.158 6.838 0.202 ;
        RECT 6.554 -0.022 6.622 0.382 ;
        RECT 6.338 -0.022 6.406 0.382 ;
        RECT 6.122 0.158 6.406 0.202 ;
        RECT 6.122 -0.022 6.19 0.382 ;
        RECT 5.906 -0.022 5.974 0.382 ;
        RECT 5.69 0.158 5.974 0.202 ;
        RECT 5.69 -0.022 5.758 0.382 ;
        RECT 5.474 -0.022 5.542 0.382 ;
        RECT 5.258 0.158 5.542 0.202 ;
        RECT 5.258 -0.022 5.326 0.382 ;
        RECT 5.042 -0.022 5.11 0.382 ;
        RECT 4.826 0.158 5.11 0.202 ;
        RECT 4.826 -0.022 4.894 0.382 ;
        RECT 4.61 -0.022 4.678 0.382 ;
        RECT 4.394 0.158 4.678 0.202 ;
        RECT 4.394 -0.022 4.462 0.382 ;
        RECT 4.178 -0.022 4.246 0.382 ;
        RECT 3.962 0.158 4.246 0.202 ;
        RECT 3.962 -0.022 4.03 0.382 ;
        RECT 3.746 -0.022 3.814 0.382 ;
        RECT 3.53 0.158 3.814 0.202 ;
        RECT 3.53 -0.022 3.598 0.382 ;
        RECT 3.314 -0.022 3.382 0.382 ;
        RECT 3.098 0.158 3.382 0.202 ;
        RECT 3.098 -0.022 3.166 0.382 ;
        RECT 2.882 -0.022 2.95 0.382 ;
        RECT 2.666 0.158 2.95 0.202 ;
        RECT 2.666 -0.022 2.734 0.382 ;
        RECT 2.45 -0.022 2.518 0.382 ;
        RECT 2.234 0.158 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.382 ;
        RECT 2.018 -0.022 2.086 0.382 ;
        RECT 1.802 0.158 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.382 ;
        RECT 1.586 -0.022 1.654 0.382 ;
        RECT 1.37 0.158 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.382 ;
        RECT 1.154 -0.022 1.222 0.382 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.382 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
        RECT 0.938 0.293 1.006 0.337 ;
        RECT 1.154 0.293 1.222 0.337 ;
        RECT 1.37 0.293 1.438 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
        RECT 1.802 0.293 1.87 0.337 ;
        RECT 2.018 0.293 2.086 0.337 ;
        RECT 2.234 0.293 2.302 0.337 ;
        RECT 2.45 0.293 2.518 0.337 ;
        RECT 2.666 0.293 2.734 0.337 ;
        RECT 2.882 0.293 2.95 0.337 ;
        RECT 3.098 0.293 3.166 0.337 ;
        RECT 3.314 0.293 3.382 0.337 ;
        RECT 3.53 0.293 3.598 0.337 ;
        RECT 3.746 0.293 3.814 0.337 ;
        RECT 3.962 0.293 4.03 0.337 ;
        RECT 4.178 0.293 4.246 0.337 ;
        RECT 4.394 0.293 4.462 0.337 ;
        RECT 4.61 0.293 4.678 0.337 ;
        RECT 4.826 0.293 4.894 0.337 ;
        RECT 5.042 0.293 5.11 0.337 ;
        RECT 5.258 0.293 5.326 0.337 ;
        RECT 5.474 0.293 5.542 0.337 ;
        RECT 5.69 0.293 5.758 0.337 ;
        RECT 5.906 0.293 5.974 0.337 ;
        RECT 6.122 0.293 6.19 0.337 ;
        RECT 6.338 0.293 6.406 0.337 ;
        RECT 6.554 0.293 6.622 0.337 ;
        RECT 6.77 0.293 6.838 0.337 ;
    END
  END vssx
END b15zdcf33an1n64x5

MACRO b15zdcf55an1n04x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf55an1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END vssx
END b15zdcf55an1n04x5

MACRO b15zdcf55an1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf55an1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END vssx
END b15zdcf55an1n08x5

MACRO b15zdcf55an1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf55an1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.654 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.222 0.472 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.382 ;
        RECT 1.37 0.158 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.382 ;
        RECT 1.154 -0.022 1.222 0.382 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.382 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
        RECT 0.938 0.293 1.006 0.337 ;
        RECT 1.154 0.293 1.222 0.337 ;
        RECT 1.37 0.293 1.438 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
    END
  END vssx
END b15zdcf55an1n16x5

MACRO b15zdcf55an1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf55an1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.382 0.472 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.95 0.472 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.518 0.472 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 2.086 0.472 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.654 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.222 0.472 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.316 0.538 3.38 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.314 -0.022 3.382 0.382 ;
        RECT 3.098 0.158 3.382 0.202 ;
        RECT 3.098 -0.022 3.166 0.382 ;
        RECT 2.882 -0.022 2.95 0.382 ;
        RECT 2.666 0.158 2.95 0.202 ;
        RECT 2.666 -0.022 2.734 0.382 ;
        RECT 2.45 -0.022 2.518 0.382 ;
        RECT 2.234 0.158 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.382 ;
        RECT 2.018 -0.022 2.086 0.382 ;
        RECT 1.802 0.158 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.382 ;
        RECT 1.586 -0.022 1.654 0.382 ;
        RECT 1.37 0.158 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.382 ;
        RECT 1.154 -0.022 1.222 0.382 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.382 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
        RECT 0.938 0.293 1.006 0.337 ;
        RECT 1.154 0.293 1.222 0.337 ;
        RECT 1.37 0.293 1.438 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
        RECT 1.802 0.293 1.87 0.337 ;
        RECT 2.018 0.293 2.086 0.337 ;
        RECT 2.234 0.293 2.302 0.337 ;
        RECT 2.45 0.293 2.518 0.337 ;
        RECT 2.666 0.293 2.734 0.337 ;
        RECT 2.882 0.293 2.95 0.337 ;
        RECT 3.098 0.293 3.166 0.337 ;
        RECT 3.314 0.293 3.382 0.337 ;
    END
  END vssx
END b15zdcf55an1n32x5

MACRO b15zdcf55an1n64x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdcf55an1n64x5 0 0 ;
  SIZE 6.912 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.946 0.652 ;
        RECT 6.77 0.428 6.838 0.652 ;
        RECT 6.554 0.428 6.838 0.472 ;
        RECT 6.554 0.428 6.622 0.652 ;
        RECT 6.338 0.428 6.406 0.652 ;
        RECT 6.122 0.428 6.406 0.472 ;
        RECT 6.122 0.428 6.19 0.652 ;
        RECT 5.906 0.428 5.974 0.652 ;
        RECT 5.69 0.428 5.974 0.472 ;
        RECT 5.69 0.428 5.758 0.652 ;
        RECT 5.474 0.428 5.542 0.652 ;
        RECT 5.258 0.428 5.542 0.472 ;
        RECT 5.258 0.428 5.326 0.652 ;
        RECT 5.042 0.428 5.11 0.652 ;
        RECT 4.826 0.428 5.11 0.472 ;
        RECT 4.826 0.428 4.894 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 4.394 0.428 4.678 0.472 ;
        RECT 4.394 0.428 4.462 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.962 0.428 4.246 0.472 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.53 0.428 3.814 0.472 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.382 0.472 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.95 0.472 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.518 0.472 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 2.086 0.472 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.654 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.222 0.472 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
        RECT 3.638 0.428 3.706 0.472 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 4.07 0.428 4.138 0.472 ;
        RECT 4.18 0.538 4.244 0.582 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 4.502 0.428 4.57 0.472 ;
        RECT 4.612 0.538 4.676 0.582 ;
        RECT 4.828 0.538 4.892 0.582 ;
        RECT 4.934 0.428 5.002 0.472 ;
        RECT 5.044 0.538 5.108 0.582 ;
        RECT 5.26 0.538 5.324 0.582 ;
        RECT 5.366 0.428 5.434 0.472 ;
        RECT 5.476 0.538 5.54 0.582 ;
        RECT 5.692 0.538 5.756 0.582 ;
        RECT 5.798 0.428 5.866 0.472 ;
        RECT 5.908 0.538 5.972 0.582 ;
        RECT 6.124 0.538 6.188 0.582 ;
        RECT 6.23 0.428 6.298 0.472 ;
        RECT 6.34 0.538 6.404 0.582 ;
        RECT 6.556 0.538 6.62 0.582 ;
        RECT 6.662 0.428 6.73 0.472 ;
        RECT 6.772 0.538 6.836 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.946 0.022 ;
        RECT 6.77 -0.022 6.838 0.382 ;
        RECT 6.554 0.158 6.838 0.202 ;
        RECT 6.554 -0.022 6.622 0.382 ;
        RECT 6.338 -0.022 6.406 0.382 ;
        RECT 6.122 0.158 6.406 0.202 ;
        RECT 6.122 -0.022 6.19 0.382 ;
        RECT 5.906 -0.022 5.974 0.382 ;
        RECT 5.69 0.158 5.974 0.202 ;
        RECT 5.69 -0.022 5.758 0.382 ;
        RECT 5.474 -0.022 5.542 0.382 ;
        RECT 5.258 0.158 5.542 0.202 ;
        RECT 5.258 -0.022 5.326 0.382 ;
        RECT 5.042 -0.022 5.11 0.382 ;
        RECT 4.826 0.158 5.11 0.202 ;
        RECT 4.826 -0.022 4.894 0.382 ;
        RECT 4.61 -0.022 4.678 0.382 ;
        RECT 4.394 0.158 4.678 0.202 ;
        RECT 4.394 -0.022 4.462 0.382 ;
        RECT 4.178 -0.022 4.246 0.382 ;
        RECT 3.962 0.158 4.246 0.202 ;
        RECT 3.962 -0.022 4.03 0.382 ;
        RECT 3.746 -0.022 3.814 0.382 ;
        RECT 3.53 0.158 3.814 0.202 ;
        RECT 3.53 -0.022 3.598 0.382 ;
        RECT 3.314 -0.022 3.382 0.382 ;
        RECT 3.098 0.158 3.382 0.202 ;
        RECT 3.098 -0.022 3.166 0.382 ;
        RECT 2.882 -0.022 2.95 0.382 ;
        RECT 2.666 0.158 2.95 0.202 ;
        RECT 2.666 -0.022 2.734 0.382 ;
        RECT 2.45 -0.022 2.518 0.382 ;
        RECT 2.234 0.158 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.382 ;
        RECT 2.018 -0.022 2.086 0.382 ;
        RECT 1.802 0.158 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.382 ;
        RECT 1.586 -0.022 1.654 0.382 ;
        RECT 1.37 0.158 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.382 ;
        RECT 1.154 -0.022 1.222 0.382 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.382 ;
        RECT 0.722 -0.022 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.382 ;
        RECT 0.29 -0.022 0.358 0.382 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
        RECT 0.938 0.293 1.006 0.337 ;
        RECT 1.154 0.293 1.222 0.337 ;
        RECT 1.37 0.293 1.438 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
        RECT 1.802 0.293 1.87 0.337 ;
        RECT 2.018 0.293 2.086 0.337 ;
        RECT 2.234 0.293 2.302 0.337 ;
        RECT 2.45 0.293 2.518 0.337 ;
        RECT 2.666 0.293 2.734 0.337 ;
        RECT 2.882 0.293 2.95 0.337 ;
        RECT 3.098 0.293 3.166 0.337 ;
        RECT 3.314 0.293 3.382 0.337 ;
        RECT 3.53 0.293 3.598 0.337 ;
        RECT 3.746 0.293 3.814 0.337 ;
        RECT 3.962 0.293 4.03 0.337 ;
        RECT 4.178 0.293 4.246 0.337 ;
        RECT 4.394 0.293 4.462 0.337 ;
        RECT 4.61 0.293 4.678 0.337 ;
        RECT 4.826 0.293 4.894 0.337 ;
        RECT 5.042 0.293 5.11 0.337 ;
        RECT 5.258 0.293 5.326 0.337 ;
        RECT 5.474 0.293 5.542 0.337 ;
        RECT 5.69 0.293 5.758 0.337 ;
        RECT 5.906 0.293 5.974 0.337 ;
        RECT 6.122 0.293 6.19 0.337 ;
        RECT 6.338 0.293 6.406 0.337 ;
        RECT 6.554 0.293 6.622 0.337 ;
        RECT 6.77 0.293 6.838 0.337 ;
    END
  END vssx
END b15zdcf55an1n64x5

MACRO b15zdnd00an1n01x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd00an1n01x5 0 0 ;
  SIZE 0.108 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.142 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.142 0.022 ;
    END
  END vssx
END b15zdnd00an1n01x5

MACRO b15zdnd00an1n02x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd00an1n02x5 0 0 ;
  SIZE 0.216 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.25 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.25 0.022 ;
    END
  END vssx
END b15zdnd00an1n02x5

MACRO b15zdnd11an1n04x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd11an1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
    END
  END vssx
END b15zdnd11an1n04x5

MACRO b15zdnd11an1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd11an1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
    END
  END vssx
END b15zdnd11an1n08x5

MACRO b15zdnd11an1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd11an1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
    END
  END vssx
END b15zdnd11an1n16x5

MACRO b15zdnd11an1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd11an1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
    END
  END vssx
END b15zdnd11an1n32x5

MACRO b15zdnd11an1n64x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd11an1n64x5 0 0 ;
  SIZE 6.912 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.946 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.946 0.022 ;
    END
  END vssx
END b15zdnd11an1n64x5

MACRO b15zdnd33an1n04x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd33an1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
    END
  END vssx
END b15zdnd33an1n04x5

MACRO b15zdnd33an1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd33an1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
    END
  END vssx
END b15zdnd33an1n08x5

MACRO b15zdnd33an1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd33an1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
    END
  END vssx
END b15zdnd33an1n16x5

MACRO b15zdnd33an1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd33an1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
    END
  END vssx
END b15zdnd33an1n32x5

MACRO b15zdnd33an1n64x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd33an1n64x5 0 0 ;
  SIZE 6.912 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.946 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.946 0.022 ;
    END
  END vssx
END b15zdnd33an1n64x5

MACRO b15zdnd55an1n03x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd55an1n03x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
    END
  END vssx
END b15zdnd55an1n03x5

MACRO b15zdnd55an1n04x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd55an1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
    END
  END vssx
END b15zdnd55an1n04x5

MACRO b15zdnd55an1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd55an1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
    END
  END vssx
END b15zdnd55an1n08x5

MACRO b15zdnd55an1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd55an1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
    END
  END vssx
END b15zdnd55an1n16x5

MACRO b15zdnd55an1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd55an1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
    END
  END vssx
END b15zdnd55an1n32x5

MACRO b15zdnd55an1n64x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnd55an1n64x5 0 0 ;
  SIZE 6.912 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.946 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.946 0.022 ;
    END
  END vssx
END b15zdnd55an1n64x5

MACRO b15zdnf11an1n04x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf11an1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
    LAYER v0 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
  END
END b15zdnf11an1n04x5

MACRO b15zdnf11an1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf11an1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
    LAYER v0 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
  END
END b15zdnf11an1n08x5

MACRO b15zdnf11an1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf11an1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.382 ;
    LAYER v0 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.438 0.158 1.586 0.202 ;
      RECT 1.586 0.068 1.654 0.382 ;
  END
END b15zdnf11an1n16x5

MACRO b15zdnf11an1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf11an1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.382 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.382 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.234 0.068 2.302 0.382 ;
      RECT 2.666 0.428 2.734 0.562 ;
      RECT 2.666 0.068 2.734 0.382 ;
      RECT 3.098 0.428 3.166 0.562 ;
      RECT 3.098 0.068 3.166 0.382 ;
    LAYER v0 ;
      RECT 3.314 0.293 3.382 0.337 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.293 3.166 0.337 ;
      RECT 2.882 0.293 2.95 0.337 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.45 0.293 2.518 0.337 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.438 0.158 1.586 0.202 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.87 0.428 2.018 0.472 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 1.87 0.158 2.018 0.202 ;
      RECT 2.018 0.068 2.086 0.382 ;
      RECT 2.302 0.428 2.45 0.472 ;
      RECT 2.45 0.428 2.518 0.562 ;
      RECT 2.302 0.158 2.45 0.202 ;
      RECT 2.45 0.068 2.518 0.382 ;
      RECT 2.734 0.428 2.882 0.472 ;
      RECT 2.882 0.428 2.95 0.562 ;
      RECT 2.734 0.158 2.882 0.202 ;
      RECT 2.882 0.068 2.95 0.382 ;
      RECT 3.166 0.428 3.314 0.472 ;
      RECT 3.314 0.428 3.382 0.562 ;
      RECT 3.166 0.158 3.314 0.202 ;
      RECT 3.314 0.068 3.382 0.382 ;
  END
END b15zdnf11an1n32x5

MACRO b15zdnf11an1n64x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf11an1n64x5 0 0 ;
  SIZE 6.912 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.946 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.946 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.382 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.382 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.234 0.068 2.302 0.382 ;
      RECT 2.666 0.428 2.734 0.562 ;
      RECT 2.666 0.068 2.734 0.382 ;
      RECT 3.098 0.428 3.166 0.562 ;
      RECT 3.098 0.068 3.166 0.382 ;
      RECT 3.53 0.428 3.598 0.562 ;
      RECT 3.53 0.068 3.598 0.382 ;
      RECT 3.962 0.428 4.03 0.562 ;
      RECT 3.962 0.068 4.03 0.382 ;
      RECT 4.394 0.428 4.462 0.562 ;
      RECT 4.394 0.068 4.462 0.382 ;
      RECT 4.826 0.428 4.894 0.562 ;
      RECT 4.826 0.068 4.894 0.382 ;
      RECT 5.258 0.428 5.326 0.562 ;
      RECT 5.258 0.068 5.326 0.382 ;
      RECT 5.69 0.428 5.758 0.562 ;
      RECT 5.69 0.068 5.758 0.382 ;
      RECT 6.122 0.428 6.19 0.562 ;
      RECT 6.122 0.068 6.19 0.382 ;
      RECT 6.554 0.428 6.622 0.562 ;
      RECT 6.554 0.068 6.622 0.382 ;
    LAYER v0 ;
      RECT 6.77 0.293 6.838 0.337 ;
      RECT 6.662 0.428 6.73 0.472 ;
      RECT 6.554 0.293 6.622 0.337 ;
      RECT 6.338 0.293 6.406 0.337 ;
      RECT 6.23 0.428 6.298 0.472 ;
      RECT 6.122 0.293 6.19 0.337 ;
      RECT 5.906 0.293 5.974 0.337 ;
      RECT 5.798 0.428 5.866 0.472 ;
      RECT 5.69 0.293 5.758 0.337 ;
      RECT 5.474 0.293 5.542 0.337 ;
      RECT 5.366 0.428 5.434 0.472 ;
      RECT 5.258 0.293 5.326 0.337 ;
      RECT 5.042 0.293 5.11 0.337 ;
      RECT 4.934 0.428 5.002 0.472 ;
      RECT 4.826 0.293 4.894 0.337 ;
      RECT 4.61 0.293 4.678 0.337 ;
      RECT 4.502 0.428 4.57 0.472 ;
      RECT 4.394 0.293 4.462 0.337 ;
      RECT 4.178 0.293 4.246 0.337 ;
      RECT 4.07 0.428 4.138 0.472 ;
      RECT 3.962 0.293 4.03 0.337 ;
      RECT 3.746 0.293 3.814 0.337 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.53 0.293 3.598 0.337 ;
      RECT 3.314 0.293 3.382 0.337 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.293 3.166 0.337 ;
      RECT 2.882 0.293 2.95 0.337 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.45 0.293 2.518 0.337 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.438 0.158 1.586 0.202 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.87 0.428 2.018 0.472 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 1.87 0.158 2.018 0.202 ;
      RECT 2.018 0.068 2.086 0.382 ;
      RECT 2.302 0.428 2.45 0.472 ;
      RECT 2.45 0.428 2.518 0.562 ;
      RECT 2.302 0.158 2.45 0.202 ;
      RECT 2.45 0.068 2.518 0.382 ;
      RECT 2.734 0.428 2.882 0.472 ;
      RECT 2.882 0.428 2.95 0.562 ;
      RECT 2.734 0.158 2.882 0.202 ;
      RECT 2.882 0.068 2.95 0.382 ;
      RECT 3.166 0.428 3.314 0.472 ;
      RECT 3.314 0.428 3.382 0.562 ;
      RECT 3.166 0.158 3.314 0.202 ;
      RECT 3.314 0.068 3.382 0.382 ;
      RECT 3.598 0.428 3.746 0.472 ;
      RECT 3.746 0.428 3.814 0.562 ;
      RECT 3.598 0.158 3.746 0.202 ;
      RECT 3.746 0.068 3.814 0.382 ;
      RECT 4.03 0.428 4.178 0.472 ;
      RECT 4.178 0.428 4.246 0.562 ;
      RECT 4.03 0.158 4.178 0.202 ;
      RECT 4.178 0.068 4.246 0.382 ;
      RECT 4.462 0.428 4.61 0.472 ;
      RECT 4.61 0.428 4.678 0.562 ;
      RECT 4.462 0.158 4.61 0.202 ;
      RECT 4.61 0.068 4.678 0.382 ;
      RECT 4.894 0.428 5.042 0.472 ;
      RECT 5.042 0.428 5.11 0.562 ;
      RECT 4.894 0.158 5.042 0.202 ;
      RECT 5.042 0.068 5.11 0.382 ;
      RECT 5.326 0.428 5.474 0.472 ;
      RECT 5.474 0.428 5.542 0.562 ;
      RECT 5.326 0.158 5.474 0.202 ;
      RECT 5.474 0.068 5.542 0.382 ;
      RECT 5.758 0.428 5.906 0.472 ;
      RECT 5.906 0.428 5.974 0.562 ;
      RECT 5.758 0.158 5.906 0.202 ;
      RECT 5.906 0.068 5.974 0.382 ;
      RECT 6.19 0.428 6.338 0.472 ;
      RECT 6.338 0.428 6.406 0.562 ;
      RECT 6.19 0.158 6.338 0.202 ;
      RECT 6.338 0.068 6.406 0.382 ;
      RECT 6.622 0.428 6.77 0.472 ;
      RECT 6.77 0.428 6.838 0.562 ;
      RECT 6.622 0.158 6.77 0.202 ;
      RECT 6.77 0.068 6.838 0.382 ;
  END
END b15zdnf11an1n64x5

MACRO b15zdnf33an1n04x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf33an1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
    LAYER v0 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
  END
END b15zdnf33an1n04x5

MACRO b15zdnf33an1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf33an1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
    LAYER v0 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
  END
END b15zdnf33an1n08x5

MACRO b15zdnf33an1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf33an1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.382 ;
    LAYER v0 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.438 0.158 1.586 0.202 ;
      RECT 1.586 0.068 1.654 0.382 ;
  END
END b15zdnf33an1n16x5

MACRO b15zdnf33an1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf33an1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.382 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.382 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.234 0.068 2.302 0.382 ;
      RECT 2.666 0.428 2.734 0.562 ;
      RECT 2.666 0.068 2.734 0.382 ;
      RECT 3.098 0.428 3.166 0.562 ;
      RECT 3.098 0.068 3.166 0.382 ;
    LAYER v0 ;
      RECT 3.314 0.293 3.382 0.337 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.293 3.166 0.337 ;
      RECT 2.882 0.293 2.95 0.337 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.45 0.293 2.518 0.337 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.438 0.158 1.586 0.202 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.87 0.428 2.018 0.472 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 1.87 0.158 2.018 0.202 ;
      RECT 2.018 0.068 2.086 0.382 ;
      RECT 2.302 0.428 2.45 0.472 ;
      RECT 2.45 0.428 2.518 0.562 ;
      RECT 2.302 0.158 2.45 0.202 ;
      RECT 2.45 0.068 2.518 0.382 ;
      RECT 2.734 0.428 2.882 0.472 ;
      RECT 2.882 0.428 2.95 0.562 ;
      RECT 2.734 0.158 2.882 0.202 ;
      RECT 2.882 0.068 2.95 0.382 ;
      RECT 3.166 0.428 3.314 0.472 ;
      RECT 3.314 0.428 3.382 0.562 ;
      RECT 3.166 0.158 3.314 0.202 ;
      RECT 3.314 0.068 3.382 0.382 ;
  END
END b15zdnf33an1n32x5

MACRO b15zdnf33an1n64x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf33an1n64x5 0 0 ;
  SIZE 6.912 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.946 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.946 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.382 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.382 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.234 0.068 2.302 0.382 ;
      RECT 2.666 0.428 2.734 0.562 ;
      RECT 2.666 0.068 2.734 0.382 ;
      RECT 3.098 0.428 3.166 0.562 ;
      RECT 3.098 0.068 3.166 0.382 ;
      RECT 3.53 0.428 3.598 0.562 ;
      RECT 3.53 0.068 3.598 0.382 ;
      RECT 3.962 0.428 4.03 0.562 ;
      RECT 3.962 0.068 4.03 0.382 ;
      RECT 4.394 0.428 4.462 0.562 ;
      RECT 4.394 0.068 4.462 0.382 ;
      RECT 4.826 0.428 4.894 0.562 ;
      RECT 4.826 0.068 4.894 0.382 ;
      RECT 5.258 0.428 5.326 0.562 ;
      RECT 5.258 0.068 5.326 0.382 ;
      RECT 5.69 0.428 5.758 0.562 ;
      RECT 5.69 0.068 5.758 0.382 ;
      RECT 6.122 0.428 6.19 0.562 ;
      RECT 6.122 0.068 6.19 0.382 ;
      RECT 6.554 0.428 6.622 0.562 ;
      RECT 6.554 0.068 6.622 0.382 ;
    LAYER v0 ;
      RECT 6.77 0.293 6.838 0.337 ;
      RECT 6.662 0.428 6.73 0.472 ;
      RECT 6.554 0.293 6.622 0.337 ;
      RECT 6.338 0.293 6.406 0.337 ;
      RECT 6.23 0.428 6.298 0.472 ;
      RECT 6.122 0.293 6.19 0.337 ;
      RECT 5.906 0.293 5.974 0.337 ;
      RECT 5.798 0.428 5.866 0.472 ;
      RECT 5.69 0.293 5.758 0.337 ;
      RECT 5.474 0.293 5.542 0.337 ;
      RECT 5.366 0.428 5.434 0.472 ;
      RECT 5.258 0.293 5.326 0.337 ;
      RECT 5.042 0.293 5.11 0.337 ;
      RECT 4.934 0.428 5.002 0.472 ;
      RECT 4.826 0.293 4.894 0.337 ;
      RECT 4.61 0.293 4.678 0.337 ;
      RECT 4.502 0.428 4.57 0.472 ;
      RECT 4.394 0.293 4.462 0.337 ;
      RECT 4.178 0.293 4.246 0.337 ;
      RECT 4.07 0.428 4.138 0.472 ;
      RECT 3.962 0.293 4.03 0.337 ;
      RECT 3.746 0.293 3.814 0.337 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.53 0.293 3.598 0.337 ;
      RECT 3.314 0.293 3.382 0.337 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.293 3.166 0.337 ;
      RECT 2.882 0.293 2.95 0.337 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.45 0.293 2.518 0.337 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.438 0.158 1.586 0.202 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.87 0.428 2.018 0.472 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 1.87 0.158 2.018 0.202 ;
      RECT 2.018 0.068 2.086 0.382 ;
      RECT 2.302 0.428 2.45 0.472 ;
      RECT 2.45 0.428 2.518 0.562 ;
      RECT 2.302 0.158 2.45 0.202 ;
      RECT 2.45 0.068 2.518 0.382 ;
      RECT 2.734 0.428 2.882 0.472 ;
      RECT 2.882 0.428 2.95 0.562 ;
      RECT 2.734 0.158 2.882 0.202 ;
      RECT 2.882 0.068 2.95 0.382 ;
      RECT 3.166 0.428 3.314 0.472 ;
      RECT 3.314 0.428 3.382 0.562 ;
      RECT 3.166 0.158 3.314 0.202 ;
      RECT 3.314 0.068 3.382 0.382 ;
      RECT 3.598 0.428 3.746 0.472 ;
      RECT 3.746 0.428 3.814 0.562 ;
      RECT 3.598 0.158 3.746 0.202 ;
      RECT 3.746 0.068 3.814 0.382 ;
      RECT 4.03 0.428 4.178 0.472 ;
      RECT 4.178 0.428 4.246 0.562 ;
      RECT 4.03 0.158 4.178 0.202 ;
      RECT 4.178 0.068 4.246 0.382 ;
      RECT 4.462 0.428 4.61 0.472 ;
      RECT 4.61 0.428 4.678 0.562 ;
      RECT 4.462 0.158 4.61 0.202 ;
      RECT 4.61 0.068 4.678 0.382 ;
      RECT 4.894 0.428 5.042 0.472 ;
      RECT 5.042 0.428 5.11 0.562 ;
      RECT 4.894 0.158 5.042 0.202 ;
      RECT 5.042 0.068 5.11 0.382 ;
      RECT 5.326 0.428 5.474 0.472 ;
      RECT 5.474 0.428 5.542 0.562 ;
      RECT 5.326 0.158 5.474 0.202 ;
      RECT 5.474 0.068 5.542 0.382 ;
      RECT 5.758 0.428 5.906 0.472 ;
      RECT 5.906 0.428 5.974 0.562 ;
      RECT 5.758 0.158 5.906 0.202 ;
      RECT 5.906 0.068 5.974 0.382 ;
      RECT 6.19 0.428 6.338 0.472 ;
      RECT 6.338 0.428 6.406 0.562 ;
      RECT 6.19 0.158 6.338 0.202 ;
      RECT 6.338 0.068 6.406 0.382 ;
      RECT 6.622 0.428 6.77 0.472 ;
      RECT 6.77 0.428 6.838 0.562 ;
      RECT 6.622 0.158 6.77 0.202 ;
      RECT 6.77 0.068 6.838 0.382 ;
  END
END b15zdnf33an1n64x5

MACRO b15zdnf55an1n04x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf55an1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
    LAYER v0 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
  END
END b15zdnf55an1n04x5

MACRO b15zdnf55an1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf55an1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
    LAYER v0 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
  END
END b15zdnf55an1n08x5

MACRO b15zdnf55an1n16x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf55an1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.382 ;
    LAYER v0 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.438 0.158 1.586 0.202 ;
      RECT 1.586 0.068 1.654 0.382 ;
  END
END b15zdnf55an1n16x5

MACRO b15zdnf55an1n32x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf55an1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.382 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.382 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.234 0.068 2.302 0.382 ;
      RECT 2.666 0.428 2.734 0.562 ;
      RECT 2.666 0.068 2.734 0.382 ;
      RECT 3.098 0.428 3.166 0.562 ;
      RECT 3.098 0.068 3.166 0.382 ;
    LAYER v0 ;
      RECT 3.314 0.293 3.382 0.337 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.293 3.166 0.337 ;
      RECT 2.882 0.293 2.95 0.337 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.45 0.293 2.518 0.337 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.438 0.158 1.586 0.202 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.87 0.428 2.018 0.472 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 1.87 0.158 2.018 0.202 ;
      RECT 2.018 0.068 2.086 0.382 ;
      RECT 2.302 0.428 2.45 0.472 ;
      RECT 2.45 0.428 2.518 0.562 ;
      RECT 2.302 0.158 2.45 0.202 ;
      RECT 2.45 0.068 2.518 0.382 ;
      RECT 2.734 0.428 2.882 0.472 ;
      RECT 2.882 0.428 2.95 0.562 ;
      RECT 2.734 0.158 2.882 0.202 ;
      RECT 2.882 0.068 2.95 0.382 ;
      RECT 3.166 0.428 3.314 0.472 ;
      RECT 3.314 0.428 3.382 0.562 ;
      RECT 3.166 0.158 3.314 0.202 ;
      RECT 3.314 0.068 3.382 0.382 ;
  END
END b15zdnf55an1n32x5

MACRO b15zdnf55an1n64x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnf55an1n64x5 0 0 ;
  SIZE 6.912 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.946 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.946 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.382 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.382 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.234 0.068 2.302 0.382 ;
      RECT 2.666 0.428 2.734 0.562 ;
      RECT 2.666 0.068 2.734 0.382 ;
      RECT 3.098 0.428 3.166 0.562 ;
      RECT 3.098 0.068 3.166 0.382 ;
      RECT 3.53 0.428 3.598 0.562 ;
      RECT 3.53 0.068 3.598 0.382 ;
      RECT 3.962 0.428 4.03 0.562 ;
      RECT 3.962 0.068 4.03 0.382 ;
      RECT 4.394 0.428 4.462 0.562 ;
      RECT 4.394 0.068 4.462 0.382 ;
      RECT 4.826 0.428 4.894 0.562 ;
      RECT 4.826 0.068 4.894 0.382 ;
      RECT 5.258 0.428 5.326 0.562 ;
      RECT 5.258 0.068 5.326 0.382 ;
      RECT 5.69 0.428 5.758 0.562 ;
      RECT 5.69 0.068 5.758 0.382 ;
      RECT 6.122 0.428 6.19 0.562 ;
      RECT 6.122 0.068 6.19 0.382 ;
      RECT 6.554 0.428 6.622 0.562 ;
      RECT 6.554 0.068 6.622 0.382 ;
    LAYER v0 ;
      RECT 6.77 0.293 6.838 0.337 ;
      RECT 6.662 0.428 6.73 0.472 ;
      RECT 6.554 0.293 6.622 0.337 ;
      RECT 6.338 0.293 6.406 0.337 ;
      RECT 6.23 0.428 6.298 0.472 ;
      RECT 6.122 0.293 6.19 0.337 ;
      RECT 5.906 0.293 5.974 0.337 ;
      RECT 5.798 0.428 5.866 0.472 ;
      RECT 5.69 0.293 5.758 0.337 ;
      RECT 5.474 0.293 5.542 0.337 ;
      RECT 5.366 0.428 5.434 0.472 ;
      RECT 5.258 0.293 5.326 0.337 ;
      RECT 5.042 0.293 5.11 0.337 ;
      RECT 4.934 0.428 5.002 0.472 ;
      RECT 4.826 0.293 4.894 0.337 ;
      RECT 4.61 0.293 4.678 0.337 ;
      RECT 4.502 0.428 4.57 0.472 ;
      RECT 4.394 0.293 4.462 0.337 ;
      RECT 4.178 0.293 4.246 0.337 ;
      RECT 4.07 0.428 4.138 0.472 ;
      RECT 3.962 0.293 4.03 0.337 ;
      RECT 3.746 0.293 3.814 0.337 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.53 0.293 3.598 0.337 ;
      RECT 3.314 0.293 3.382 0.337 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.293 3.166 0.337 ;
      RECT 2.882 0.293 2.95 0.337 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.45 0.293 2.518 0.337 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.438 0.158 1.586 0.202 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.87 0.428 2.018 0.472 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 1.87 0.158 2.018 0.202 ;
      RECT 2.018 0.068 2.086 0.382 ;
      RECT 2.302 0.428 2.45 0.472 ;
      RECT 2.45 0.428 2.518 0.562 ;
      RECT 2.302 0.158 2.45 0.202 ;
      RECT 2.45 0.068 2.518 0.382 ;
      RECT 2.734 0.428 2.882 0.472 ;
      RECT 2.882 0.428 2.95 0.562 ;
      RECT 2.734 0.158 2.882 0.202 ;
      RECT 2.882 0.068 2.95 0.382 ;
      RECT 3.166 0.428 3.314 0.472 ;
      RECT 3.314 0.428 3.382 0.562 ;
      RECT 3.166 0.158 3.314 0.202 ;
      RECT 3.314 0.068 3.382 0.382 ;
      RECT 3.598 0.428 3.746 0.472 ;
      RECT 3.746 0.428 3.814 0.562 ;
      RECT 3.598 0.158 3.746 0.202 ;
      RECT 3.746 0.068 3.814 0.382 ;
      RECT 4.03 0.428 4.178 0.472 ;
      RECT 4.178 0.428 4.246 0.562 ;
      RECT 4.03 0.158 4.178 0.202 ;
      RECT 4.178 0.068 4.246 0.382 ;
      RECT 4.462 0.428 4.61 0.472 ;
      RECT 4.61 0.428 4.678 0.562 ;
      RECT 4.462 0.158 4.61 0.202 ;
      RECT 4.61 0.068 4.678 0.382 ;
      RECT 4.894 0.428 5.042 0.472 ;
      RECT 5.042 0.428 5.11 0.562 ;
      RECT 4.894 0.158 5.042 0.202 ;
      RECT 5.042 0.068 5.11 0.382 ;
      RECT 5.326 0.428 5.474 0.472 ;
      RECT 5.474 0.428 5.542 0.562 ;
      RECT 5.326 0.158 5.474 0.202 ;
      RECT 5.474 0.068 5.542 0.382 ;
      RECT 5.758 0.428 5.906 0.472 ;
      RECT 5.906 0.428 5.974 0.562 ;
      RECT 5.758 0.158 5.906 0.202 ;
      RECT 5.906 0.068 5.974 0.382 ;
      RECT 6.19 0.428 6.338 0.472 ;
      RECT 6.338 0.428 6.406 0.562 ;
      RECT 6.19 0.158 6.338 0.202 ;
      RECT 6.338 0.068 6.406 0.382 ;
      RECT 6.622 0.428 6.77 0.472 ;
      RECT 6.77 0.428 6.838 0.562 ;
      RECT 6.622 0.158 6.77 0.202 ;
      RECT 6.77 0.068 6.838 0.382 ;
  END
END b15zdnf55an1n64x5

MACRO b15zdnnvian1d03x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnnvian1d03x5 0 0 ;
  SIZE 0.324 BY 1.26 ;
  SYMMETRY Y ;
  SITE core ;
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.202 ;
        RECT -0.034 1.238 0.358 1.282 ;
      LAYER v0 ;
        RECT 0.074 0.118 0.142 0.162 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 1.058 0.142 1.192 ;
    LAYER v0 ;
      RECT 0.074 1.103 0.142 1.147 ;
  END
END b15zdnnvian1d03x5

MACRO b15zdnnvian1n03x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15zdnnvian1n03x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.074 0.068 0.142 0.202 ;
    LAYER v0 ;
      RECT 0.074 0.113 0.142 0.157 ;
      RECT 0.074 0.473 0.142 0.517 ;
  END
END b15zdnnvian1n03x5

MACRO b15ztp015an1n05x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15ztp015an1n05x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.202 ;
    LAYER v0 ;
      RECT 0.182 0.118 0.25 0.162 ;
  END
END b15ztp015an1n05x5

MACRO b15ztp051an1n05x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15ztp051an1n05x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.428 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.182 0.473 0.25 0.517 ;
  END
END b15ztp051an1n05x5

MACRO b15ztpn00an1d03x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15ztpn00an1d03x5 0 0 ;
  SIZE 0.324 BY 1.26 ;
  SYMMETRY Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.608 0.142 0.832 ;
      LAYER v0 ;
        RECT 0.076 0.678 0.14 0.722 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
        RECT -0.034 1.238 0.358 1.282 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 1.058 0.142 1.192 ;
    LAYER v0 ;
      RECT 0.074 1.103 0.142 1.147 ;
  END
END b15ztpn00an1d03x5

MACRO b15ztpn00an1n08x5
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN b15ztpn00an1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY Y ;
  SITE core ;
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
END b15ztpn00an1n08x5

END LIBRARY
